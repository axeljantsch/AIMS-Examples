/* Verilog module written by vlog2Verilog (qflow) */

module multiplierBeh(
    input [31:0] a,
    input [31:0] b,
    input clk,
    output [63:0] y
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _11689_ ;
wire _11269_ ;
wire _9837_ ;
wire _9417_ ;
wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _9590_ ;
wire _9170_ ;
wire [31:0] a ;
wire [31:0] b ;
wire _1677_ ;
wire _1257_ ;
wire _7903_ ;
wire [63:0] y ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _11901_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _10293_ ;
wire _4608_ ;
wire _8861_ ;
wire _8441_ ;
wire _8021_ ;
wire _11498_ ;
wire _11078_ ;
wire _9646_ ;
wire _9226_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _7712_ ;
wire _10769_ ;
wire _10349_ ;
wire _397_ ;
wire _11710_ ;
wire _8917_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _8670_ ;
wire _8250_ ;
wire _9875_ ;
wire _9455_ ;
wire _9035_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _7941_ ;
wire _7521_ ;
wire _7101_ ;
wire _10998_ ;
wire _10578_ ;
wire _10158_ ;
wire _8726_ ;
wire _8306_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _9684_ ;
wire _9264_ ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _7750_ ;
wire _7330_ ;
wire _10387_ ;
wire _8955_ ;
wire _8535_ ;
wire _8115_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _9493_ ;
wire _9073_ ;
wire _7806_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _11804_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _10196_ ;
wire _8764_ ;
wire _8344_ ;
wire _9969_ ;
wire _9549_ ;
wire _9129_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _7615_ ;
wire _2750_ ;
wire _2330_ ;
wire _11613_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _8993_ ;
wire _8573_ ;
wire _8153_ ;
wire _19_ ;
wire _1601_ ;
wire _9778_ ;
wire _9358_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _7844_ ;
wire _7424_ ;
wire _7004_ ;
wire _11842_ ;
wire _11422_ ;
wire _11002_ ;
wire _8629_ ;
wire _8209_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _8382_ ;
wire _1830_ ;
wire _1410_ ;
wire _9587_ ;
wire _9167_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _7653_ ;
wire _7233_ ;
wire _11651_ ;
wire _11231_ ;
wire _8858_ ;
wire _8438_ ;
wire _8018_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _8191_ ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire _9396_ ;
wire _10922_ ;
wire _10502_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _7709_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _11707_ ;
wire _3629_ ;
wire _3209_ ;
wire _7882_ ;
wire _7462_ ;
wire _7042_ ;
wire _10099_ ;
wire _11880_ ;
wire _11460_ ;
wire _11040_ ;
wire _8667_ ;
wire _8247_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _10731_ ;
wire _10311_ ;
wire _7938_ ;
wire _7518_ ;
wire _2653_ ;
wire _2233_ ;
wire _11516_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _7691_ ;
wire _7271_ ;
wire _8896_ ;
wire _8476_ ;
wire _8056_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _10960_ ;
wire _10540_ ;
wire _10120_ ;
wire _7747_ ;
wire _7327_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _11745_ ;
wire _11325_ ;
wire _3667_ ;
wire _3247_ ;
wire _7080_ ;
wire _5813_ ;
wire _8285_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6771_ ;
wire _6351_ ;
wire _7976_ ;
wire _7556_ ;
wire _7136_ ;
wire _2691_ ;
wire _2271_ ;
wire _11554_ ;
wire _11134_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _9702_ ;
wire _5622_ ;
wire _5202_ ;
wire _8094_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _9299_ ;
wire _10825_ ;
wire _10405_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _7785_ ;
wire _7365_ ;
wire _2080_ ;
wire _11783_ ;
wire _11363_ ;
wire _3285_ ;
wire _9931_ ;
wire _9511_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _10634_ ;
wire _10214_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _11839_ ;
wire _11419_ ;
wire _4702_ ;
wire _7594_ ;
wire _7174_ ;
wire _11592_ ;
wire _11172_ ;
wire _5907_ ;
wire _8799_ ;
wire _8379_ ;
wire _3094_ ;
wire _9740_ ;
wire _9320_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _10863_ ;
wire _10443_ ;
wire _10023_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _11648_ ;
wire _11228_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _8188_ ;
wire _1636_ ;
wire _1216_ ;
wire _10919_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _10672_ ;
wire _10252_ ;
wire _7879_ ;
wire _7459_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _8820_ ;
wire _8400_ ;
wire _11877_ ;
wire _11457_ ;
wire _11037_ ;
wire _3799_ ;
wire _3379_ ;
wire _9605_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _10728_ ;
wire _10308_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _10481_ ;
wire _10061_ ;
wire _7688_ ;
wire _7268_ ;
wire _11686_ ;
wire _11266_ ;
wire _3188_ ;
wire _9834_ ;
wire _9414_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _7900_ ;
wire _10957_ ;
wire _10537_ ;
wire _10117_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _10290_ ;
wire _4605_ ;
wire _7497_ ;
wire _7077_ ;
wire _11495_ ;
wire _11075_ ;
wire _9643_ ;
wire _9223_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire areg_25_bF$buf0 ;
wire areg_25_bF$buf1 ;
wire areg_25_bF$buf2 ;
wire areg_25_bF$buf3 ;
wire areg_25_bF$buf4 ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _10766_ ;
wire _10346_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _8914_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _9872_ ;
wire _9452_ ;
wire _9032_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _10995_ ;
wire _10575_ ;
wire _10155_ ;
wire _2497_ ;
wire _2077_ ;
wire _8723_ ;
wire _8303_ ;
wire _9928_ ;
wire _9508_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _9681_ ;
wire _9261_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire _10384_ ;
wire _8952_ ;
wire _8532_ ;
wire _8112_ ;
wire _11589_ ;
wire _11169_ ;
wire _9737_ ;
wire _9317_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _9490_ ;
wire _9070_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _7803_ ;
wire _488_ ;
wire _11801_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _10193_ ;
wire _4928_ ;
wire _4508_ ;
wire _8761_ ;
wire _8341_ ;
wire _11398_ ;
wire _9966_ ;
wire _9546_ ;
wire _9126_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _7612_ ;
wire _10669_ ;
wire _10249_ ;
wire _297_ ;
wire _11610_ ;
wire _8817_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire areg_7_bF$buf0 ;
wire areg_7_bF$buf1 ;
wire areg_7_bF$buf2 ;
wire areg_7_bF$buf3 ;
wire areg_7_bF$buf4 ;
wire _4737_ ;
wire _4317_ ;
wire _8990_ ;
wire _8570_ ;
wire _8150_ ;
wire _16_ ;
wire _9775_ ;
wire _9355_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7841_ ;
wire _7421_ ;
wire _7001_ ;
wire _10898_ ;
wire _10478_ ;
wire _10058_ ;
wire _8626_ ;
wire _8206_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _9584_ ;
wire _9164_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _7650_ ;
wire _7230_ ;
wire _10287_ ;
wire _8855_ ;
wire _8435_ ;
wire _8015_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire _9393_ ;
wire _7706_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _11704_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _10096_ ;
wire _8664_ ;
wire _8244_ ;
wire _9869_ ;
wire _9449_ ;
wire _9029_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _7935_ ;
wire _7515_ ;
wire _2650_ ;
wire _2230_ ;
wire _11513_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _8893_ ;
wire _8473_ ;
wire _8053_ ;
wire _1921_ ;
wire _1501_ ;
wire _9678_ ;
wire _9258_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _7744_ ;
wire _7324_ ;
wire _11742_ ;
wire _11322_ ;
wire _8949_ ;
wire _8529_ ;
wire _8109_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _8282_ ;
wire _1730_ ;
wire _1310_ ;
wire _9487_ ;
wire _9067_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _7973_ ;
wire _7553_ ;
wire _7133_ ;
wire _11551_ ;
wire _11131_ ;
wire _8758_ ;
wire _8338_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _8091_ ;
wire _6824_ ;
wire _6404_ ;
wire _9296_ ;
wire _10822_ ;
wire _10402_ ;
wire _870_ ;
wire _450_ ;
wire _7609_ ;
wire _2744_ ;
wire _2324_ ;
wire _11607_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _7782_ ;
wire _7362_ ;
wire _11780_ ;
wire _11360_ ;
wire _8987_ ;
wire _8567_ ;
wire _8147_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _10631_ ;
wire _10211_ ;
wire _7838_ ;
wire _7418_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _11836_ ;
wire _11416_ ;
wire _3758_ ;
wire _3338_ ;
wire _7591_ ;
wire _7171_ ;
wire _5904_ ;
wire _8796_ ;
wire _8376_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire _10860_ ;
wire _10440_ ;
wire _10020_ ;
wire _7647_ ;
wire _7227_ ;
wire _2782_ ;
wire _2362_ ;
wire _11645_ ;
wire _11225_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _8185_ ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire _10916_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _7876_ ;
wire _7456_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire _11874_ ;
wire _11454_ ;
wire _11034_ ;
wire _3796_ ;
wire _3376_ ;
wire _9602_ ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _9199_ ;
wire _10725_ ;
wire _10305_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _7685_ ;
wire _7265_ ;
wire _11683_ ;
wire _11263_ ;
wire _3185_ ;
wire _9831_ ;
wire _9411_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire breg_27_bF$buf0 ;
wire breg_27_bF$buf1 ;
wire breg_27_bF$buf2 ;
wire _89_ ;
wire breg_27_bF$buf3 ;
wire breg_27_bF$buf4 ;
wire _6956_ ;
wire breg_27_bF$buf5 ;
wire _6536_ ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _10954_ ;
wire _10534_ ;
wire _10114_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _11739_ ;
wire _11319_ ;
wire _4602_ ;
wire _7494_ ;
wire _7074_ ;
wire _11492_ ;
wire _11072_ ;
wire _5807_ ;
wire _8699_ ;
wire _8279_ ;
wire breg_5_bF$buf0 ;
wire breg_5_bF$buf1 ;
wire breg_5_bF$buf2 ;
wire breg_5_bF$buf3 ;
wire _9640_ ;
wire _9220_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _10763_ ;
wire _10343_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _8911_ ;
wire _11548_ ;
wire _11128_ ;
wire _3146__bF$buf0 ;
wire _3146__bF$buf1 ;
wire _3146__bF$buf2 ;
wire _3146__bF$buf3 ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _8088_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _10819_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _10992_ ;
wire _10572_ ;
wire _10152_ ;
wire _7779_ ;
wire _7359_ ;
wire _2494_ ;
wire _2074_ ;
wire _8720_ ;
wire _8300_ ;
wire _11777_ ;
wire _11357_ ;
wire _3699_ ;
wire _3279_ ;
wire _9925_ ;
wire _9505_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _10628_ ;
wire _10208_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _10381_ ;
wire _7588_ ;
wire _7168_ ;
wire _11586_ ;
wire _11166_ ;
wire _3088_ ;
wire _9734_ ;
wire _9314_ ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _7800_ ;
wire _10857_ ;
wire _10437_ ;
wire _10017_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _10190_ ;
wire _4925_ ;
wire _4505_ ;
wire _7397_ ;
wire _11395_ ;
wire _9963_ ;
wire _9543_ ;
wire _9123_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _10666_ ;
wire _10246_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _8814_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _9772_ ;
wire _9352_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _10895_ ;
wire _10475_ ;
wire _10055_ ;
wire _2397_ ;
wire _8623_ ;
wire _8203_ ;
wire _9828_ ;
wire _9408_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _9581_ ;
wire _9161_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _10284_ ;
wire _8852_ ;
wire _8432_ ;
wire _8012_ ;
wire _11489_ ;
wire _11069_ ;
wire _9637_ ;
wire _9217_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _9390_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _7703_ ;
wire _388_ ;
wire _11701_ ;
wire _8908_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _10093_ ;
wire _4828_ ;
wire _4408_ ;
wire _8661_ ;
wire _8241_ ;
wire _11298_ ;
wire _9866_ ;
wire _9446_ ;
wire _9026_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _7932_ ;
wire _7512_ ;
wire _10989_ ;
wire _10569_ ;
wire _10149_ ;
wire _197_ ;
wire _11510_ ;
wire _8717_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _8890_ ;
wire _8470_ ;
wire _8050_ ;
wire _9675_ ;
wire _9255_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _7741_ ;
wire _7321_ ;
wire _10798_ ;
wire _10378_ ;
wire _8946_ ;
wire _8526_ ;
wire _8106_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _9484_ ;
wire _9064_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _7970_ ;
wire _7550_ ;
wire _7130_ ;
wire _10187_ ;
wire _8755_ ;
wire _8335_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire areg_20_bF$buf0 ;
wire areg_20_bF$buf1 ;
wire areg_20_bF$buf2 ;
wire areg_20_bF$buf3 ;
wire areg_20_bF$buf4 ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _9293_ ;
wire _7606_ ;
wire _2741_ ;
wire _2321_ ;
wire _11604_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _8984_ ;
wire _8564_ ;
wire _8144_ ;
wire _9769_ ;
wire _9349_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _7835_ ;
wire _7415_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _11833_ ;
wire _11413_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _8793_ ;
wire _8373_ ;
wire _1821_ ;
wire _1401_ ;
wire _9998_ ;
wire _9578_ ;
wire _9158_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _7644_ ;
wire _7224_ ;
wire _11642_ ;
wire _11222_ ;
wire _8849_ ;
wire _8429_ ;
wire _8009_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _8182_ ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _9387_ ;
wire _10913_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _7873_ ;
wire _7453_ ;
wire _7033_ ;
wire _11871_ ;
wire _11451_ ;
wire _11031_ ;
wire _8658_ ;
wire _8238_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire areg_2_bF$buf0 ;
wire areg_2_bF$buf1 ;
wire areg_2_bF$buf2 ;
wire areg_2_bF$buf3 ;
wire areg_2_bF$buf4 ;
wire _6724_ ;
wire _6304_ ;
wire _9196_ ;
wire _10722_ ;
wire _10302_ ;
wire _770_ ;
wire _350_ ;
wire _7929_ ;
wire _7509_ ;
wire _2644_ ;
wire _2224_ ;
wire _11507_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _7682_ ;
wire _7262_ ;
wire _11680_ ;
wire _11260_ ;
wire _8887_ ;
wire _8467_ ;
wire _8047_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire _10951_ ;
wire _10531_ ;
wire _10111_ ;
wire _7738_ ;
wire _7318_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _11736_ ;
wire _11316_ ;
wire _3658_ ;
wire _3238_ ;
wire _7491_ ;
wire _7071_ ;
wire _5804_ ;
wire _8696_ ;
wire _8276_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _10760_ ;
wire _10340_ ;
wire _7967_ ;
wire _7547_ ;
wire _7127_ ;
wire _2682_ ;
wire _2262_ ;
wire _11545_ ;
wire _11125_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _8085_ ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _10816_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _7776_ ;
wire _7356_ ;
wire _2491_ ;
wire _2071_ ;
wire _11774_ ;
wire _11354_ ;
wire _3696_ ;
wire _3276_ ;
wire _9922_ ;
wire _9502_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire breg_19_bF$buf0 ;
wire _6627_ ;
wire breg_19_bF$buf1 ;
wire _6207_ ;
wire breg_19_bF$buf2 ;
wire breg_19_bF$buf3 ;
wire breg_19_bF$buf4 ;
wire _1762_ ;
wire breg_19_bF$buf5 ;
wire _1342_ ;
wire _9099_ ;
wire _10625_ ;
wire _10205_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _7585_ ;
wire _7165_ ;
wire _11583_ ;
wire _11163_ ;
wire _3085_ ;
wire _9731_ ;
wire _9311_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _10854_ ;
wire _10434_ ;
wire _10014_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _11639_ ;
wire _11219_ ;
wire _4922_ ;
wire _4502_ ;
wire _7394_ ;
wire _11392_ ;
wire _5707_ ;
wire _8599_ ;
wire _8179_ ;
wire _9960_ ;
wire _9540_ ;
wire _9120_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _10663_ ;
wire _10243_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _8811_ ;
wire _11868_ ;
wire _11448_ ;
wire _11028_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _10719_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _10892_ ;
wire _10472_ ;
wire _10052_ ;
wire _7679_ ;
wire _7259_ ;
wire _2394_ ;
wire _8620_ ;
wire _8200_ ;
wire _11677_ ;
wire _11257_ ;
wire _3599_ ;
wire _3179_ ;
wire _9825_ ;
wire _9405_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _10948_ ;
wire _10528_ ;
wire _10108_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _10281_ ;
wire _7488_ ;
wire _7068_ ;
wire _11486_ ;
wire _11066_ ;
wire _9634_ ;
wire _9214_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _7700_ ;
wire _10757_ ;
wire _10337_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _8905_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4116__bF$buf0 ;
wire _4116__bF$buf1 ;
wire _4116__bF$buf2 ;
wire _4116__bF$buf3 ;
wire _4116__bF$buf4 ;
wire _10090_ ;
wire _4825_ ;
wire _4405_ ;
wire _7297_ ;
wire _11295_ ;
wire _9863_ ;
wire _9443_ ;
wire _9023_ ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _10986_ ;
wire _10566_ ;
wire _10146_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _8714_ ;
wire _9919_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _9672_ ;
wire _9252_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _10795_ ;
wire _10375_ ;
wire _2297_ ;
wire _8943_ ;
wire _8523_ ;
wire _8103_ ;
wire breg_22_bF$buf0 ;
wire breg_22_bF$buf1 ;
wire breg_22_bF$buf2 ;
wire breg_22_bF$buf3 ;
wire breg_22_bF$buf4 ;
wire _9728_ ;
wire _9308_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _9481_ ;
wire _9061_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire breg_0_bF$buf0 ;
wire breg_0_bF$buf1 ;
wire breg_0_bF$buf2 ;
wire breg_0_bF$buf3 ;
wire breg_0_bF$buf4 ;
wire _3714_ ;
wire breg_0_bF$buf5 ;
wire breg_0_bF$buf6 ;
wire _6186_ ;
wire _10184_ ;
wire _4919_ ;
wire _8752_ ;
wire _8332_ ;
wire _11389_ ;
wire _9957_ ;
wire _9537_ ;
wire _9117_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _9290_ ;
wire _1797_ ;
wire _1377_ ;
wire _7603_ ;
wire _288_ ;
wire _11601_ ;
wire _8808_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _8981_ ;
wire _8561_ ;
wire _8141_ ;
wire _11198_ ;
wire _9766_ ;
wire _9346_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _7832_ ;
wire _7412_ ;
wire _10889_ ;
wire _10469_ ;
wire _10049_ ;
wire _11830_ ;
wire _11410_ ;
wire _8617_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _8790_ ;
wire _8370_ ;
wire _9995_ ;
wire _9575_ ;
wire _9155_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _7641_ ;
wire _7221_ ;
wire _10698_ ;
wire _10278_ ;
wire _8846_ ;
wire _8426_ ;
wire _8006_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire areg_31_bF$buf0 ;
wire areg_31_bF$buf1 ;
wire areg_31_bF$buf2 ;
wire areg_31_bF$buf3 ;
wire areg_31_bF$buf4 ;
wire _45_ ;
wire _6912_ ;
wire _9384_ ;
wire _10910_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire _7870_ ;
wire _7450_ ;
wire _7030_ ;
wire _10087_ ;
wire _8655_ ;
wire _8235_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _9193_ ;
wire _7926_ ;
wire _7506_ ;
wire _2641_ ;
wire _2221_ ;
wire _11504_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _8884_ ;
wire _8464_ ;
wire _8044_ ;
wire _1912_ ;
wire _9669_ ;
wire _9249_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5315__bF$buf0 ;
wire _5589_ ;
wire _5315__bF$buf1 ;
wire _5169_ ;
wire _5315__bF$buf2 ;
wire _5315__bF$buf3 ;
wire _5315__bF$buf4 ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _7735_ ;
wire _7315_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _11733_ ;
wire _11313_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _8693_ ;
wire _8273_ ;
wire _1721_ ;
wire _1301_ ;
wire _9898_ ;
wire _9478_ ;
wire _9058_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _7964_ ;
wire _7544_ ;
wire _7124_ ;
wire _11542_ ;
wire _11122_ ;
wire _8749_ ;
wire _8329_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _8082_ ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _9287_ ;
wire _10813_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _7773_ ;
wire _7353_ ;
wire _11771_ ;
wire _11351_ ;
wire _8978_ ;
wire _8558_ ;
wire _8138_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _9096_ ;
wire _10622_ ;
wire _10202_ ;
wire _670_ ;
wire _250_ ;
wire _7829_ ;
wire _7409_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _11827_ ;
wire _11407_ ;
wire _3749_ ;
wire _3329_ ;
wire _7582_ ;
wire _7162_ ;
wire _11580_ ;
wire _11160_ ;
wire _8787_ ;
wire _8367_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire _10851_ ;
wire _10431_ ;
wire _10011_ ;
wire _7638_ ;
wire _7218_ ;
wire _2773_ ;
wire _2353_ ;
wire _11636_ ;
wire _11216_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _7391_ ;
wire _5704_ ;
wire _8596_ ;
wire _8176_ ;
wire _5453__bF$buf0 ;
wire _5453__bF$buf1 ;
wire _5453__bF$buf2 ;
wire _5453__bF$buf3 ;
wire _5453__bF$buf4 ;
wire _5453__bF$buf5 ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _10907_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _10660_ ;
wire _10240_ ;
wire _7867_ ;
wire _7447_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _11865_ ;
wire _11445_ ;
wire _11025_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _10716_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire _7676_ ;
wire _7256_ ;
wire _2391_ ;
wire _11674_ ;
wire _11254_ ;
wire _3596_ ;
wire _3176_ ;
wire _9822_ ;
wire _9402_ ;
wire _2287__bF$buf0 ;
wire _2287__bF$buf1 ;
wire _2287__bF$buf2 ;
wire _2287__bF$buf3 ;
wire _1909_ ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _10945_ ;
wire _10525_ ;
wire _10105_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _7485_ ;
wire _7065_ ;
wire _11483_ ;
wire _11063_ ;
wire _9631_ ;
wire _9211_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _10754_ ;
wire _10334_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _8902_ ;
wire _11539_ ;
wire _11119_ ;
wire _4822_ ;
wire _4402_ ;
wire _7294_ ;
wire _11292_ ;
wire _5607_ ;
wire _8499_ ;
wire _8079_ ;
wire _9860_ ;
wire _9440_ ;
wire _9020_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _10983_ ;
wire _10563_ ;
wire _10143_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _8711_ ;
wire _11768_ ;
wire _11348_ ;
wire _9916_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _10619_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _10792_ ;
wire _10372_ ;
wire _7999_ ;
wire _7579_ ;
wire _7159_ ;
wire _2294_ ;
wire _8940_ ;
wire _8520_ ;
wire _8100_ ;
wire _11577_ ;
wire _11157_ ;
wire _3499_ ;
wire _3079_ ;
wire _9725_ ;
wire _9305_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _4434__bF$buf0 ;
wire _4434__bF$buf1 ;
wire _4434__bF$buf2 ;
wire _4434__bF$buf3 ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _10848_ ;
wire _10428_ ;
wire _10008_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _10181_ ;
wire _4916_ ;
wire _7388_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _11386_ ;
wire _9954_ ;
wire _9534_ ;
wire _9114_ ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _7600_ ;
wire _10657_ ;
wire _10237_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _8805_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _7197_ ;
wire _11195_ ;
wire _9763_ ;
wire _9343_ ;
wire _5683_ ;
wire _5263_ ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _10886_ ;
wire _10466_ ;
wire _10046_ ;
wire _2388_ ;
wire _8614_ ;
wire breg_14_bF$buf0 ;
wire breg_14_bF$buf1 ;
wire breg_14_bF$buf2 ;
wire breg_14_bF$buf3 ;
wire _9819_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _9992_ ;
wire _9572_ ;
wire _9152_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _10695_ ;
wire _10275_ ;
wire _2197_ ;
wire _8843_ ;
wire _8423_ ;
wire _8003_ ;
wire _9628_ ;
wire _9208_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _9381_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _10084_ ;
wire _4819_ ;
wire _8652_ ;
wire _8232_ ;
wire _11289_ ;
wire _9857_ ;
wire _9437_ ;
wire _9017_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _9190_ ;
wire _1697_ ;
wire _1277_ ;
wire _7923_ ;
wire _7503_ ;
wire _188_ ;
wire _11501_ ;
wire _8708_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _8881_ ;
wire _8461_ ;
wire _8041_ ;
wire _11098_ ;
wire _9666_ ;
wire _9246_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _7732_ ;
wire _7312_ ;
wire _10789_ ;
wire _10369_ ;
wire _11730_ ;
wire _11310_ ;
wire _8937_ ;
wire _8517_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _8690_ ;
wire _8270_ ;
wire _9895_ ;
wire _9475_ ;
wire _9055_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _7961_ ;
wire _7541_ ;
wire _7121_ ;
wire _10598_ ;
wire _10178_ ;
wire _2586__bF$buf0 ;
wire _2586__bF$buf1 ;
wire _2586__bF$buf2 ;
wire _2586__bF$buf3 ;
wire _2586__bF$buf4 ;
wire _8746_ ;
wire _8326_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _6812_ ;
wire _9284_ ;
wire _10810_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _7770_ ;
wire _7350_ ;
wire _8975_ ;
wire _8555_ ;
wire _8135_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _9093_ ;
wire _7826_ ;
wire _7406_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _11824_ ;
wire _11404_ ;
wire _3746_ ;
wire _3326_ ;
wire _8784_ ;
wire _8364_ ;
wire _1812_ ;
wire _9989_ ;
wire _9569_ ;
wire _9149_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire _7635_ ;
wire _7215_ ;
wire _2770_ ;
wire _2350_ ;
wire _11633_ ;
wire _11213_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _8593_ ;
wire _8173_ ;
wire _39_ ;
wire _6906_ ;
wire _1621_ ;
wire _1201_ ;
wire _9798_ ;
wire _9378_ ;
wire _4093_ ;
wire _10904_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _7864_ ;
wire _7444_ ;
wire _7024_ ;
wire _11862_ ;
wire _11442_ ;
wire _11022_ ;
wire _8649_ ;
wire _8229_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _9187_ ;
wire _10713_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire _7673_ ;
wire _7253_ ;
wire clk ;
wire _11671_ ;
wire _11251_ ;
wire _8878_ ;
wire _8458_ ;
wire _8038_ ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _10942_ ;
wire _10522_ ;
wire _10102_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _7729_ ;
wire _7309_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _11727_ ;
wire _11307_ ;
wire _3649_ ;
wire _3229_ ;
wire _7225__bF$buf0 ;
wire _7225__bF$buf1 ;
wire _7225__bF$buf2 ;
wire _7225__bF$buf3 ;
wire _7225__bF$buf4 ;
wire _7482_ ;
wire _7062_ ;
wire _11480_ ;
wire _11060_ ;
wire _8687_ ;
wire _8267_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _10751_ ;
wire _10331_ ;
wire _7958_ ;
wire _7538_ ;
wire _7118_ ;
wire _2673_ ;
wire _2253_ ;
wire areg_16_bF$buf0 ;
wire areg_16_bF$buf1 ;
wire areg_16_bF$buf2 ;
wire areg_16_bF$buf3 ;
wire areg_16_bF$buf4 ;
wire areg_16_bF$buf5 ;
wire _11536_ ;
wire _11116_ ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _7291_ ;
wire _5604_ ;
wire _8496_ ;
wire _8076_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _10807_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire _10980_ ;
wire _10560_ ;
wire _10140_ ;
wire _7767_ ;
wire _7347_ ;
wire _2482_ ;
wire _2062_ ;
wire _11765_ ;
wire _11345_ ;
wire _3687_ ;
wire _3267_ ;
wire _9913_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _10616_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _7996_ ;
wire _7576_ ;
wire _7156_ ;
wire _2291_ ;
wire _11574_ ;
wire _11154_ ;
wire _3496_ ;
wire _3076_ ;
wire _9722_ ;
wire _9302_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _10845_ ;
wire _10425_ ;
wire _10005_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _7385_ ;
wire _11383_ ;
wire _9951_ ;
wire _9531_ ;
wire _9111_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _10654_ ;
wire _10234_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _8802_ ;
wire _11859_ ;
wire _11439_ ;
wire _11019_ ;
wire _4722_ ;
wire _4302_ ;
wire _7194_ ;
wire _11192_ ;
wire _5927_ ;
wire _5507_ ;
wire _8399_ ;
wire _9760_ ;
wire _9340_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _10883_ ;
wire _10463_ ;
wire _10043_ ;
wire _2385_ ;
wire _8611_ ;
wire _11668_ ;
wire _11248_ ;
wire _9816_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _10939_ ;
wire _10519_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _10692_ ;
wire _10272_ ;
wire _7899_ ;
wire _7479_ ;
wire _7059_ ;
wire _2194_ ;
wire _8840_ ;
wire _8420_ ;
wire _8000_ ;
wire _11897_ ;
wire _11477_ ;
wire _11057_ ;
wire _3399_ ;
wire _9625_ ;
wire _9205_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _10748_ ;
wire _10328_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _10081_ ;
wire _4816_ ;
wire _7288_ ;
wire _11286_ ;
wire _9854_ ;
wire _9434_ ;
wire _9014_ ;
wire _5774_ ;
wire _5354_ ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _7920_ ;
wire _7500_ ;
wire _10977_ ;
wire _10557_ ;
wire _10137_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _8705_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire _7097_ ;
wire _11095_ ;
wire _9663_ ;
wire _9243_ ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _10786_ ;
wire _10366_ ;
wire _2288_ ;
wire _8934_ ;
wire _8514_ ;
wire _9719_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _9892_ ;
wire _9472_ ;
wire _9052_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _10595_ ;
wire _10175_ ;
wire _2097_ ;
wire _8743_ ;
wire _8323_ ;
wire _9948_ ;
wire _9528_ ;
wire _9108_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _9281_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _8972_ ;
wire _8552_ ;
wire _8132_ ;
wire _11189_ ;
wire _9757_ ;
wire _9337_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _9090_ ;
wire _1597_ ;
wire _1177_ ;
wire _7823_ ;
wire _7403_ ;
wire _11821_ ;
wire _11401_ ;
wire _8608_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _8781_ ;
wire _8361_ ;
wire _9986_ ;
wire _9566_ ;
wire _9146_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _7632_ ;
wire _7212_ ;
wire _10689_ ;
wire _10269_ ;
wire _11630_ ;
wire _11210_ ;
wire _8837_ ;
wire _8417_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _8590_ ;
wire _8170_ ;
wire _36_ ;
wire _6903_ ;
wire _9795_ ;
wire _9375_ ;
wire _4090_ ;
wire _10901_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _7861_ ;
wire _7441_ ;
wire _7021_ ;
wire _10498_ ;
wire _10078_ ;
wire _8646_ ;
wire _8226_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _9184_ ;
wire _10710_ ;
wire _7917_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _7670_ ;
wire _7250_ ;
wire _8875_ ;
wire _8455_ ;
wire _8035_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _7726_ ;
wire _7306_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _11724_ ;
wire _11304_ ;
wire _3646_ ;
wire _3226_ ;
wire _2376__bF$buf0 ;
wire _2376__bF$buf1 ;
wire _2376__bF$buf2 ;
wire _2376__bF$buf3 ;
wire _8684_ ;
wire _8264_ ;
wire _1712_ ;
wire _9889_ ;
wire _9469_ ;
wire _9049_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _7955_ ;
wire _7535_ ;
wire _7115_ ;
wire _2670_ ;
wire _2250_ ;
wire _11533_ ;
wire _11113_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire _5601_ ;
wire _8493_ ;
wire _8073_ ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _9698_ ;
wire _9278_ ;
wire _10804_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _7764_ ;
wire _7344_ ;
wire _11762_ ;
wire _11342_ ;
wire _8969_ ;
wire _8549_ ;
wire _8129_ ;
wire _3684_ ;
wire _3264_ ;
wire _9910_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _9087_ ;
wire _10613_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _11818_ ;
wire _7993_ ;
wire _7573_ ;
wire _7153_ ;
wire _11571_ ;
wire _11151_ ;
wire _8778_ ;
wire _8358_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _10842_ ;
wire _10422_ ;
wire _10002_ ;
wire _890_ ;
wire _470_ ;
wire _7629_ ;
wire _7209_ ;
wire _2764_ ;
wire _2344_ ;
wire _11627_ ;
wire _11207_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire areg_27_bF$buf0 ;
wire areg_27_bF$buf1 ;
wire areg_27_bF$buf2 ;
wire areg_27_bF$buf3 ;
wire areg_27_bF$buf4 ;
wire areg_27_bF$buf5 ;
wire _7382_ ;
wire _11380_ ;
wire _8587_ ;
wire _8167_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _10651_ ;
wire _10231_ ;
wire _7858_ ;
wire _7438_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _11856_ ;
wire _11436_ ;
wire _11016_ ;
wire _3778_ ;
wire _3358_ ;
wire _7191_ ;
wire _5924_ ;
wire _5504_ ;
wire _8396_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _10707_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire _10880_ ;
wire _10460_ ;
wire _10040_ ;
wire _7667_ ;
wire _7247_ ;
wire _2382_ ;
wire _11665_ ;
wire _11245_ ;
wire _3587_ ;
wire _3167_ ;
wire _9813_ ;
wire _5733_ ;
wire _5313_ ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _10936_ ;
wire _10516_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7896_ ;
wire _7476_ ;
wire _7056_ ;
wire _2191_ ;
wire _11894_ ;
wire _11474_ ;
wire _11054_ ;
wire _3396_ ;
wire _9622_ ;
wire _9202_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _10745_ ;
wire _10325_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _7285_ ;
wire _11283_ ;
wire _9851_ ;
wire _9431_ ;
wire _9011_ ;
wire areg_9_bF$buf0 ;
wire areg_9_bF$buf1 ;
wire areg_9_bF$buf2 ;
wire areg_9_bF$buf3 ;
wire areg_9_bF$buf4 ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _10974_ ;
wire _10554_ ;
wire _10134_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _8702_ ;
wire _11759_ ;
wire _11339_ ;
wire _9907_ ;
wire _4622_ ;
wire _4202_ ;
wire _7094_ ;
wire _11092_ ;
wire _5827_ ;
wire _5407_ ;
wire _8299_ ;
wire _9660_ ;
wire _9240_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _10783_ ;
wire _10363_ ;
wire _2285_ ;
wire _8931_ ;
wire _8511_ ;
wire _11568_ ;
wire _11148_ ;
wire _9716_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _10839_ ;
wire _10419_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _10592_ ;
wire _10172_ ;
wire _4907_ ;
wire _7799_ ;
wire _7379_ ;
wire _2094_ ;
wire _8740_ ;
wire _8320_ ;
wire _11797_ ;
wire _11377_ ;
wire _3299_ ;
wire _9945_ ;
wire _9525_ ;
wire _9105_ ;
wire _4660_ ;
wire _4240_ ;
wire areg_11_bF$buf0 ;
wire areg_11_bF$buf1 ;
wire areg_11_bF$buf2 ;
wire areg_11_bF$buf3 ;
wire _5865_ ;
wire areg_11_bF$buf4 ;
wire _5445_ ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _10648_ ;
wire _10228_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _7188_ ;
wire _11186_ ;
wire _9754_ ;
wire _9334_ ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _7820_ ;
wire _7400_ ;
wire _10877_ ;
wire _10457_ ;
wire _10037_ ;
wire _2799_ ;
wire _2379_ ;
wire _8605_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire _9983_ ;
wire _9563_ ;
wire _9143_ ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _10686_ ;
wire _10266_ ;
wire _2188_ ;
wire _8834_ ;
wire _8414_ ;
wire _9619_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _6900_ ;
wire _9792_ ;
wire _9372_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _10495_ ;
wire _10075_ ;
wire _8643_ ;
wire _8223_ ;
wire _9848_ ;
wire _9428_ ;
wire _9008_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _9181_ ;
wire _1688_ ;
wire _1268_ ;
wire _7914_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _8872_ ;
wire _8452_ ;
wire _8032_ ;
wire _11089_ ;
wire _1900_ ;
wire _9657_ ;
wire _9237_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _7723_ ;
wire _7303_ ;
wire _11721_ ;
wire _11301_ ;
wire _8928_ ;
wire _8508_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _8681_ ;
wire _8261_ ;
wire _9886_ ;
wire _9466_ ;
wire _9046_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _7952_ ;
wire _7532_ ;
wire _7112_ ;
wire _10589_ ;
wire _10169_ ;
wire _11530_ ;
wire _11110_ ;
wire _8737_ ;
wire _8317_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _8490_ ;
wire _8070_ ;
wire _6803_ ;
wire _9695_ ;
wire _9275_ ;
wire _10801_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _7761_ ;
wire _7341_ ;
wire _10398_ ;
wire _8966_ ;
wire _8546_ ;
wire _8126_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _9084_ ;
wire _10610_ ;
wire _7817_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _11815_ ;
wire _3737_ ;
wire _3317_ ;
wire breg_29_bF$buf0 ;
wire breg_29_bF$buf1 ;
wire breg_29_bF$buf2 ;
wire breg_29_bF$buf3 ;
wire breg_29_bF$buf4 ;
wire _7990_ ;
wire _7570_ ;
wire _7150_ ;
wire _8775_ ;
wire _8355_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire breg_7_bF$buf0 ;
wire breg_7_bF$buf1 ;
wire breg_7_bF$buf2 ;
wire breg_7_bF$buf3 ;
wire breg_7_bF$buf4 ;
wire breg_7_bF$buf5 ;
wire _7626_ ;
wire _7206_ ;
wire _2761_ ;
wire _2341_ ;
wire _11624_ ;
wire _11204_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _8584_ ;
wire _8164_ ;
wire _1612_ ;
wire _9789_ ;
wire _9369_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7855_ ;
wire _7435_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _11853_ ;
wire _11433_ ;
wire _11013_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _8393_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _9598_ ;
wire _9178_ ;
wire _10704_ ;
wire _5190__bF$buf0 ;
wire _5190__bF$buf1 ;
wire _5190__bF$buf2 ;
wire _5190__bF$buf3 ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire [63:0] _11909_ ;
wire _7664_ ;
wire _7244_ ;
wire _11662_ ;
wire _11242_ ;
wire _8869_ ;
wire _8449_ ;
wire _8029_ ;
wire _3584_ ;
wire _3164_ ;
wire _9810_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _10933_ ;
wire _10513_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _11718_ ;
wire _7893_ ;
wire _7473_ ;
wire _7053_ ;
wire _11891_ ;
wire _11471_ ;
wire _11051_ ;
wire _8678_ ;
wire _8258_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _10742_ ;
wire _10322_ ;
wire _790_ ;
wire _370_ ;
wire _7949_ ;
wire _7529_ ;
wire _7109_ ;
wire _2664_ ;
wire _2244_ ;
wire _11527_ ;
wire _11107_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _7282_ ;
wire _11280_ ;
wire _8487_ ;
wire _8067_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _10971_ ;
wire _10551_ ;
wire _10131_ ;
wire _7758_ ;
wire _7338_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _11756_ ;
wire _11336_ ;
wire _3678_ ;
wire _3258_ ;
wire _9904_ ;
wire _7091_ ;
wire _5824_ ;
wire _5404_ ;
wire _8296_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _10607_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _10780_ ;
wire _10360_ ;
wire _7987_ ;
wire _7567_ ;
wire _7147_ ;
wire _2282_ ;
wire _11565_ ;
wire _11145_ ;
wire _3487_ ;
wire _3067_ ;
wire _9713_ ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _10836_ ;
wire _10416_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _7796_ ;
wire _7376_ ;
wire _2091_ ;
wire _11794_ ;
wire _11374_ ;
wire _3296_ ;
wire _9942_ ;
wire _9522_ ;
wire _9102_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _10645_ ;
wire _10225_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _7185_ ;
wire _11183_ ;
wire _5918_ ;
wire _9751_ ;
wire _9331_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire _10874_ ;
wire _10454_ ;
wire _10034_ ;
wire _2796_ ;
wire _2376_ ;
wire _8602_ ;
wire _11659_ ;
wire _11239_ ;
wire _9807_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _8199_ ;
wire _9980_ ;
wire _9560_ ;
wire _9140_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _10683_ ;
wire _10263_ ;
wire _2185_ ;
wire _8831_ ;
wire _8411_ ;
wire _11888_ ;
wire _11468_ ;
wire _11048_ ;
wire _9616_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire areg_22_bF$buf0 ;
wire areg_22_bF$buf1 ;
wire _1876_ ;
wire areg_22_bF$buf2 ;
wire _1456_ ;
wire areg_22_bF$buf3 ;
wire _1036_ ;
wire areg_22_bF$buf4 ;
wire _10739_ ;
wire _10319_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _10492_ ;
wire _10072_ ;
wire _4807_ ;
wire _7699_ ;
wire _7279_ ;
wire _8640_ ;
wire _8220_ ;
wire _11697_ ;
wire _11277_ ;
wire _3199_ ;
wire _9845_ ;
wire _9425_ ;
wire _9005_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _7911_ ;
wire _10968_ ;
wire _10548_ ;
wire _10128_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _7088_ ;
wire _11086_ ;
wire _9654_ ;
wire _9234_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _7720_ ;
wire _7300_ ;
wire _10777_ ;
wire _10357_ ;
wire _2699_ ;
wire _2279_ ;
wire _8925_ ;
wire _8505_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _9883_ ;
wire _9463_ ;
wire _9043_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire _10586_ ;
wire _10166_ ;
wire _2088_ ;
wire _8734_ ;
wire _8314_ ;
wire _9939_ ;
wire _9519_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _9692_ ;
wire _9272_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire areg_4_bF$buf0 ;
wire areg_4_bF$buf1 ;
wire areg_4_bF$buf2 ;
wire areg_4_bF$buf3 ;
wire areg_4_bF$buf4 ;
wire _10395_ ;
wire _8963_ ;
wire _8543_ ;
wire _8123_ ;
wire _9748_ ;
wire _9328_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _9081_ ;
wire _1588_ ;
wire _1168_ ;
wire _7814_ ;
wire _499_ ;
wire _11812_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _8772_ ;
wire _8352_ ;
wire _1800_ ;
wire _9977_ ;
wire _9557_ ;
wire _9137_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _7623_ ;
wire _7203_ ;
wire _11621_ ;
wire _11201_ ;
wire _8828_ ;
wire _8408_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _8581_ ;
wire _8161_ ;
wire _27_ ;
wire _9786_ ;
wire _9366_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _7852_ ;
wire _7432_ ;
wire _7012_ ;
wire _10489_ ;
wire _10069_ ;
wire _11850_ ;
wire _11430_ ;
wire _11010_ ;
wire _8637_ ;
wire _8217_ ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _8390_ ;
wire _6703_ ;
wire _9595_ ;
wire _9175_ ;
wire _10701_ ;
wire _7908_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _11906_ ;
wire _3828_ ;
wire _3408_ ;
wire _7661_ ;
wire _7241_ ;
wire _10298_ ;
wire _8866_ ;
wire _8446_ ;
wire _8026_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _10930_ ;
wire _10510_ ;
wire _7717_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _11715_ ;
wire _3637_ ;
wire _3217_ ;
wire _7890_ ;
wire _7470_ ;
wire _7050_ ;
wire _8675_ ;
wire _8255_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _7946_ ;
wire _7526_ ;
wire _7106_ ;
wire _2661_ ;
wire _2241_ ;
wire _11524_ ;
wire _11104_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _8484_ ;
wire _8064_ ;
wire _1932_ ;
wire _1512_ ;
wire _9689_ ;
wire _9269_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _7755_ ;
wire _7335_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _11753_ ;
wire _11333_ ;
wire _3675_ ;
wire _3255_ ;
wire _9901_ ;
wire _5821_ ;
wire _5401_ ;
wire _8293_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _9498_ ;
wire _9078_ ;
wire _10604_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _11809_ ;
wire _7984_ ;
wire _7564_ ;
wire _7144_ ;
wire _11562_ ;
wire _11142_ ;
wire _8769_ ;
wire _8349_ ;
wire _3484_ ;
wire _3064_ ;
wire _9710_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _10833_ ;
wire _10413_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _11618_ ;
wire _4901_ ;
wire _7793_ ;
wire _7373_ ;
wire _11791_ ;
wire _11371_ ;
wire _8998_ ;
wire _8578_ ;
wire _8158_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _10642_ ;
wire _10222_ ;
wire _690_ ;
wire _270_ ;
wire _7849_ ;
wire _7429_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _11847_ ;
wire _11427_ ;
wire _11007_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _7182_ ;
wire _11180_ ;
wire _5915_ ;
wire _8387_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire _10871_ ;
wire _10451_ ;
wire _10031_ ;
wire _7658_ ;
wire _7238_ ;
wire _2793_ ;
wire _2373_ ;
wire _11656_ ;
wire _11236_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _9804_ ;
wire _5724_ ;
wire _5304_ ;
wire _8196_ ;
wire _6929_ ;
wire _6509_ ;
wire breg_24_bF$buf0 ;
wire breg_24_bF$buf1 ;
wire _1644_ ;
wire breg_24_bF$buf2 ;
wire _1224_ ;
wire breg_24_bF$buf3 ;
wire breg_24_bF$buf4 ;
wire breg_24_bF$buf5 ;
wire _10927_ ;
wire _10507_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _10680_ ;
wire _10260_ ;
wire _7887_ ;
wire _7467_ ;
wire _7047_ ;
wire _2182_ ;
wire _11885_ ;
wire _11465_ ;
wire _11045_ ;
wire _3387_ ;
wire breg_2_bF$buf0 ;
wire breg_2_bF$buf1 ;
wire _9613_ ;
wire breg_2_bF$buf2 ;
wire breg_2_bF$buf3 ;
wire breg_2_bF$buf4 ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _10736_ ;
wire _10316_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _7696_ ;
wire _7276_ ;
wire _11694_ ;
wire _11274_ ;
wire _3196_ ;
wire _9842_ ;
wire _9422_ ;
wire _9002_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _10965_ ;
wire _10545_ ;
wire _10125_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _7085_ ;
wire _11083_ ;
wire _5818_ ;
wire _9651_ ;
wire _9231_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _10774_ ;
wire _10354_ ;
wire _2696_ ;
wire _2276_ ;
wire _8922_ ;
wire _8502_ ;
wire _11559_ ;
wire _11139_ ;
wire _9707_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _8099_ ;
wire _9880_ ;
wire _9460_ ;
wire _9040_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _10583_ ;
wire _10163_ ;
wire _2085_ ;
wire _8731_ ;
wire _8311_ ;
wire _11788_ ;
wire _11368_ ;
wire _9936_ ;
wire _9516_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _10639_ ;
wire _10219_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _10392_ ;
wire _4707_ ;
wire _7599_ ;
wire _7179_ ;
wire _8960_ ;
wire _8540_ ;
wire _8120_ ;
wire _11597_ ;
wire _11177_ ;
wire _3099_ ;
wire _9745_ ;
wire _9325_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _7811_ ;
wire _10868_ ;
wire _10448_ ;
wire _10028_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _9974_ ;
wire _9554_ ;
wire _9134_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _7620_ ;
wire _7200_ ;
wire _10677_ ;
wire _10257_ ;
wire _2599_ ;
wire _2179_ ;
wire _8825_ ;
wire _8405_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _9783_ ;
wire _9363_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _10486_ ;
wire _10066_ ;
wire _8634_ ;
wire _8214_ ;
wire _9839_ ;
wire _9419_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _9592_ ;
wire _9172_ ;
wire _1679_ ;
wire _1259_ ;
wire _7905_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _11903_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _10295_ ;
wire _8863_ ;
wire _8443_ ;
wire _8023_ ;
wire _9648_ ;
wire _9228_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _7714_ ;
wire _399_ ;
wire _11712_ ;
wire _8919_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _8672_ ;
wire _8252_ ;
wire _1700_ ;
wire _9877_ ;
wire _9457_ ;
wire _9037_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _7943_ ;
wire _7523_ ;
wire _7103_ ;
wire _11521_ ;
wire _11101_ ;
wire _8728_ ;
wire _8308_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _8481_ ;
wire _8061_ ;
wire _9686_ ;
wire _9266_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _7752_ ;
wire _7332_ ;
wire _10389_ ;
wire _11750_ ;
wire _11330_ ;
wire _8957_ ;
wire _8537_ ;
wire _8117_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _8290_ ;
wire _6603_ ;
wire _9495_ ;
wire _9075_ ;
wire _10601_ ;
wire _7808_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _11806_ ;
wire _3728_ ;
wire _3308_ ;
wire _7981_ ;
wire _7561_ ;
wire _7141_ ;
wire _10198_ ;
wire _8766_ ;
wire _8346_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _10830_ ;
wire _10410_ ;
wire _7617_ ;
wire _2752_ ;
wire _2332_ ;
wire _11615_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _7790_ ;
wire _7370_ ;
wire _8995_ ;
wire _8575_ ;
wire _8155_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire _7846_ ;
wire _7426_ ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _11844_ ;
wire _11424_ ;
wire _11004_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _8384_ ;
wire _1832_ ;
wire _1412_ ;
wire _9589_ ;
wire _9169_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire _7655_ ;
wire _7235_ ;
wire _2790_ ;
wire _2370_ ;
wire _11653_ ;
wire _11233_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _9801_ ;
wire _5721_ ;
wire _5301_ ;
wire _8193_ ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _9398_ ;
wire _10924_ ;
wire _10504_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _11709_ ;
wire _7884_ ;
wire _7464_ ;
wire _7044_ ;
wire _11882_ ;
wire _11462_ ;
wire _11042_ ;
wire _8669_ ;
wire _8249_ ;
wire _3384_ ;
wire _9610_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _10733_ ;
wire _10313_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _11518_ ;
wire _2669__bF$buf0 ;
wire _2669__bF$buf1 ;
wire _2669__bF$buf2 ;
wire _2669__bF$buf3 ;
wire _4801_ ;
wire _7693_ ;
wire _7273_ ;
wire _11691_ ;
wire _11271_ ;
wire _8898_ ;
wire _8478_ ;
wire _8058_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _10962_ ;
wire _10542_ ;
wire _10122_ ;
wire _590_ ;
wire _170_ ;
wire _7749_ ;
wire _7329_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _11747_ ;
wire _11327_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _7082_ ;
wire _11080_ ;
wire _5815_ ;
wire _8287_ ;
wire _1735_ ;
wire _1315_ ;
wire breg_16_bF$buf0 ;
wire breg_16_bF$buf1 ;
wire breg_16_bF$buf2 ;
wire breg_16_bF$buf3 ;
wire breg_16_bF$buf4 ;
wire breg_16_bF$buf5 ;
wire _646_ ;
wire _226_ ;
wire _6773_ ;
wire _6353_ ;
wire _10771_ ;
wire _10351_ ;
wire _7978_ ;
wire _7558_ ;
wire _7138_ ;
wire _2693_ ;
wire _2273_ ;
wire _11556_ ;
wire _11136_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _9704_ ;
wire _5624_ ;
wire _5204_ ;
wire _8096_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _10827_ ;
wire _10407_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _10580_ ;
wire _10160_ ;
wire _7787_ ;
wire _7367_ ;
wire _2082_ ;
wire _11785_ ;
wire _11365_ ;
wire _3287_ ;
wire _9933_ ;
wire _9513_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _10636_ ;
wire _10216_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire _7596_ ;
wire _7176_ ;
wire _11594_ ;
wire _11174_ ;
wire _5909_ ;
wire _3096_ ;
wire _9742_ ;
wire _9322_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _10865_ ;
wire _10445_ ;
wire _10025_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _9971_ ;
wire _9551_ ;
wire _9131_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _10674_ ;
wire _10254_ ;
wire _2596_ ;
wire _2176_ ;
wire _8822_ ;
wire _8402_ ;
wire _11879_ ;
wire _11459_ ;
wire _11039_ ;
wire _9607_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _9780_ ;
wire _9360_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _10483_ ;
wire _10063_ ;
wire _8631_ ;
wire _8211_ ;
wire _11688_ ;
wire _11268_ ;
wire _9836_ ;
wire _9416_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _7902_ ;
wire _10959_ ;
wire _10539_ ;
wire _10119_ ;
wire _587_ ;
wire _167_ ;
wire _11900_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _10292_ ;
wire _4607_ ;
wire _7499_ ;
wire _7079_ ;
wire _8860_ ;
wire _8440_ ;
wire _8020_ ;
wire _11497_ ;
wire _11077_ ;
wire _9645_ ;
wire _9225_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _2519__bF$buf0 ;
wire _2519__bF$buf1 ;
wire _2519__bF$buf2 ;
wire _2519__bF$buf3 ;
wire _1485_ ;
wire _1065_ ;
wire _7711_ ;
wire _10768_ ;
wire _10348_ ;
wire _396_ ;
wire _8916_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _9874_ ;
wire _9454_ ;
wire _9034_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _7940_ ;
wire _7520_ ;
wire _7100_ ;
wire _10997_ ;
wire _10577_ ;
wire _10157_ ;
wire _2499_ ;
wire _2079_ ;
wire _8725_ ;
wire _8305_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _9683_ ;
wire _9263_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire _10386_ ;
wire _8954_ ;
wire _8534_ ;
wire _8114_ ;
wire _9739_ ;
wire _9319_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _9492_ ;
wire _9072_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _7805_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _11803_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _10195_ ;
wire _8763_ ;
wire _8343_ ;
wire _9968_ ;
wire _9548_ ;
wire _9128_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _5921__bF$buf0 ;
wire _5921__bF$buf1 ;
wire _5921__bF$buf2 ;
wire _5921__bF$buf3 ;
wire _1388_ ;
wire _7614_ ;
wire _299_ ;
wire _11612_ ;
wire _8819_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _8992_ ;
wire _8572_ ;
wire _8152_ ;
wire areg_18_bF$buf0 ;
wire areg_18_bF$buf1 ;
wire areg_18_bF$buf2 ;
wire areg_18_bF$buf3 ;
wire areg_18_bF$buf4 ;
wire areg_18_bF$buf5 ;
wire _18_ ;
wire _1600_ ;
wire _9777_ ;
wire _9357_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7843_ ;
wire _7423_ ;
wire _7003_ ;
wire _11841_ ;
wire _11421_ ;
wire _11001_ ;
wire _8628_ ;
wire _8208_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _8381_ ;
wire _9586_ ;
wire _9166_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _7652_ ;
wire _7232_ ;
wire _10289_ ;
wire _11650_ ;
wire _11230_ ;
wire _8857_ ;
wire _8437_ ;
wire _8017_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _8190_ ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire _9395_ ;
wire _10921_ ;
wire _10501_ ;
wire _7708_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _11706_ ;
wire _3628_ ;
wire _3208_ ;
wire _7881_ ;
wire _7461_ ;
wire _7041_ ;
wire _10098_ ;
wire _8666_ ;
wire _8246_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _10730_ ;
wire _10310_ ;
wire _7937_ ;
wire _7517_ ;
wire _2652_ ;
wire _2232_ ;
wire _11515_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _7690_ ;
wire _7270_ ;
wire _8895_ ;
wire _8475_ ;
wire _8055_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _7746_ ;
wire _7326_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _11744_ ;
wire _11324_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _8284_ ;
wire _1732_ ;
wire _1312_ ;
wire _9489_ ;
wire _9069_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire _7975_ ;
wire _7555_ ;
wire _7135_ ;
wire _2690_ ;
wire _2270_ ;
wire _11553_ ;
wire _11133_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _9701_ ;
wire _5621_ ;
wire _5201_ ;
wire _8093_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _9298_ ;
wire _10824_ ;
wire _10404_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _11609_ ;
wire _7784_ ;
wire _7364_ ;
wire _11782_ ;
wire _11362_ ;
wire _8989_ ;
wire _8569_ ;
wire _8149_ ;
wire _3284_ ;
wire _9930_ ;
wire _9510_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _10633_ ;
wire _10213_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _11838_ ;
wire _11418_ ;
wire _4701_ ;
wire _7593_ ;
wire _7173_ ;
wire _11591_ ;
wire _11171_ ;
wire _5906_ ;
wire _8798_ ;
wire _8378_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _10862_ ;
wire _10442_ ;
wire _10022_ ;
wire _490_ ;
wire _7649_ ;
wire _7229_ ;
wire _2784_ ;
wire _2364_ ;
wire _11647_ ;
wire _11227_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _8187_ ;
wire _1635_ ;
wire _1215_ ;
wire _10918_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _10671_ ;
wire _10251_ ;
wire _7878_ ;
wire _7458_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _11876_ ;
wire _11456_ ;
wire _11036_ ;
wire _3798_ ;
wire _3378_ ;
wire _9604_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _10727_ ;
wire _10307_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _10480_ ;
wire _10060_ ;
wire _7687_ ;
wire _7267_ ;
wire _11685_ ;
wire _11265_ ;
wire _3187_ ;
wire _9833_ ;
wire _9413_ ;
wire _5753_ ;
wire _5333_ ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _10956_ ;
wire _10536_ ;
wire _10116_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _7496_ ;
wire _7076_ ;
wire _11494_ ;
wire _11074_ ;
wire _5809_ ;
wire _9642_ ;
wire _9222_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _10765_ ;
wire _10345_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _8913_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _9871_ ;
wire _9451_ ;
wire _9031_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _10994_ ;
wire _10574_ ;
wire _10154_ ;
wire _2496_ ;
wire _2076_ ;
wire _8722_ ;
wire _8302_ ;
wire _11779_ ;
wire _11359_ ;
wire _9927_ ;
wire _9507_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _9680_ ;
wire _9260_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _10383_ ;
wire _8951_ ;
wire _8531_ ;
wire _8111_ ;
wire _11588_ ;
wire _11168_ ;
wire _9736_ ;
wire _9316_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _7802_ ;
wire _10859_ ;
wire _10439_ ;
wire _10019_ ;
wire _487_ ;
wire _11800_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire breg_11_bF$buf0 ;
wire breg_11_bF$buf1 ;
wire breg_11_bF$buf2 ;
wire breg_11_bF$buf3 ;
wire _10192_ ;
wire breg_11_bF$buf4 ;
wire _4927_ ;
wire _4507_ ;
wire _7399_ ;
wire _8760_ ;
wire _8340_ ;
wire _11397_ ;
wire _9965_ ;
wire _9545_ ;
wire _9125_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _7611_ ;
wire _10668_ ;
wire _10248_ ;
wire _296_ ;
wire _8816_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _9774_ ;
wire _9354_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7840_ ;
wire _7420_ ;
wire _7000_ ;
wire _10897_ ;
wire _10477_ ;
wire _10057_ ;
wire _2399_ ;
wire _8625_ ;
wire _8205_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _9583_ ;
wire _9163_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _10286_ ;
wire _8854_ ;
wire _8434_ ;
wire _8014_ ;
wire _9639_ ;
wire _9219_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _9392_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _7705_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _11703_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _10095_ ;
wire _8663_ ;
wire _8243_ ;
wire _9868_ ;
wire _9448_ ;
wire _9028_ ;
wire _4583_ ;
wire _4163_ ;
wire areg_29_bF$buf0 ;
wire areg_29_bF$buf1 ;
wire areg_29_bF$buf2 ;
wire areg_29_bF$buf3 ;
wire areg_29_bF$buf4 ;
wire areg_29_bF$buf5 ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire [31:0] breg ;
wire _1288_ ;
wire _7934_ ;
wire _7514_ ;
wire _199_ ;
wire _11512_ ;
wire _8719_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _8892_ ;
wire _8472_ ;
wire _8052_ ;
wire _1920_ ;
wire _1500_ ;
wire _9677_ ;
wire _9257_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _6300__bF$buf0 ;
wire _6300__bF$buf1 ;
wire _6300__bF$buf2 ;
wire _6300__bF$buf3 ;
wire _5597_ ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _7743_ ;
wire _7323_ ;
wire _11741_ ;
wire _11321_ ;
wire _8948_ ;
wire _8528_ ;
wire _8108_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _8281_ ;
wire _9486_ ;
wire _9066_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _7972_ ;
wire _7552_ ;
wire _7132_ ;
wire _10189_ ;
wire _11550_ ;
wire _11130_ ;
wire _8757_ ;
wire _8337_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _8090_ ;
wire _6823_ ;
wire _6403_ ;
wire _9295_ ;
wire _10821_ ;
wire _10401_ ;
wire _7608_ ;
wire _2743_ ;
wire _2323_ ;
wire _11606_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _7781_ ;
wire _7361_ ;
wire _8986_ ;
wire _8566_ ;
wire _8146_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _10630_ ;
wire _10210_ ;
wire _7837_ ;
wire _7417_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _11835_ ;
wire _11415_ ;
wire _3757_ ;
wire _3337_ ;
wire _7590_ ;
wire _7170_ ;
wire _5903_ ;
wire _8795_ ;
wire _8375_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire _7646_ ;
wire _7226_ ;
wire _2781_ ;
wire _2361_ ;
wire _11644_ ;
wire _11224_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _8184_ ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _9389_ ;
wire _10915_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7875_ ;
wire _7455_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _11873_ ;
wire _11453_ ;
wire _11033_ ;
wire _3795_ ;
wire _3375_ ;
wire _9601_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _9198_ ;
wire _10724_ ;
wire _10304_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire areg_13_bF$buf0 ;
wire areg_13_bF$buf1 ;
wire _11509_ ;
wire areg_13_bF$buf2 ;
wire areg_13_bF$buf3 ;
wire areg_13_bF$buf4 ;
wire _7684_ ;
wire _7264_ ;
wire _11682_ ;
wire _11262_ ;
wire _8889_ ;
wire _8469_ ;
wire _8049_ ;
wire _3184_ ;
wire _9830_ ;
wire _9410_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _2825__bF$buf0 ;
wire _6955_ ;
wire _2825__bF$buf1 ;
wire _6535_ ;
wire _2825__bF$buf2 ;
wire _6115_ ;
wire _2825__bF$buf3 ;
wire _2825__bF$buf4 ;
wire _1670_ ;
wire _1250_ ;
wire _10953_ ;
wire _10533_ ;
wire _10113_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _11738_ ;
wire _11318_ ;
wire _4601_ ;
wire _7493_ ;
wire _7073_ ;
wire _11491_ ;
wire _11071_ ;
wire _5806_ ;
wire _8698_ ;
wire _8278_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6764_ ;
wire _6344_ ;
wire _10762_ ;
wire _10342_ ;
wire _390_ ;
wire _7969_ ;
wire _7549_ ;
wire _7129_ ;
wire _2684_ ;
wire _2264_ ;
wire _8910_ ;
wire _11547_ ;
wire _11127_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _8087_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _10818_ ;
wire _866_ ;
wire _446_ ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _10991_ ;
wire _10571_ ;
wire _10151_ ;
wire _7778_ ;
wire _7358_ ;
wire _2493_ ;
wire _2073_ ;
wire _11776_ ;
wire _11356_ ;
wire _3698_ ;
wire _3278_ ;
wire _9924_ ;
wire _9504_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _3961__bF$buf0 ;
wire _3961__bF$buf1 ;
wire _3961__bF$buf2 ;
wire _3961__bF$buf3 ;
wire _3961__bF$buf4 ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _10627_ ;
wire _10207_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _10380_ ;
wire _7587_ ;
wire _7167_ ;
wire _11585_ ;
wire _11165_ ;
wire _3087_ ;
wire _3646__bF$buf0 ;
wire _3646__bF$buf1 ;
wire _3646__bF$buf2 ;
wire _9733_ ;
wire _3646__bF$buf3 ;
wire _9313_ ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _10856_ ;
wire _10436_ ;
wire _10016_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _7396_ ;
wire _11394_ ;
wire _5709_ ;
wire _9962_ ;
wire _9542_ ;
wire _9122_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _10665_ ;
wire _10245_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _8813_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _9771_ ;
wire _9351_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _10894_ ;
wire _10474_ ;
wire _10054_ ;
wire _2396_ ;
wire _8622_ ;
wire _8202_ ;
wire _11679_ ;
wire _11259_ ;
wire _9827_ ;
wire _9407_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _9580_ ;
wire _9160_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _10283_ ;
wire _8851_ ;
wire _8431_ ;
wire _8011_ ;
wire _11488_ ;
wire _11068_ ;
wire _9636_ ;
wire _9216_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _7702_ ;
wire _10759_ ;
wire _10339_ ;
wire _387_ ;
wire _11700_ ;
wire _8907_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire breg_9_bF$buf0 ;
wire breg_9_bF$buf1 ;
wire _10092_ ;
wire breg_9_bF$buf2 ;
wire breg_9_bF$buf3 ;
wire breg_9_bF$buf4 ;
wire _4827_ ;
wire breg_9_bF$buf5 ;
wire _4407_ ;
wire _7299_ ;
wire _8660_ ;
wire _8240_ ;
wire _11297_ ;
wire _9865_ ;
wire _9445_ ;
wire _9025_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _7931_ ;
wire _7511_ ;
wire _10988_ ;
wire _10568_ ;
wire _10148_ ;
wire _196_ ;
wire _8716_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _9674_ ;
wire _9254_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _7740_ ;
wire _7320_ ;
wire _10797_ ;
wire _10377_ ;
wire _2299_ ;
wire _8945_ ;
wire _8525_ ;
wire _8105_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _9483_ ;
wire _9063_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire _10186_ ;
wire _8754_ ;
wire _8334_ ;
wire _9959_ ;
wire _9539_ ;
wire _9119_ ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _9292_ ;
wire _1799_ ;
wire _1379_ ;
wire _7605_ ;
wire _2740_ ;
wire _2320_ ;
wire _11603_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _8983_ ;
wire _8563_ ;
wire _8143_ ;
wire _9768_ ;
wire _9348_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire [31:0] areg ;
wire _1188_ ;
wire _7834_ ;
wire _7414_ ;
wire _11832_ ;
wire _11412_ ;
wire _8619_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _8792_ ;
wire _8372_ ;
wire _1820_ ;
wire _1400_ ;
wire _9997_ ;
wire _9577_ ;
wire _9157_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _7643_ ;
wire _7223_ ;
wire _11641_ ;
wire _11221_ ;
wire _8848_ ;
wire _8428_ ;
wire _8008_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _8181_ ;
wire _47_ ;
wire _6914_ ;
wire _9386_ ;
wire _10912_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire _7872_ ;
wire _7452_ ;
wire _7032_ ;
wire _10089_ ;
wire _11870_ ;
wire _11450_ ;
wire _11030_ ;
wire _8657_ ;
wire _8237_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _9195_ ;
wire _10721_ ;
wire _10301_ ;
wire _7928_ ;
wire _7508_ ;
wire _2643_ ;
wire _2223_ ;
wire _11506_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _7681_ ;
wire _7261_ ;
wire _8886_ ;
wire _8466_ ;
wire _8046_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _10950_ ;
wire _10530_ ;
wire _10110_ ;
wire _7737_ ;
wire _7317_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _11735_ ;
wire _11315_ ;
wire _3657_ ;
wire _3237_ ;
wire _7490_ ;
wire _7070_ ;
wire _5803_ ;
wire _8695_ ;
wire _8275_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _7966_ ;
wire _7546_ ;
wire _7126_ ;
wire _2681_ ;
wire _2261_ ;
wire _11544_ ;
wire _11124_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _8084_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _9289_ ;
wire _10815_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _7775_ ;
wire _7355_ ;
wire areg_24_bF$buf0 ;
wire areg_24_bF$buf1 ;
wire areg_24_bF$buf2 ;
wire areg_24_bF$buf3 ;
wire _2490_ ;
wire areg_24_bF$buf4 ;
wire _2070_ ;
wire _11773_ ;
wire _11353_ ;
wire _3695_ ;
wire _3275_ ;
wire _9921_ ;
wire _9501_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _9098_ ;
wire _10624_ ;
wire _10204_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _11829_ ;
wire _11409_ ;
wire _7584_ ;
wire _7164_ ;
wire _11582_ ;
wire _11162_ ;
wire _8789_ ;
wire _8369_ ;
wire _3084_ ;
wire _9730_ ;
wire _9310_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _10853_ ;
wire _10433_ ;
wire _10013_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _11638_ ;
wire _11218_ ;
wire _4921_ ;
wire _4501_ ;
wire _7393_ ;
wire _11391_ ;
wire _5706_ ;
wire _8598_ ;
wire _8178_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _10909_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6815__bF$buf0 ;
wire _6815__bF$buf1 ;
wire _6815__bF$buf2 ;
wire _6815__bF$buf3 ;
wire _6815__bF$buf4 ;
wire _6664_ ;
wire _6244_ ;
wire _10662_ ;
wire _10242_ ;
wire _290_ ;
wire _7869_ ;
wire _7449_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _8810_ ;
wire _11867_ ;
wire _11447_ ;
wire _11027_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _10718_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _10891_ ;
wire _10471_ ;
wire _10051_ ;
wire _7678_ ;
wire _7258_ ;
wire _2393_ ;
wire _11676_ ;
wire _11256_ ;
wire _3598_ ;
wire _3178_ ;
wire _9824_ ;
wire _9404_ ;
wire areg_6_bF$buf0 ;
wire areg_6_bF$buf1 ;
wire areg_6_bF$buf2 ;
wire areg_6_bF$buf3 ;
wire areg_6_bF$buf4 ;
wire _5744_ ;
wire _5324_ ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _10947_ ;
wire _10527_ ;
wire _10107_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _10280_ ;
wire _7487_ ;
wire _7067_ ;
wire _11485_ ;
wire _11065_ ;
wire _9633_ ;
wire _9213_ ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _10756_ ;
wire _10336_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _8904_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _7296_ ;
wire _11294_ ;
wire _5609_ ;
wire _9862_ ;
wire _9442_ ;
wire _9022_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _10985_ ;
wire _10565_ ;
wire _10145_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _8713_ ;
wire _9918_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _9671_ ;
wire _9251_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _10794_ ;
wire _10374_ ;
wire _2296_ ;
wire _8942_ ;
wire _8522_ ;
wire _8102_ ;
wire _11579_ ;
wire _11159_ ;
wire _9727_ ;
wire _9307_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _9480_ ;
wire _9060_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _10183_ ;
wire _4918_ ;
wire _8751_ ;
wire _8331_ ;
wire _11388_ ;
wire _9956_ ;
wire _9536_ ;
wire _9116_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _7602_ ;
wire _10659_ ;
wire _10239_ ;
wire _287_ ;
wire _11600_ ;
wire _8807_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _7199_ ;
wire _8980_ ;
wire _8560_ ;
wire _8140_ ;
wire _11197_ ;
wire _9765_ ;
wire _9345_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _7831_ ;
wire _7411_ ;
wire _10888_ ;
wire _10468_ ;
wire _10048_ ;
wire _8616_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _9994_ ;
wire _9574_ ;
wire _9154_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _7640_ ;
wire _7220_ ;
wire _10697_ ;
wire _10277_ ;
wire _2199_ ;
wire _8845_ ;
wire _8425_ ;
wire _8005_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _6911_ ;
wire _9383_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _10086_ ;
wire _8654_ ;
wire _8234_ ;
wire _9859_ ;
wire _9439_ ;
wire _9019_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _9192_ ;
wire _1699_ ;
wire _1279_ ;
wire _7925_ ;
wire _7505_ ;
wire _2640_ ;
wire _2220_ ;
wire _11503_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _8883_ ;
wire _8463_ ;
wire _8043_ ;
wire _1911_ ;
wire _9668_ ;
wire _9248_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _7734_ ;
wire _7314_ ;
wire _11732_ ;
wire _11312_ ;
wire _8939_ ;
wire _8519_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _8692_ ;
wire _8272_ ;
wire _1720_ ;
wire _1300_ ;
wire _9897_ ;
wire _9477_ ;
wire _9057_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _7963_ ;
wire _7543_ ;
wire _7123_ ;
wire breg_26_bF$buf0 ;
wire breg_26_bF$buf1 ;
wire breg_26_bF$buf2 ;
wire breg_26_bF$buf3 ;
wire breg_26_bF$buf4 ;
wire _4541__bF$buf0 ;
wire _4541__bF$buf1 ;
wire _4541__bF$buf2 ;
wire _4541__bF$buf3 ;
wire _4541__bF$buf4 ;
wire _11541_ ;
wire _11121_ ;
wire _8748_ ;
wire _8328_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _8081_ ;
wire _6814_ ;
wire _9286_ ;
wire breg_4_bF$buf0 ;
wire breg_4_bF$buf1 ;
wire breg_4_bF$buf2 ;
wire _10812_ ;
wire breg_4_bF$buf3 ;
wire breg_4_bF$buf4 ;
wire breg_4_bF$buf5 ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _7772_ ;
wire _7352_ ;
wire _11770_ ;
wire _11350_ ;
wire _8977_ ;
wire _8557_ ;
wire _8137_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _9095_ ;
wire _10621_ ;
wire _10201_ ;
wire _7828_ ;
wire _7408_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _11826_ ;
wire _11406_ ;
wire _3748_ ;
wire _3328_ ;
wire _7581_ ;
wire _7161_ ;
wire _8786_ ;
wire _8366_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire _10850_ ;
wire _10430_ ;
wire _10010_ ;
wire _7637_ ;
wire _7217_ ;
wire _2772_ ;
wire _2352_ ;
wire _11635_ ;
wire _11215_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _7390_ ;
wire _5703_ ;
wire _8595_ ;
wire _8175_ ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _10906_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7866_ ;
wire _7446_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _11864_ ;
wire _11444_ ;
wire _11024_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _9189_ ;
wire _10715_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire _7675_ ;
wire _7255_ ;
wire _2390_ ;
wire _11673_ ;
wire _11253_ ;
wire _3595_ ;
wire _3175_ ;
wire _9821_ ;
wire _9401_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _10944_ ;
wire _10524_ ;
wire _10104_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _11729_ ;
wire _11309_ ;
wire _7484_ ;
wire _7064_ ;
wire _11482_ ;
wire _11062_ ;
wire _8689_ ;
wire _8269_ ;
wire _9630_ ;
wire _9210_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _10753_ ;
wire _10333_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _8901_ ;
wire _11538_ ;
wire _11118_ ;
wire _4821_ ;
wire _4401_ ;
wire _7293_ ;
wire _11291_ ;
wire _5606_ ;
wire _8498_ ;
wire _8078_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _10809_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire _10982_ ;
wire _10562_ ;
wire _10142_ ;
wire _190_ ;
wire _7769_ ;
wire _7349_ ;
wire _2484_ ;
wire _2064_ ;
wire _8710_ ;
wire _11767_ ;
wire _11347_ ;
wire _3689_ ;
wire _3269_ ;
wire _9915_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _10618_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _10791_ ;
wire _10371_ ;
wire _7998_ ;
wire _7578_ ;
wire _7158_ ;
wire _2293_ ;
wire _11576_ ;
wire _11156_ ;
wire _3498_ ;
wire _3078_ ;
wire _9724_ ;
wire _9304_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _10847_ ;
wire _10427_ ;
wire _10007_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _10180_ ;
wire _4915_ ;
wire _7387_ ;
wire _11385_ ;
wire _9953_ ;
wire _9533_ ;
wire _9113_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _10656_ ;
wire _10236_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _8804_ ;
wire [63:0] _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _7196_ ;
wire _11194_ ;
wire _5929_ ;
wire _5509_ ;
wire _9762_ ;
wire _9342_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _10885_ ;
wire _10465_ ;
wire _10045_ ;
wire _2387_ ;
wire _8613_ ;
wire _9818_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _9991_ ;
wire _9571_ ;
wire _9151_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _10694_ ;
wire _10274_ ;
wire _2196_ ;
wire _8842_ ;
wire _8422_ ;
wire _8002_ ;
wire _11899_ ;
wire _11479_ ;
wire _11059_ ;
wire _9627_ ;
wire _9207_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _9380_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _10083_ ;
wire _4818_ ;
wire _8651_ ;
wire _8231_ ;
wire _11288_ ;
wire _9856_ ;
wire _9436_ ;
wire _9016_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _7922_ ;
wire _7502_ ;
wire _10979_ ;
wire _10559_ ;
wire _10139_ ;
wire _187_ ;
wire _11500_ ;
wire _8707_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _7099_ ;
wire _8880_ ;
wire _8460_ ;
wire _8040_ ;
wire _11097_ ;
wire _9665_ ;
wire _9245_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _7731_ ;
wire _7311_ ;
wire areg_1_bF$buf0 ;
wire areg_1_bF$buf1 ;
wire areg_1_bF$buf2 ;
wire areg_1_bF$buf3 ;
wire areg_1_bF$buf4 ;
wire _10788_ ;
wire _10368_ ;
wire _8936_ ;
wire _8516_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _9894_ ;
wire _9474_ ;
wire _9054_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _7960_ ;
wire _7540_ ;
wire _7120_ ;
wire _10597_ ;
wire _10177_ ;
wire _2099_ ;
wire _8745_ ;
wire _8325_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _9283_ ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire _8974_ ;
wire _8554_ ;
wire _8134_ ;
wire _9759_ ;
wire _9339_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _9092_ ;
wire _1599_ ;
wire _1179_ ;
wire _7825_ ;
wire _7405_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _11823_ ;
wire _11403_ ;
wire _3745_ ;
wire _3325_ ;
wire _8783_ ;
wire _8363_ ;
wire _1811_ ;
wire _9988_ ;
wire _9568_ ;
wire _9148_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _7634_ ;
wire _7214_ ;
wire breg_18_bF$buf0 ;
wire breg_18_bF$buf1 ;
wire breg_18_bF$buf2 ;
wire breg_18_bF$buf3 ;
wire breg_18_bF$buf4 ;
wire breg_18_bF$buf5 ;
wire _11632_ ;
wire _11212_ ;
wire _8839_ ;
wire _8419_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _8592_ ;
wire _8172_ ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _9797_ ;
wire _9377_ ;
wire _4092_ ;
wire _10903_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7863_ ;
wire _7443_ ;
wire _7023_ ;
wire _11861_ ;
wire _11441_ ;
wire _11021_ ;
wire _8648_ ;
wire _8228_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _9186_ ;
wire _10712_ ;
wire _760_ ;
wire _340_ ;
wire _7919_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _7672_ ;
wire _7252_ ;
wire _11670_ ;
wire _11250_ ;
wire _8877_ ;
wire _8457_ ;
wire _8037_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _10941_ ;
wire _10521_ ;
wire _10101_ ;
wire _7728_ ;
wire _7308_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _11726_ ;
wire _11306_ ;
wire _3648_ ;
wire _3228_ ;
wire _7481_ ;
wire _7061_ ;
wire _8686_ ;
wire _8266_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _10750_ ;
wire _10330_ ;
wire _7957_ ;
wire _7537_ ;
wire _2562__bF$buf0 ;
wire _7117_ ;
wire _2562__bF$buf1 ;
wire _2562__bF$buf2 ;
wire _2562__bF$buf3 ;
wire _2672_ ;
wire _2562__bF$buf4 ;
wire _2252_ ;
wire clk_bF$buf10 ;
wire _11535_ ;
wire _11115_ ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _7290_ ;
wire _5603_ ;
wire _8495_ ;
wire _8075_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _10806_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire _7766_ ;
wire _7346_ ;
wire _2481_ ;
wire _2061_ ;
wire _11764_ ;
wire _11344_ ;
wire _3686_ ;
wire _3266_ ;
wire _9912_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _9089_ ;
wire _10615_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _7995_ ;
wire _7575_ ;
wire _7155_ ;
wire _2290_ ;
wire _11573_ ;
wire _11153_ ;
wire _3495_ ;
wire _3075_ ;
wire _9721_ ;
wire _9301_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _10844_ ;
wire _10424_ ;
wire _10004_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _11629_ ;
wire _11209_ ;
wire _4912_ ;
wire _7384_ ;
wire _11382_ ;
wire _8589_ ;
wire _8169_ ;
wire _9950_ ;
wire _9530_ ;
wire _9110_ ;
wire _1617_ ;
wire breg_21_bF$buf0 ;
wire breg_21_bF$buf1 ;
wire breg_21_bF$buf2 ;
wire _4089_ ;
wire breg_21_bF$buf3 ;
wire breg_21_bF$buf4 ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _10653_ ;
wire _10233_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _8801_ ;
wire _11858_ ;
wire _11438_ ;
wire _11018_ ;
wire _4721_ ;
wire _4301_ ;
wire _7193_ ;
wire _11191_ ;
wire _5926_ ;
wire _5506_ ;
wire _8398_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _10709_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire _10882_ ;
wire _10462_ ;
wire _10042_ ;
wire _7669_ ;
wire _7249_ ;
wire _2384_ ;
wire _8610_ ;
wire _11667_ ;
wire _11247_ ;
wire _3589_ ;
wire _3169_ ;
wire _9815_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _10938_ ;
wire _10518_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _10691_ ;
wire _10271_ ;
wire _7898_ ;
wire _7478_ ;
wire _7058_ ;
wire _2193_ ;
wire _11896_ ;
wire _11476_ ;
wire _11056_ ;
wire _3398_ ;
wire _9624_ ;
wire _9204_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _10747_ ;
wire _10327_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _10080_ ;
wire _4815_ ;
wire _7287_ ;
wire _11285_ ;
wire _9853_ ;
wire _9433_ ;
wire _9013_ ;
wire _5773_ ;
wire _5353_ ;
wire areg_30_bF$buf0 ;
wire areg_30_bF$buf1 ;
wire areg_30_bF$buf2 ;
wire areg_30_bF$buf3 ;
wire areg_30_bF$buf4 ;
wire areg_30_bF$buf5 ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _10976_ ;
wire _10556_ ;
wire _10136_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _8704_ ;
wire _9909_ ;
wire _4624_ ;
wire _4204_ ;
wire _7096_ ;
wire _11094_ ;
wire _5829_ ;
wire _5409_ ;
wire _9662_ ;
wire _9242_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _10785_ ;
wire _10365_ ;
wire _2287_ ;
wire _8933_ ;
wire _8513_ ;
wire _9718_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _9891_ ;
wire _9471_ ;
wire _9051_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _10594_ ;
wire _10174_ ;
wire _4909_ ;
wire _2096_ ;
wire _8742_ ;
wire _8322_ ;
wire _11799_ ;
wire _11379_ ;
wire _9947_ ;
wire _9527_ ;
wire _9107_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _9280_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _8971_ ;
wire _8551_ ;
wire _8131_ ;
wire _11188_ ;
wire _9756_ ;
wire _9336_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _7822_ ;
wire _7402_ ;
wire _10879_ ;
wire _10459_ ;
wire _10039_ ;
wire _11820_ ;
wire _11400_ ;
wire _8607_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _8780_ ;
wire _8360_ ;
wire _9985_ ;
wire _9565_ ;
wire _9145_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _7631_ ;
wire _7211_ ;
wire _10688_ ;
wire _10268_ ;
wire _8836_ ;
wire _8416_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _6902_ ;
wire _9794_ ;
wire _9374_ ;
wire _10900_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7860_ ;
wire _7440_ ;
wire _7020_ ;
wire _10497_ ;
wire _10077_ ;
wire _8645_ ;
wire _8225_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _9183_ ;
wire _7916_ ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _8874_ ;
wire _8454_ ;
wire _8034_ ;
wire _1902_ ;
wire _9659_ ;
wire _9239_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _7725_ ;
wire _7305_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _11723_ ;
wire _11303_ ;
wire _3645_ ;
wire _3225_ ;
wire _8683_ ;
wire _8263_ ;
wire _1711_ ;
wire _9888_ ;
wire _9468_ ;
wire _9048_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _7954_ ;
wire _7534_ ;
wire _7114_ ;
wire _11532_ ;
wire _11112_ ;
wire _8739_ ;
wire _8319_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _8492_ ;
wire _8072_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _9697_ ;
wire _9277_ ;
wire _10803_ ;
wire _4551__bF$buf0 ;
wire _4551__bF$buf1 ;
wire _4551__bF$buf2 ;
wire _4551__bF$buf3 ;
wire _4551__bF$buf4 ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3958__bF$buf0 ;
wire _3958__bF$buf1 ;
wire _3958__bF$buf2 ;
wire _7763_ ;
wire _3958__bF$buf3 ;
wire _7343_ ;
wire _11761_ ;
wire _11341_ ;
wire _8968_ ;
wire _8548_ ;
wire _8128_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _9086_ ;
wire _10612_ ;
wire _660_ ;
wire _240_ ;
wire _7819_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _11817_ ;
wire _3739_ ;
wire _3319_ ;
wire _7992_ ;
wire _7572_ ;
wire _7152_ ;
wire _11570_ ;
wire _11150_ ;
wire _8777_ ;
wire _8357_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _10841_ ;
wire _10421_ ;
wire _10001_ ;
wire _7628_ ;
wire _7208_ ;
wire _2763_ ;
wire _2343_ ;
wire _11626_ ;
wire _11206_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _7381_ ;
wire _8586_ ;
wire _8166_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _10650_ ;
wire _10230_ ;
wire _7857_ ;
wire _7437_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _11855_ ;
wire _11435_ ;
wire _11015_ ;
wire _3777_ ;
wire _3357_ ;
wire _7190_ ;
wire _5923_ ;
wire _5503_ ;
wire _8395_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _10706_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire _7666_ ;
wire _7246_ ;
wire _2381_ ;
wire _11664_ ;
wire _11244_ ;
wire _3586_ ;
wire _3166_ ;
wire _9812_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _10935_ ;
wire _10515_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _7895_ ;
wire _7475_ ;
wire _7055_ ;
wire _2190_ ;
wire _11893_ ;
wire _11473_ ;
wire _11053_ ;
wire _3395_ ;
wire _9621_ ;
wire _9201_ ;
wire _1708_ ;
wire breg_13_bF$buf0 ;
wire breg_13_bF$buf1 ;
wire breg_13_bF$buf2 ;
wire breg_13_bF$buf3 ;
wire breg_13_bF$buf4 ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _10744_ ;
wire _10324_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _11529_ ;
wire _11109_ ;
wire _4812_ ;
wire _7284_ ;
wire _11282_ ;
wire _8489_ ;
wire _8069_ ;
wire _9850_ ;
wire _9430_ ;
wire _9010_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _10973_ ;
wire _10553_ ;
wire _10133_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _8701_ ;
wire _11758_ ;
wire _11338_ ;
wire _9906_ ;
wire _4621_ ;
wire _4201_ ;
wire _7093_ ;
wire _11091_ ;
wire _5826_ ;
wire _5406_ ;
wire _8298_ ;
wire _1746_ ;
wire _1326_ ;
wire _10609_ ;
wire _657_ ;
wire _237_ ;
wire _6686__bF$buf0 ;
wire _6686__bF$buf1 ;
wire _6686__bF$buf2 ;
wire _6686__bF$buf3 ;
wire _6784_ ;
wire _6364_ ;
wire _10782_ ;
wire _10362_ ;
wire _7989_ ;
wire _7569_ ;
wire _7149_ ;
wire _2284_ ;
wire _8930_ ;
wire _8510_ ;
wire _11567_ ;
wire _11147_ ;
wire _3489_ ;
wire _3069_ ;
wire _9715_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _10838_ ;
wire _10418_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _10591_ ;
wire _10171_ ;
wire _4906_ ;
wire _7798_ ;
wire _7378_ ;
wire _2093_ ;
wire _11796_ ;
wire _11376_ ;
wire _3298_ ;
wire _9944_ ;
wire _9524_ ;
wire _9104_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _10647_ ;
wire _10227_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _7187_ ;
wire _11185_ ;
wire _9753_ ;
wire _9333_ ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _10876_ ;
wire _10456_ ;
wire _10036_ ;
wire _2798_ ;
wire _2378_ ;
wire _8604_ ;
wire _9809_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _9982_ ;
wire _9562_ ;
wire _9142_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _10685_ ;
wire _10265_ ;
wire _2187_ ;
wire _8833_ ;
wire _8413_ ;
wire _9618_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _9791_ ;
wire _9371_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _10494_ ;
wire _10074_ ;
wire _4809_ ;
wire _8642_ ;
wire _8222_ ;
wire _11699_ ;
wire _11279_ ;
wire _9847_ ;
wire _9427_ ;
wire _9007_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _9180_ ;
wire _1687_ ;
wire _1267_ ;
wire _7913_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _8871_ ;
wire _8451_ ;
wire _8031_ ;
wire _11088_ ;
wire _9656_ ;
wire _9236_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _7722_ ;
wire _7302_ ;
wire _10779_ ;
wire _10359_ ;
wire _11720_ ;
wire _11300_ ;
wire _8927_ ;
wire _8507_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _8680_ ;
wire _8260_ ;
wire _9885_ ;
wire _9465_ ;
wire _9045_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _7951_ ;
wire _7531_ ;
wire _7111_ ;
wire _10588_ ;
wire _10168_ ;
wire _8736_ ;
wire _8316_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _9694_ ;
wire _9274_ ;
wire _10800_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _7760_ ;
wire _7340_ ;
wire _10397_ ;
wire _8965_ ;
wire _8545_ ;
wire _8125_ ;
wire _3680_ ;
wire _3260_ ;
wire areg_15_bF$buf0 ;
wire areg_15_bF$buf1 ;
wire areg_15_bF$buf2 ;
wire areg_15_bF$buf3 ;
wire areg_15_bF$buf4 ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _9083_ ;
wire _7816_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _11814_ ;
wire _3736_ ;
wire _3316_ ;
wire _8774_ ;
wire _8354_ ;
wire _1802_ ;
wire _9979_ ;
wire _9559_ ;
wire _9139_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _7625_ ;
wire _7205_ ;
wire _2760_ ;
wire _2340_ ;
wire _11623_ ;
wire _11203_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _8583_ ;
wire _8163_ ;
wire _29_ ;
wire _1611_ ;
wire _9788_ ;
wire _9368_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7854_ ;
wire _7434_ ;
wire _7014_ ;
wire _11852_ ;
wire _11432_ ;
wire _11012_ ;
wire _8639_ ;
wire _8219_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _8392_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _9597_ ;
wire _9177_ ;
wire _10703_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire _11908_ ;
wire _7663_ ;
wire _7243_ ;
wire _11661_ ;
wire _11241_ ;
wire _8868_ ;
wire _8448_ ;
wire _8028_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _10932_ ;
wire _10512_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _7719_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _11717_ ;
wire _3639_ ;
wire _3219_ ;
wire _7892_ ;
wire _7472_ ;
wire _7052_ ;
wire _11890_ ;
wire _11470_ ;
wire _11050_ ;
wire _8677_ ;
wire _8257_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _10741_ ;
wire _10321_ ;
wire _7948_ ;
wire _7528_ ;
wire _7108_ ;
wire _2663_ ;
wire _2243_ ;
wire _11526_ ;
wire _11106_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _7281_ ;
wire _8486_ ;
wire _8066_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _10970_ ;
wire _10550_ ;
wire _10130_ ;
wire _7757_ ;
wire _7337_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _11755_ ;
wire _11335_ ;
wire _3677_ ;
wire _3257_ ;
wire _9903_ ;
wire _7090_ ;
wire _5823_ ;
wire _5403_ ;
wire _8295_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _10606_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _7986_ ;
wire _7566_ ;
wire _7146_ ;
wire _2281_ ;
wire _11564_ ;
wire _11144_ ;
wire _3486_ ;
wire _3066_ ;
wire _9712_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _10835_ ;
wire _10415_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _7795_ ;
wire _7375_ ;
wire _2090_ ;
wire _11793_ ;
wire _11373_ ;
wire _3295_ ;
wire _9941_ ;
wire _9521_ ;
wire _9101_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _10644_ ;
wire _10224_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _11849_ ;
wire _11429_ ;
wire _11009_ ;
wire _4712_ ;
wire _7184_ ;
wire _11182_ ;
wire _5917_ ;
wire _8389_ ;
wire _9750_ ;
wire _9330_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire _10873_ ;
wire _10453_ ;
wire _10033_ ;
wire _2795_ ;
wire _2375_ ;
wire _8601_ ;
wire _11658_ ;
wire _11238_ ;
wire _9806_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _8198_ ;
wire _1646_ ;
wire _1226_ ;
wire _4258__bF$buf0 ;
wire _4258__bF$buf1 ;
wire _4258__bF$buf2 ;
wire _4258__bF$buf3 ;
wire _10929_ ;
wire _10509_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _10682_ ;
wire _10262_ ;
wire _7889_ ;
wire _7469_ ;
wire _7049_ ;
wire _2184_ ;
wire _8830_ ;
wire _8410_ ;
wire _11887_ ;
wire _11467_ ;
wire _11047_ ;
wire _3389_ ;
wire _9615_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _10738_ ;
wire _10318_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _10491_ ;
wire _10071_ ;
wire _4806_ ;
wire _7698_ ;
wire _7278_ ;
wire _11696_ ;
wire _11276_ ;
wire _3198_ ;
wire _9844_ ;
wire _9424_ ;
wire _9004_ ;
wire _5764_ ;
wire _5344_ ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _7910_ ;
wire _10967_ ;
wire _10547_ ;
wire _10127_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _7087_ ;
wire _11085_ ;
wire _9653_ ;
wire _9233_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _10776_ ;
wire _10356_ ;
wire _2698_ ;
wire _2278_ ;
wire _8924_ ;
wire _8504_ ;
wire _9709_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _9882_ ;
wire _9462_ ;
wire _9042_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _10585_ ;
wire _10165_ ;
wire _2087_ ;
wire _8733_ ;
wire _8313_ ;
wire _9938_ ;
wire _9518_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _9691_ ;
wire _9271_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _10394_ ;
wire _4709_ ;
wire _8962_ ;
wire _8542_ ;
wire _8122_ ;
wire _11599_ ;
wire _11179_ ;
wire _9747_ ;
wire _9327_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _9080_ ;
wire _1587_ ;
wire _1167_ ;
wire _7813_ ;
wire _498_ ;
wire _11811_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _8771_ ;
wire _8351_ ;
wire _9976_ ;
wire _9556_ ;
wire _9136_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _7622_ ;
wire _7202_ ;
wire _10679_ ;
wire _10259_ ;
wire _11620_ ;
wire _11200_ ;
wire _8827_ ;
wire _8407_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _8580_ ;
wire _8160_ ;
wire _26_ ;
wire _9785_ ;
wire _9365_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _6050__bF$buf0 ;
wire _6050__bF$buf1 ;
wire _6050__bF$buf2 ;
wire _6050__bF$buf3 ;
wire _7851_ ;
wire _7431_ ;
wire _7011_ ;
wire _10488_ ;
wire _10068_ ;
wire _8636_ ;
wire _8216_ ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire areg_26_bF$buf0 ;
wire areg_26_bF$buf1 ;
wire areg_26_bF$buf2 ;
wire areg_26_bF$buf3 ;
wire areg_26_bF$buf4 ;
wire _6702_ ;
wire _9594_ ;
wire _9174_ ;
wire _10700_ ;
wire _7907_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _11905_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _7660_ ;
wire _7240_ ;
wire _10297_ ;
wire _8865_ ;
wire _8445_ ;
wire _8025_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _7716_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _11714_ ;
wire _3636_ ;
wire _3216_ ;
wire _8674_ ;
wire _8254_ ;
wire _1702_ ;
wire _9879_ ;
wire _9459_ ;
wire _9039_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _7945_ ;
wire _7525_ ;
wire _7105_ ;
wire _2660_ ;
wire _2240_ ;
wire _11523_ ;
wire _11103_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _8483_ ;
wire _8063_ ;
wire _1931_ ;
wire _1511_ ;
wire _9688_ ;
wire _9268_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _7754_ ;
wire _7334_ ;
wire _11752_ ;
wire _11332_ ;
wire _8959_ ;
wire _8539_ ;
wire _8119_ ;
wire _3674_ ;
wire _3254_ ;
wire _9900_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _8292_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _9497_ ;
wire _9077_ ;
wire _10603_ ;
wire _651_ ;
wire _231_ ;
wire areg_8_bF$buf0 ;
wire _2945_ ;
wire areg_8_bF$buf1 ;
wire _2525_ ;
wire areg_8_bF$buf2 ;
wire _2105_ ;
wire areg_8_bF$buf3 ;
wire areg_8_bF$buf4 ;
wire _11808_ ;
wire _7983_ ;
wire _7563_ ;
wire _7143_ ;
wire _11561_ ;
wire _11141_ ;
wire _8768_ ;
wire _8348_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _10832_ ;
wire _10412_ ;
wire _880_ ;
wire _460_ ;
wire _7619_ ;
wire _2754_ ;
wire _2334_ ;
wire _11617_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _7792_ ;
wire _7372_ ;
wire _11790_ ;
wire _11370_ ;
wire _8997_ ;
wire _8577_ ;
wire _8157_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _10641_ ;
wire _10221_ ;
wire _7848_ ;
wire _7428_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _11846_ ;
wire _11426_ ;
wire _11006_ ;
wire _3768_ ;
wire _3348_ ;
wire _7181_ ;
wire _5914_ ;
wire _8386_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire areg_10_bF$buf0 ;
wire areg_10_bF$buf1 ;
wire areg_10_bF$buf2 ;
wire areg_10_bF$buf3 ;
wire areg_10_bF$buf4 ;
wire _10870_ ;
wire _10450_ ;
wire _10030_ ;
wire _7657_ ;
wire _7237_ ;
wire _2792_ ;
wire _2372_ ;
wire _11655_ ;
wire _11235_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _9803_ ;
wire _5723_ ;
wire _5303_ ;
wire _8195_ ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _10926_ ;
wire _10506_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7886_ ;
wire _7466_ ;
wire _7046_ ;
wire _2181_ ;
wire _11884_ ;
wire _11464_ ;
wire _11044_ ;
wire _3386_ ;
wire _9612_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _10735_ ;
wire _10315_ ;
wire _783_ ;
wire _363_ ;
wire _2362__bF$buf0 ;
wire _2657_ ;
wire _2362__bF$buf1 ;
wire _2237_ ;
wire _2362__bF$buf2 ;
wire _2362__bF$buf3 ;
wire _2362__bF$buf4 ;
wire _2362__bF$buf5 ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _7695_ ;
wire _7275_ ;
wire _11693_ ;
wire _11273_ ;
wire _3195_ ;
wire _9841_ ;
wire _9421_ ;
wire _9001_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _10964_ ;
wire _10544_ ;
wire _10124_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _11749_ ;
wire _11329_ ;
wire _4612_ ;
wire _7084_ ;
wire _11082_ ;
wire _5817_ ;
wire _8289_ ;
wire _9650_ ;
wire _9230_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _10773_ ;
wire _10353_ ;
wire _2695_ ;
wire _2275_ ;
wire _8921_ ;
wire _8501_ ;
wire _11558_ ;
wire _11138_ ;
wire _9706_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _8098_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _10829_ ;
wire _10409_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _10582_ ;
wire _10162_ ;
wire _7789_ ;
wire _7369_ ;
wire _2084_ ;
wire _8730_ ;
wire _8310_ ;
wire _11787_ ;
wire _11367_ ;
wire _3289_ ;
wire _9935_ ;
wire _9515_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _10638_ ;
wire _10218_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _10391_ ;
wire _4706_ ;
wire _7598_ ;
wire _7178_ ;
wire _11596_ ;
wire _11176_ ;
wire _3098_ ;
wire _9744_ ;
wire _9324_ ;
wire _5664_ ;
wire _5244_ ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _7810_ ;
wire _10867_ ;
wire _10447_ ;
wire _10027_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _9973_ ;
wire _9553_ ;
wire _9133_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _10676_ ;
wire _10256_ ;
wire _2598_ ;
wire _2178_ ;
wire _8824_ ;
wire _8404_ ;
wire _9609_ ;
wire _4744_ ;
wire _4324_ ;
wire breg_28_bF$buf0 ;
wire breg_28_bF$buf1 ;
wire breg_28_bF$buf2 ;
wire breg_28_bF$buf3 ;
wire breg_28_bF$buf4 ;
wire breg_28_bF$buf5 ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _9782_ ;
wire _9362_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _10485_ ;
wire _10065_ ;
wire breg_6_bF$buf0 ;
wire breg_6_bF$buf1 ;
wire breg_6_bF$buf2 ;
wire breg_6_bF$buf3 ;
wire breg_6_bF$buf4 ;
wire breg_6_bF$buf5 ;
wire _8633_ ;
wire _8213_ ;
wire _9838_ ;
wire _9418_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _9591_ ;
wire _9171_ ;
wire _1678_ ;
wire _1258_ ;
wire _7904_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _11902_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _10294_ ;
wire _4609_ ;
wire _8862_ ;
wire _8442_ ;
wire _8022_ ;
wire _11499_ ;
wire _11079_ ;
wire _9647_ ;
wire _9227_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _7713_ ;
wire _398_ ;
wire _11711_ ;
wire _8918_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _8671_ ;
wire _8251_ ;
wire _9876_ ;
wire _9456_ ;
wire _9036_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _7942_ ;
wire _7522_ ;
wire _7102_ ;
wire _10999_ ;
wire _10579_ ;
wire _10159_ ;
wire _11520_ ;
wire _11100_ ;
wire _8727_ ;
wire _8307_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _8480_ ;
wire _8060_ ;
wire _9685_ ;
wire _9265_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _7751_ ;
wire _7331_ ;
wire _10388_ ;
wire _8956_ ;
wire _8536_ ;
wire _8116_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _9494_ ;
wire _9074_ ;
wire _10600_ ;
wire _7807_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _11805_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _7980_ ;
wire _7560_ ;
wire _7140_ ;
wire _10197_ ;
wire _8765_ ;
wire _8345_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _7616_ ;
wire _2751_ ;
wire _2331_ ;
wire _11614_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _8994_ ;
wire _8574_ ;
wire _8154_ ;
wire _1602_ ;
wire _9779_ ;
wire _9359_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7845_ ;
wire _7425_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _11843_ ;
wire _11423_ ;
wire _11003_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _8383_ ;
wire _1831_ ;
wire _1411_ ;
wire _9588_ ;
wire _9168_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _7654_ ;
wire _7234_ ;
wire _11652_ ;
wire _11232_ ;
wire _8859_ ;
wire _8439_ ;
wire _8019_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _9800_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _8192_ ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _9397_ ;
wire _10923_ ;
wire _10503_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _11708_ ;
wire _7883_ ;
wire _7463_ ;
wire _7043_ ;
wire _11881_ ;
wire _11461_ ;
wire _11041_ ;
wire _8668_ ;
wire _8248_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _10732_ ;
wire _10312_ ;
wire _780_ ;
wire _360_ ;
wire _7939_ ;
wire _7519_ ;
wire _2654_ ;
wire _2234_ ;
wire _11517_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _7692_ ;
wire _7272_ ;
wire _11690_ ;
wire _11270_ ;
wire _8897_ ;
wire _8477_ ;
wire _8057_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _10961_ ;
wire _10541_ ;
wire _10121_ ;
wire _7748_ ;
wire _7328_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire areg_21_bF$buf0 ;
wire areg_21_bF$buf1 ;
wire areg_21_bF$buf2 ;
wire areg_21_bF$buf3 ;
wire areg_21_bF$buf4 ;
wire _11746_ ;
wire _11326_ ;
wire _3668_ ;
wire _3248_ ;
wire _7081_ ;
wire _5814_ ;
wire _8286_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _10770_ ;
wire _10350_ ;
wire _7977_ ;
wire _7557_ ;
wire _7137_ ;
wire _2692_ ;
wire _2272_ ;
wire _11555_ ;
wire _11135_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _9703_ ;
wire _5623_ ;
wire _5203_ ;
wire _8095_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _10826_ ;
wire _10406_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _7786_ ;
wire _7366_ ;
wire _2081_ ;
wire _11784_ ;
wire _11364_ ;
wire _3286_ ;
wire _9932_ ;
wire _9512_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _10635_ ;
wire _10215_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _7595_ ;
wire _7175_ ;
wire _11593_ ;
wire _11173_ ;
wire _5908_ ;
wire _3095_ ;
wire _9741_ ;
wire _9321_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _10864_ ;
wire _10444_ ;
wire _10024_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _11649_ ;
wire _11229_ ;
wire _4932_ ;
wire _4512_ ;
wire areg_3_bF$buf0 ;
wire areg_3_bF$buf1 ;
wire areg_3_bF$buf2 ;
wire areg_3_bF$buf3 ;
wire areg_3_bF$buf4 ;
wire _5717_ ;
wire _8189_ ;
wire _9970_ ;
wire _9550_ ;
wire _9130_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _10673_ ;
wire _10253_ ;
wire _2595_ ;
wire _2175_ ;
wire _8821_ ;
wire _8401_ ;
wire _11878_ ;
wire _11458_ ;
wire _11038_ ;
wire _9606_ ;
wire _4741_ ;
wire _4321_ ;
wire _7217__bF$buf0 ;
wire _7217__bF$buf1 ;
wire _7217__bF$buf2 ;
wire _7217__bF$buf3 ;
wire _7217__bF$buf4 ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _10729_ ;
wire _10309_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _10482_ ;
wire _10062_ ;
wire _7689_ ;
wire _7269_ ;
wire _8630_ ;
wire _8210_ ;
wire _11687_ ;
wire _11267_ ;
wire _3189_ ;
wire _9835_ ;
wire _9415_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _7901_ ;
wire _10958_ ;
wire _10538_ ;
wire _10118_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _10291_ ;
wire _4606_ ;
wire _7498_ ;
wire _7078_ ;
wire _11496_ ;
wire _11076_ ;
wire _9644_ ;
wire _9224_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _7710_ ;
wire _10767_ ;
wire _10347_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _8915_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _9873_ ;
wire _9453_ ;
wire _9033_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _3781__bF$buf0 ;
wire _3781__bF$buf1 ;
wire _6998_ ;
wire _3781__bF$buf2 ;
wire _6578_ ;
wire _3781__bF$buf3 ;
wire _6158_ ;
wire _1293_ ;
wire _10996_ ;
wire _10576_ ;
wire _10156_ ;
wire _2498_ ;
wire _2078_ ;
wire _8724_ ;
wire _8304_ ;
wire _9929_ ;
wire _9509_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _9682_ ;
wire _9262_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _10385_ ;
wire _8953_ ;
wire _8533_ ;
wire _8113_ ;
wire _9738_ ;
wire _9318_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _9491_ ;
wire _9071_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _7804_ ;
wire _489_ ;
wire _11802_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _10194_ ;
wire _4929_ ;
wire _4509_ ;
wire _8762_ ;
wire _8342_ ;
wire _11399_ ;
wire _9967_ ;
wire _9547_ ;
wire _9127_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _7613_ ;
wire _298_ ;
wire _11611_ ;
wire _8818_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _8991_ ;
wire _8571_ ;
wire _8151_ ;
wire _17_ ;
wire _9776_ ;
wire _9356_ ;
wire _4491_ ;
wire _4071_ ;
wire _3253__bF$buf0 ;
wire _3253__bF$buf1 ;
wire _3253__bF$buf2 ;
wire _3253__bF$buf3 ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7842_ ;
wire _7422_ ;
wire _7002_ ;
wire _10899_ ;
wire _10479_ ;
wire _10059_ ;
wire _11840_ ;
wire _11420_ ;
wire _11000_ ;
wire _8627_ ;
wire _8207_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _8380_ ;
wire _9585_ ;
wire _9165_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire _7651_ ;
wire _7231_ ;
wire _10288_ ;
wire _8856_ ;
wire _8436_ ;
wire _8016_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire _9394_ ;
wire _10920_ ;
wire _10500_ ;
wire _7707_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _11705_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7880_ ;
wire _7460_ ;
wire _7040_ ;
wire _10097_ ;
wire _8665_ ;
wire _8245_ ;
wire _3380_ ;
wire _3529__bF$buf0 ;
wire _3529__bF$buf1 ;
wire _3529__bF$buf2 ;
wire _3529__bF$buf3 ;
wire _3529__bF$buf4 ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _7936_ ;
wire _7516_ ;
wire _2651_ ;
wire _2231_ ;
wire breg_23_bF$buf0 ;
wire breg_23_bF$buf1 ;
wire breg_23_bF$buf2 ;
wire breg_23_bF$buf3 ;
wire _11514_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _8894_ ;
wire _8474_ ;
wire _8054_ ;
wire _1922_ ;
wire _1502_ ;
wire _9679_ ;
wire _9259_ ;
wire _4394_ ;
wire breg_1_bF$buf0 ;
wire breg_1_bF$buf1 ;
wire breg_1_bF$buf2 ;
wire breg_1_bF$buf3 ;
wire breg_1_bF$buf4 ;
wire _833_ ;
wire breg_1_bF$buf5 ;
wire _413_ ;
wire breg_1_bF$buf6 ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _7745_ ;
wire _7325_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _11743_ ;
wire _11323_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _8283_ ;
wire _1731_ ;
wire _1311_ ;
wire _9488_ ;
wire _9068_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _7974_ ;
wire _7520__bF$buf0 ;
wire _7554_ ;
wire _7520__bF$buf1 ;
wire _7134_ ;
wire _7520__bF$buf2 ;
wire _7520__bF$buf3 ;
wire _11552_ ;
wire _11132_ ;
wire _8759_ ;
wire _8339_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _9700_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _8092_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _9297_ ;
wire _10823_ ;
wire _10403_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _11608_ ;
wire _7783_ ;
wire _7363_ ;
wire _11781_ ;
wire _11361_ ;
wire _8988_ ;
wire _8568_ ;
wire _8148_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _10632_ ;
wire _10212_ ;
wire _680_ ;
wire _260_ ;
wire _7839_ ;
wire _7419_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _11837_ ;
wire _11417_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _7592_ ;
wire _7172_ ;
wire _11590_ ;
wire _11170_ ;
wire _5905_ ;
wire _8797_ ;
wire _8377_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire _10861_ ;
wire _10441_ ;
wire _10021_ ;
wire _7648_ ;
wire _7228_ ;
wire _2783_ ;
wire _2363_ ;
wire _11646_ ;
wire _11226_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _8186_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire _10917_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _10670_ ;
wire _10250_ ;
wire _7877_ ;
wire _7457_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _11875_ ;
wire _11455_ ;
wire _11035_ ;
wire _3797_ ;
wire _3377_ ;
wire _9603_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _10726_ ;
wire _10306_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _7686_ ;
wire _7266_ ;
wire _11684_ ;
wire _11264_ ;
wire _3186_ ;
wire _9832_ ;
wire _9412_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _10955_ ;
wire _10535_ ;
wire _10115_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _7495_ ;
wire _7075_ ;
wire _11493_ ;
wire _11073_ ;
wire _5808_ ;
wire _5668__bF$buf0 ;
wire _5668__bF$buf1 ;
wire _5668__bF$buf2 ;
wire _5668__bF$buf3 ;
wire _5668__bF$buf4 ;
wire _9641_ ;
wire _5668__bF$buf5 ;
wire _9221_ ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _10764_ ;
wire _10344_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _8912_ ;
wire _11549_ ;
wire _11129_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _8089_ ;
wire _9870_ ;
wire _9450_ ;
wire _9030_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _10993_ ;
wire _10573_ ;
wire _10153_ ;
wire _6044__bF$buf0 ;
wire _6044__bF$buf1 ;
wire _6044__bF$buf2 ;
wire _6044__bF$buf3 ;
wire _6044__bF$buf4 ;
wire _6044__bF$buf5 ;
wire _2495_ ;
wire _2075_ ;
wire _8721_ ;
wire _8301_ ;
wire _11778_ ;
wire _11358_ ;
wire _9926_ ;
wire _9506_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _10629_ ;
wire _10209_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _10382_ ;
wire _7589_ ;
wire _7169_ ;
wire _8950_ ;
wire _8530_ ;
wire _8110_ ;
wire _11587_ ;
wire _11167_ ;
wire _3089_ ;
wire _9735_ ;
wire _9315_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _7801_ ;
wire _10858_ ;
wire _10438_ ;
wire _10018_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _10191_ ;
wire _4926_ ;
wire _4506_ ;
wire _7398_ ;
wire _11396_ ;
wire _9964_ ;
wire _9544_ ;
wire _9124_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _7610_ ;
wire _10667_ ;
wire _10247_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _8815_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _9773_ ;
wire _9353_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _10896_ ;
wire _10476_ ;
wire _10056_ ;
wire _2398_ ;
wire _8624_ ;
wire _8204_ ;
wire _9829_ ;
wire _9409_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _9582_ ;
wire _9162_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _10285_ ;
wire _8853_ ;
wire _8433_ ;
wire _8013_ ;
wire _9638_ ;
wire _9218_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _9391_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _7704_ ;
wire _389_ ;
wire _11702_ ;
wire _8909_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _10094_ ;
wire _4829_ ;
wire _4409_ ;
wire _2884__bF$buf0 ;
wire _8662_ ;
wire _2884__bF$buf1 ;
wire _8242_ ;
wire _2884__bF$buf2 ;
wire _2884__bF$buf3 ;
wire _11299_ ;
wire _9867_ ;
wire _9447_ ;
wire _9027_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _3402__bF$buf0 ;
wire _3402__bF$buf1 ;
wire _3402__bF$buf2 ;
wire _3402__bF$buf3 ;
wire _7933_ ;
wire _7513_ ;
wire _198_ ;
wire _11511_ ;
wire _8718_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _8891_ ;
wire _8471_ ;
wire _8051_ ;
wire _9676_ ;
wire _9256_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _7742_ ;
wire _7322_ ;
wire _10799_ ;
wire _10379_ ;
wire _11740_ ;
wire _11320_ ;
wire _8947_ ;
wire _8527_ ;
wire _8107_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _8280_ ;
wire _9485_ ;
wire _9065_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _7971_ ;
wire _7551_ ;
wire _7131_ ;
wire _10188_ ;
wire _8756_ ;
wire _8336_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _9294_ ;
wire _10820_ ;
wire _10400_ ;
wire _7607_ ;
wire _2742_ ;
wire _2322_ ;
wire breg_15_bF$buf0 ;
wire breg_15_bF$buf1 ;
wire breg_15_bF$buf2 ;
wire breg_15_bF$buf3 ;
wire breg_15_bF$buf4 ;
wire breg_15_bF$buf5 ;
wire _11605_ ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _7780_ ;
wire _7360_ ;
wire _8985_ ;
wire _8565_ ;
wire _8145_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _7836_ ;
wire _7416_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _11834_ ;
wire _11414_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _8794_ ;
wire _8374_ ;
wire _1822_ ;
wire _1402_ ;
wire _9999_ ;
wire _9579_ ;
wire _9159_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire _7645_ ;
wire _7225_ ;
wire _2780_ ;
wire _2360_ ;
wire _11643_ ;
wire _11223_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _8183_ ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _9388_ ;
wire _10914_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _7874_ ;
wire _7454_ ;
wire _7034_ ;
wire _11872_ ;
wire _11452_ ;
wire _11032_ ;
wire _8659_ ;
wire _8239_ ;
wire _3794_ ;
wire _3374_ ;
wire _9600_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _9197_ ;
wire _10723_ ;
wire _10303_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _11508_ ;
wire _7683_ ;
wire _7263_ ;
wire _11681_ ;
wire _11261_ ;
wire _8888_ ;
wire _8468_ ;
wire _8048_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire _10952_ ;
wire _10532_ ;
wire _10112_ ;
wire _580_ ;
wire _160_ ;
wire _7739_ ;
wire _7319_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _11737_ ;
wire _11317_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _7492_ ;
wire _7072_ ;
wire _11490_ ;
wire _11070_ ;
wire _5805_ ;
wire _8697_ ;
wire _8277_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _10761_ ;
wire _10341_ ;
wire _7968_ ;
wire _7548_ ;
wire _7128_ ;
wire _2683_ ;
wire _2263_ ;
wire _11546_ ;
wire _11126_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _8086_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _10817_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _10990_ ;
wire _10570_ ;
wire _10150_ ;
wire _7777_ ;
wire _7357_ ;
wire _2492_ ;
wire _2072_ ;
wire _11775_ ;
wire _11355_ ;
wire _3697_ ;
wire _3277_ ;
wire _9923_ ;
wire _9503_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _10626_ ;
wire _10206_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _7586_ ;
wire _7166_ ;
wire _11584_ ;
wire _11164_ ;
wire _3086_ ;
wire _9732_ ;
wire _9312_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _10855_ ;
wire _10435_ ;
wire _10015_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _7395_ ;
wire _11393_ ;
wire _5708_ ;
wire _9961_ ;
wire _9541_ ;
wire _9121_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _10664_ ;
wire _10244_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _8812_ ;
wire _11869_ ;
wire _11449_ ;
wire _11029_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _9770_ ;
wire _9350_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _10893_ ;
wire _10473_ ;
wire _10053_ ;
wire _2395_ ;
wire _8621_ ;
wire _8201_ ;
wire _11678_ ;
wire _11258_ ;
wire _9826_ ;
wire _9406_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire areg_17_bF$buf0 ;
wire _1666_ ;
wire areg_17_bF$buf1 ;
wire _1246_ ;
wire areg_17_bF$buf2 ;
wire areg_17_bF$buf3 ;
wire areg_17_bF$buf4 ;
wire areg_17_bF$buf5 ;
wire _10949_ ;
wire _10529_ ;
wire _10109_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _10282_ ;
wire _7489_ ;
wire _7069_ ;
wire _8850_ ;
wire _8430_ ;
wire _8010_ ;
wire _11487_ ;
wire _11067_ ;
wire _9635_ ;
wire _9215_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _7701_ ;
wire _10758_ ;
wire _10338_ ;
wire _386_ ;
wire _8906_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _10091_ ;
wire _4826_ ;
wire _4406_ ;
wire _7298_ ;
wire _11296_ ;
wire _9864_ ;
wire _9444_ ;
wire _9024_ ;
wire _5784_ ;
wire _5364_ ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _7930_ ;
wire _7510_ ;
wire _10987_ ;
wire _10567_ ;
wire _10147_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _8715_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _9673_ ;
wire _9253_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _10796_ ;
wire _10376_ ;
wire _2298_ ;
wire _8944_ ;
wire _8524_ ;
wire _8104_ ;
wire _9729_ ;
wire _9309_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _9482_ ;
wire _9062_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _10185_ ;
wire _8753_ ;
wire _8333_ ;
wire _9958_ ;
wire _9538_ ;
wire _9118_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _9291_ ;
wire _1798_ ;
wire _1378_ ;
wire _7604_ ;
wire _289_ ;
wire _11602_ ;
wire _8809_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _8982_ ;
wire _8562_ ;
wire _8142_ ;
wire _11199_ ;
wire _9767_ ;
wire _9347_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _7833_ ;
wire _7413_ ;
wire _11831_ ;
wire _11411_ ;
wire _8618_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _8791_ ;
wire _8371_ ;
wire _9996_ ;
wire _9576_ ;
wire _9156_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _7642_ ;
wire _7222_ ;
wire _10699_ ;
wire _10279_ ;
wire _11640_ ;
wire _11220_ ;
wire _8847_ ;
wire _8427_ ;
wire _8007_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _8180_ ;
wire _46_ ;
wire _6913_ ;
wire _9385_ ;
wire _10911_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _7871_ ;
wire _7451_ ;
wire _7031_ ;
wire _10088_ ;
wire _8656_ ;
wire _8236_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _9194_ ;
wire _10720_ ;
wire _10300_ ;
wire _7927_ ;
wire _7507_ ;
wire _2642_ ;
wire _2222_ ;
wire _11505_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _7680_ ;
wire _7260_ ;
wire _8885_ ;
wire _8465_ ;
wire _8045_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire _7736_ ;
wire _7316_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _11734_ ;
wire _11314_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _8694_ ;
wire _8274_ ;
wire _1722_ ;
wire _1302_ ;
wire _9899_ ;
wire _9479_ ;
wire _9059_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _7965_ ;
wire _7545_ ;
wire _7125_ ;
wire _2680_ ;
wire _2260_ ;
wire _11543_ ;
wire _11123_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _8083_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _9288_ ;
wire _10814_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _7774_ ;
wire _7354_ ;
wire _11772_ ;
wire _11352_ ;
wire _8979_ ;
wire _8559_ ;
wire _8139_ ;
wire _3694_ ;
wire _3274_ ;
wire _9920_ ;
wire _9500_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _9097_ ;
wire _10623_ ;
wire _10203_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _11828_ ;
wire _11408_ ;
wire _7583_ ;
wire _7163_ ;
wire _11581_ ;
wire _11161_ ;
wire _8788_ ;
wire _8368_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire _10852_ ;
wire _10432_ ;
wire _10012_ ;
wire _480_ ;
wire _7639_ ;
wire _7219_ ;
wire _2774_ ;
wire _2354_ ;
wire _11637_ ;
wire _11217_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _7392_ ;
wire _11390_ ;
wire _5705_ ;
wire _8597_ ;
wire _8177_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _10908_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _10661_ ;
wire _10241_ ;
wire _7868_ ;
wire _7448_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _11866_ ;
wire _11446_ ;
wire _11026_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire breg_10_bF$buf0 ;
wire _5514_ ;
wire breg_10_bF$buf1 ;
wire breg_10_bF$buf2 ;
wire breg_10_bF$buf3 ;
wire breg_10_bF$buf4 ;
wire breg_10_bF$buf5 ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _10717_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire _6052_ ;
wire _6582__bF$buf0 ;
wire _6582__bF$buf1 ;
wire _6582__bF$buf2 ;
wire _6582__bF$buf3 ;
wire _10890_ ;
wire _10470_ ;
wire _10050_ ;
wire _7677_ ;
wire _7257_ ;
wire _2392_ ;
wire _11675_ ;
wire _11255_ ;
wire _3597_ ;
wire _3177_ ;
wire _9823_ ;
wire _9403_ ;
wire _5743_ ;
wire _5323_ ;
wire _7100__bF$buf0 ;
wire _7100__bF$buf1 ;
wire _7100__bF$buf2 ;
wire _7100__bF$buf3 ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _10946_ ;
wire _10526_ ;
wire _10106_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _7486_ ;
wire _7066_ ;
wire _11484_ ;
wire _11064_ ;
wire _9632_ ;
wire _9212_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _10755_ ;
wire _10335_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _8903_ ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _7295_ ;
wire _11293_ ;
wire _5608_ ;
wire _9861_ ;
wire _9441_ ;
wire _9021_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _10984_ ;
wire _10564_ ;
wire _10144_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _8712_ ;
wire _11769_ ;
wire _11349_ ;
wire _9917_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _9670_ ;
wire _9250_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire areg_28_bF$buf0 ;
wire areg_28_bF$buf1 ;
wire areg_28_bF$buf2 ;
wire areg_28_bF$buf3 ;
wire areg_28_bF$buf4 ;
wire areg_28_bF$buf5 ;
wire _3903_ ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _10793_ ;
wire _10373_ ;
wire _2295_ ;
wire _8941_ ;
wire _8521_ ;
wire _8101_ ;
wire _11578_ ;
wire _11158_ ;
wire _9726_ ;
wire _9306_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _10849_ ;
wire _10429_ ;
wire _10009_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _10182_ ;
wire _4917_ ;
wire _7389_ ;
wire _8750_ ;
wire _8330_ ;
wire _11387_ ;
wire _9955_ ;
wire _9535_ ;
wire _9115_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _7601_ ;
wire _10658_ ;
wire _10238_ ;
wire _286_ ;
wire _8806_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _7198_ ;
wire _11196_ ;
wire _9764_ ;
wire _9344_ ;
wire _5684_ ;
wire _5264_ ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _7830_ ;
wire _7410_ ;
wire _10887_ ;
wire _10467_ ;
wire _10047_ ;
wire _2389_ ;
wire _8615_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _9993_ ;
wire _9573_ ;
wire _9153_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _10696_ ;
wire _10276_ ;
wire _2198_ ;
wire _8844_ ;
wire _8424_ ;
wire _8004_ ;
wire _9629_ ;
wire _9209_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _6910_ ;
wire _9382_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _10085_ ;
wire _8653_ ;
wire _8233_ ;
wire _9858_ ;
wire _9438_ ;
wire _9018_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _9191_ ;
wire _1698_ ;
wire _1278_ ;
wire _7924_ ;
wire _7504_ ;
wire _189_ ;
wire _11502_ ;
wire _8709_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _8882_ ;
wire _8462_ ;
wire _8042_ ;
wire _11099_ ;
wire _1910_ ;
wire _9667_ ;
wire _9247_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _7733_ ;
wire _7313_ ;
wire _11731_ ;
wire _11311_ ;
wire _8938_ ;
wire _8518_ ;
wire _3653_ ;
wire _3233_ ;
wire areg_12_bF$buf0 ;
wire areg_12_bF$buf1 ;
wire areg_12_bF$buf2 ;
wire areg_12_bF$buf3 ;
wire areg_12_bF$buf4 ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _8691_ ;
wire _8271_ ;
wire _9896_ ;
wire _9476_ ;
wire _9056_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _7962_ ;
wire _7542_ ;
wire _7122_ ;
wire _10599_ ;
wire _10179_ ;
wire _11540_ ;
wire _11120_ ;
wire _8747_ ;
wire _8327_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _8080_ ;
wire _6813_ ;
wire _9285_ ;
wire _10811_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _7771_ ;
wire _7351_ ;
wire _8976_ ;
wire _8556_ ;
wire _8136_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _9094_ ;
wire _10620_ ;
wire _10200_ ;
wire _7827_ ;
wire _7407_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _11825_ ;
wire _11405_ ;
wire _3747_ ;
wire _3327_ ;
wire _7580_ ;
wire _7160_ ;
wire _8785_ ;
wire _8365_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire _7636_ ;
wire _7216_ ;
wire _2771_ ;
wire _2351_ ;
wire _11634_ ;
wire _11214_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _8594_ ;
wire _8174_ ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _9799_ ;
wire _9379_ ;
wire _4094_ ;
wire _10905_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7865_ ;
wire _7445_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _11863_ ;
wire _11443_ ;
wire _11023_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _9188_ ;
wire _10714_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _7674_ ;
wire _7254_ ;
wire _11672_ ;
wire _11252_ ;
wire _8879_ ;
wire _8459_ ;
wire _8039_ ;
wire _3594_ ;
wire _3174_ ;
wire _9820_ ;
wire _9400_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _10943_ ;
wire _10523_ ;
wire _10103_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _11728_ ;
wire _11308_ ;
wire _7483_ ;
wire _7063_ ;
wire _11481_ ;
wire _11061_ ;
wire _8688_ ;
wire _8268_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _10752_ ;
wire _10332_ ;
wire _380_ ;
wire _7959_ ;
wire _7539_ ;
wire _7119_ ;
wire _2674_ ;
wire _2254_ ;
wire _8900_ ;
wire _11537_ ;
wire _11117_ ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _7292_ ;
wire _11290_ ;
wire _5605_ ;
wire _8497_ ;
wire _8077_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _10808_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire _10981_ ;
wire _10561_ ;
wire _10141_ ;
wire _7768_ ;
wire _7348_ ;
wire _2483_ ;
wire _2063_ ;
wire _11766_ ;
wire _11346_ ;
wire _3688_ ;
wire _3268_ ;
wire _9914_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _10617_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _10790_ ;
wire _10370_ ;
wire _7997_ ;
wire _7577_ ;
wire _7157_ ;
wire _2292_ ;
wire _11575_ ;
wire _11155_ ;
wire _3497_ ;
wire _3077_ ;
wire _9723_ ;
wire _9303_ ;
wire _5643_ ;
wire _5223_ ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _10846_ ;
wire _10426_ ;
wire _10006_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _7386_ ;
wire _11384_ ;
wire _9952_ ;
wire _9532_ ;
wire _9112_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _10655_ ;
wire _10235_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _8803_ ;
wire _4723_ ;
wire _4303_ ;
wire _7195_ ;
wire _11193_ ;
wire _5928_ ;
wire _5508_ ;
wire _9761_ ;
wire _9341_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire _10884_ ;
wire _10464_ ;
wire _10044_ ;
wire _2386_ ;
wire _8612_ ;
wire _11669_ ;
wire _11249_ ;
wire _9817_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _9990_ ;
wire _9570_ ;
wire _9150_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _10693_ ;
wire _10273_ ;
wire _2195_ ;
wire _8841_ ;
wire _8421_ ;
wire _8001_ ;
wire _9104__bF$buf0 ;
wire _9104__bF$buf1 ;
wire _9104__bF$buf2 ;
wire _11898_ ;
wire _9104__bF$buf3 ;
wire _11478_ ;
wire _11058_ ;
wire _9626_ ;
wire _9206_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _10749_ ;
wire _10329_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _10082_ ;
wire _4817_ ;
wire _7289_ ;
wire _8650_ ;
wire _8230_ ;
wire _11287_ ;
wire _9855_ ;
wire _9435_ ;
wire _9015_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _7921_ ;
wire _7501_ ;
wire _10978_ ;
wire _10558_ ;
wire _10138_ ;
wire _186_ ;
wire _8706_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _7098_ ;
wire _11096_ ;
wire _9664_ ;
wire _9244_ ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _7730_ ;
wire _7310_ ;
wire _10787_ ;
wire _10367_ ;
wire _2289_ ;
wire _8935_ ;
wire _8515_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _9893_ ;
wire _9473_ ;
wire _9053_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _10596_ ;
wire _10176_ ;
wire _2098_ ;
wire _8744_ ;
wire _8324_ ;
wire _9949_ ;
wire _9529_ ;
wire _9109_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _9282_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _8973_ ;
wire _8553_ ;
wire _8133_ ;
wire _9758_ ;
wire _9338_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _9091_ ;
wire _1598_ ;
wire _1178_ ;
wire _7824_ ;
wire _7404_ ;
wire _11822_ ;
wire _11402_ ;
wire _8609_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _8782_ ;
wire _8362_ ;
wire areg_23_bF$buf0 ;
wire areg_23_bF$buf1 ;
wire areg_23_bF$buf2 ;
wire areg_23_bF$buf3 ;
wire areg_23_bF$buf4 ;
wire _1810_ ;
wire _9987_ ;
wire _9567_ ;
wire _9147_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _7633_ ;
wire _7213_ ;
wire _11631_ ;
wire _11211_ ;
wire _8838_ ;
wire _8418_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _8591_ ;
wire _8171_ ;
wire _37_ ;
wire _6904_ ;
wire _9796_ ;
wire _9376_ ;
wire _4091_ ;
wire _10902_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7862_ ;
wire _7442_ ;
wire _7022_ ;
wire _10499_ ;
wire _10079_ ;
wire _11860_ ;
wire _11440_ ;
wire _11020_ ;
wire _8647_ ;
wire _8227_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire _9185_ ;
wire _10711_ ;
wire _7918_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _7671_ ;
wire _7251_ ;
wire _8876_ ;
wire _8456_ ;
wire _8036_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _10940_ ;
wire _10520_ ;
wire _10100_ ;
wire _7727_ ;
wire _7307_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _11725_ ;
wire _11305_ ;
wire _3647_ ;
wire _3227_ ;
wire _7480_ ;
wire _7060_ ;
wire _8685_ ;
wire _8265_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire areg_5_bF$buf0 ;
wire areg_5_bF$buf1 ;
wire areg_5_bF$buf2 ;
wire areg_5_bF$buf3 ;
wire areg_5_bF$buf4 ;
wire _6751_ ;
wire _6331_ ;
wire _7956_ ;
wire _7536_ ;
wire _7116_ ;
wire _2671_ ;
wire _2251_ ;
wire _11534_ ;
wire _11114_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5420__bF$buf0 ;
wire _5420__bF$buf1 ;
wire _5420__bF$buf2 ;
wire _5420__bF$buf3 ;
wire _5602_ ;
wire _8494_ ;
wire _8074_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _9699_ ;
wire _9279_ ;
wire _10805_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire _7765_ ;
wire _7345_ ;
wire _2480_ ;
wire _2060_ ;
wire _11763_ ;
wire _11343_ ;
wire _3685_ ;
wire _3265_ ;
wire _9911_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _9088_ ;
wire _10614_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _11819_ ;
wire _7994_ ;
wire _7574_ ;
wire _7154_ ;
wire _11572_ ;
wire _11152_ ;
wire _8779_ ;
wire _8359_ ;
wire _3494_ ;
wire _3074_ ;
wire _9720_ ;
wire _9300_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _10843_ ;
wire _10423_ ;
wire _10003_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _11628_ ;
wire _11208_ ;
wire _4911_ ;
wire _7383_ ;
wire _11381_ ;
wire _8588_ ;
wire _8168_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _10652_ ;
wire _10232_ ;
wire _280_ ;
wire _7859_ ;
wire _7439_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _8800_ ;
wire _11857_ ;
wire _11437_ ;
wire _11017_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _7192_ ;
wire _11190_ ;
wire _5925_ ;
wire _5505_ ;
wire _8397_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _10708_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire _10881_ ;
wire _10461_ ;
wire _10041_ ;
wire _7668_ ;
wire _7248_ ;
wire _2383_ ;
wire _11666_ ;
wire _11246_ ;
wire _3588_ ;
wire _3168_ ;
wire _9814_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _10937_ ;
wire _10517_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _10690_ ;
wire _10270_ ;
wire _7897_ ;
wire _7477_ ;
wire _7057_ ;
wire _2192_ ;
wire _11895_ ;
wire _11475_ ;
wire _11055_ ;
wire _3397_ ;
wire _9623_ ;
wire _9203_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _10746_ ;
wire _10326_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _7286_ ;
wire _11284_ ;
wire _9852_ ;
wire _9432_ ;
wire _9012_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _10975_ ;
wire _10555_ ;
wire _10135_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _8703_ ;
wire _9908_ ;
wire _4623_ ;
wire _4203_ ;
wire _7095_ ;
wire _11093_ ;
wire _5828_ ;
wire _5408_ ;
wire _9661_ ;
wire _9241_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _10784_ ;
wire _10364_ ;
wire _2286_ ;
wire _8932_ ;
wire _8512_ ;
wire _11569_ ;
wire _11149_ ;
wire _9717_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _9890_ ;
wire _9470_ ;
wire _9050_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _10593_ ;
wire _10173_ ;
wire _4908_ ;
wire _2095_ ;
wire _8741_ ;
wire _8321_ ;
wire _11798_ ;
wire _11378_ ;
wire _9946_ ;
wire _9526_ ;
wire _9106_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _10649_ ;
wire _10229_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _7189_ ;
wire _8970_ ;
wire _8550_ ;
wire _8130_ ;
wire breg_25_bF$buf0 ;
wire _11187_ ;
wire breg_25_bF$buf1 ;
wire breg_25_bF$buf2 ;
wire breg_25_bF$buf3 ;
wire breg_25_bF$buf4 ;
wire breg_25_bF$buf5 ;
wire _9755_ ;
wire _9335_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _7821_ ;
wire _7401_ ;
wire _10878_ ;
wire _10458_ ;
wire _10038_ ;
wire breg_3_bF$buf0 ;
wire breg_3_bF$buf1 ;
wire breg_3_bF$buf2 ;
wire breg_3_bF$buf3 ;
wire breg_3_bF$buf4 ;
wire breg_3_bF$buf5 ;
wire _8606_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _9984_ ;
wire _9564_ ;
wire _9144_ ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _7630_ ;
wire _7210_ ;
wire _10687_ ;
wire _10267_ ;
wire _2189_ ;
wire _8835_ ;
wire _8415_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _6901_ ;
wire _9793_ ;
wire _9373_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _10496_ ;
wire _10076_ ;
wire _8644_ ;
wire _8224_ ;
wire _9849_ ;
wire _9429_ ;
wire _9009_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _9182_ ;
wire _1689_ ;
wire _1269_ ;
wire _7915_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _8873_ ;
wire _8453_ ;
wire _8033_ ;
wire _1901_ ;
wire _9658_ ;
wire _9238_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _7724_ ;
wire _7304_ ;
wire _11722_ ;
wire _11302_ ;
wire _8929_ ;
wire _8509_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _8682_ ;
wire _8262_ ;
wire _1710_ ;
wire _9887_ ;
wire _9467_ ;
wire _9047_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _7953_ ;
wire _7533_ ;
wire _7113_ ;
wire _11531_ ;
wire _11111_ ;
wire _8738_ ;
wire _8318_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _8491_ ;
wire _8071_ ;
wire _6804_ ;
wire _9696_ ;
wire _9276_ ;
wire _10802_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _7762_ ;
wire _7342_ ;
wire _10399_ ;
wire _11760_ ;
wire _11340_ ;
wire _8967_ ;
wire _8547_ ;
wire _8127_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _6613_ ;
wire _9085_ ;
wire _10611_ ;
wire _7818_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _11816_ ;
wire _3738_ ;
wire _3318_ ;
wire _7991_ ;
wire _7571_ ;
wire _7151_ ;
wire _8776_ ;
wire _8356_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _10840_ ;
wire _10420_ ;
wire _10000_ ;
wire _7627_ ;
wire _7207_ ;
wire _2762_ ;
wire _2342_ ;
wire _11625_ ;
wire _11205_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _7380_ ;
wire _8585_ ;
wire _8165_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7856_ ;
wire _7436_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _11854_ ;
wire _11434_ ;
wire _11014_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _8394_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _9599_ ;
wire _9179_ ;
wire _10705_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire _7665_ ;
wire _7245_ ;
wire _2380_ ;
wire _11663_ ;
wire _11243_ ;
wire _3585_ ;
wire _3165_ ;
wire _9811_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _10934_ ;
wire _10514_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _11719_ ;
wire _7894_ ;
wire _7474_ ;
wire _7054_ ;
wire _11892_ ;
wire _11472_ ;
wire _11052_ ;
wire _8679_ ;
wire _8259_ ;
wire _3394_ ;
wire _9620_ ;
wire _9200_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _10743_ ;
wire _10323_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _11528_ ;
wire _11108_ ;
wire _4811_ ;
wire _7283_ ;
wire _11281_ ;
wire _8488_ ;
wire _8068_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _10972_ ;
wire _10552_ ;
wire _10132_ ;
wire _180_ ;
wire _7759_ ;
wire _7339_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _8700_ ;
wire _11757_ ;
wire _11337_ ;
wire _3679_ ;
wire _3259_ ;
wire _9905_ ;
wire _4620_ ;
wire _4200_ ;
wire _7092_ ;
wire _11090_ ;
wire _5825_ ;
wire _5405_ ;
wire _8297_ ;
wire _1745_ ;
wire _1325_ ;
wire _10608_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _10781_ ;
wire _10361_ ;
wire _7988_ ;
wire _7568_ ;
wire _7148_ ;
wire _2283_ ;
wire _11566_ ;
wire _11146_ ;
wire _3488_ ;
wire _3068_ ;
wire _9714_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _10837_ ;
wire _10417_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _10590_ ;
wire _10170_ ;
wire _4905_ ;
wire _7797_ ;
wire _7377_ ;
wire _2092_ ;
wire _11795_ ;
wire _11375_ ;
wire _3297_ ;
wire _9943_ ;
wire _9523_ ;
wire _9103_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _10646_ ;
wire _10226_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _7186_ ;
wire _11184_ ;
wire _5919_ ;
wire _9752_ ;
wire _9332_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire _10875_ ;
wire _10455_ ;
wire _10035_ ;
wire _2797_ ;
wire _2377_ ;
wire _549__bF$buf0 ;
wire _549__bF$buf1 ;
wire _549__bF$buf2 ;
wire _549__bF$buf3 ;
wire _549__bF$buf4 ;
wire _8603_ ;
wire _9808_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _9981_ ;
wire _9561_ ;
wire _9141_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _10684_ ;
wire _10264_ ;
wire _2186_ ;
wire _8832_ ;
wire _8412_ ;
wire _11889_ ;
wire _11469_ ;
wire _11049_ ;
wire _9617_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _9790_ ;
wire _9370_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _10493_ ;
wire _10073_ ;
wire _4808_ ;
wire _8641_ ;
wire _8221_ ;
wire _11698_ ;
wire _11278_ ;
wire breg_17_bF$buf0 ;
wire breg_17_bF$buf1 ;
wire breg_17_bF$buf2 ;
wire breg_17_bF$buf3 ;
wire breg_17_bF$buf4 ;
wire _9846_ ;
wire _9426_ ;
wire _9006_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _7912_ ;
wire _10969_ ;
wire _10549_ ;
wire _10129_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _7089_ ;
wire _8870_ ;
wire _8450_ ;
wire _8030_ ;
wire _11087_ ;
wire _9655_ ;
wire _9235_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _7721_ ;
wire _7301_ ;
wire _10778_ ;
wire _10358_ ;
wire _8926_ ;
wire _8506_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _9884_ ;
wire _9464_ ;
wire _9044_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _7950_ ;
wire _7530_ ;
wire _7110_ ;
wire _10587_ ;
wire _10167_ ;
wire _2089_ ;
wire _8735_ ;
wire _8315_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _9693_ ;
wire _9273_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _2560__bF$buf0 ;
wire _2560__bF$buf1 ;
wire _2560__bF$buf2 ;
wire _10396_ ;
wire _2560__bF$buf3 ;
wire _2560__bF$buf4 ;
wire _8964_ ;
wire _8544_ ;
wire _8124_ ;
wire _9749_ ;
wire _9329_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _9082_ ;
wire _1589_ ;
wire _1169_ ;
wire _7815_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _11813_ ;
wire _3735_ ;
wire _3315_ ;
wire _8773_ ;
wire _8353_ ;
wire _1801_ ;
wire _9978_ ;
wire _9558_ ;
wire _9138_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _7624_ ;
wire _7204_ ;
wire _11622_ ;
wire _11202_ ;
wire _8829_ ;
wire _8409_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _8582_ ;
wire _8162_ ;
wire _28_ ;
wire _1610_ ;
wire _9787_ ;
wire _9367_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _7853_ ;
wire _7433_ ;
wire _7013_ ;
wire _11851_ ;
wire _11431_ ;
wire _11011_ ;
wire _8638_ ;
wire _8218_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _8391_ ;
wire _6704_ ;
wire _9596_ ;
wire _9176_ ;
wire _10702_ ;
wire _750_ ;
wire _330_ ;
wire _7909_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire breg_20_bF$buf0 ;
wire breg_20_bF$buf1 ;
wire _11907_ ;
wire breg_20_bF$buf2 ;
wire breg_20_bF$buf3 ;
wire breg_20_bF$buf4 ;
wire _3829_ ;
wire _3409_ ;
wire _7662_ ;
wire _7242_ ;
wire _10299_ ;
wire _11660_ ;
wire _11240_ ;
wire _8867_ ;
wire _8447_ ;
wire _8027_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _10931_ ;
wire _10511_ ;
wire _7718_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _11716_ ;
wire _3638_ ;
wire _3218_ ;
wire _7891_ ;
wire _7471_ ;
wire _7051_ ;
wire _8676_ ;
wire _8256_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _10740_ ;
wire _10320_ ;
wire _7947_ ;
wire _7527_ ;
wire _7107_ ;
wire _2662_ ;
wire _2242_ ;
wire _11525_ ;
wire _11105_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _7280_ ;
wire _8485_ ;
wire _8065_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _7756_ ;
wire _7336_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _11754_ ;
wire _11334_ ;
wire _3676_ ;
wire _3256_ ;
wire _9902_ ;
wire _5822_ ;
wire _5402_ ;
wire _8294_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _9499_ ;
wire _9079_ ;
wire _10605_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _7985_ ;
wire _7565_ ;
wire _7145_ ;
wire areg_19_bF$buf0 ;
wire areg_19_bF$buf1 ;
wire areg_19_bF$buf2 ;
wire _2280_ ;
wire areg_19_bF$buf3 ;
wire areg_19_bF$buf4 ;
wire areg_19_bF$buf5 ;
wire _11563_ ;
wire _11143_ ;
wire _3485_ ;
wire _3065_ ;
wire _9711_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _10834_ ;
wire _10414_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _11619_ ;
wire _4902_ ;
wire _7794_ ;
wire _7374_ ;
wire _11792_ ;
wire _11372_ ;
wire _8999_ ;
wire _8579_ ;
wire _8159_ ;
wire _3294_ ;
wire _9940_ ;
wire _9520_ ;
wire _9100_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _10643_ ;
wire _10223_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _11848_ ;
wire _11428_ ;
wire _11008_ ;
wire _4711_ ;
wire _7183_ ;
wire _11181_ ;
wire _5916_ ;
wire _8388_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire _10872_ ;
wire _10452_ ;
wire _10032_ ;
wire _7659_ ;
wire _7239_ ;
wire _2794_ ;
wire _2374_ ;
wire _8600_ ;
wire _11657_ ;
wire _11237_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _9805_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _8197_ ;
wire _1645_ ;
wire _1225_ ;
wire _10928_ ;
wire _10508_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _10681_ ;
wire _10261_ ;
wire _7888_ ;
wire _7468_ ;
wire _7048_ ;
wire _2183_ ;
wire _11886_ ;
wire _11466_ ;
wire _11046_ ;
wire _3388_ ;
wire _9614_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _10737_ ;
wire _10317_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _10490_ ;
wire _10070_ ;
wire _4805_ ;
wire _7697_ ;
wire _7277_ ;
wire _11695_ ;
wire _11275_ ;
wire _3197_ ;
wire _9843_ ;
wire _9423_ ;
wire _9003_ ;
wire _5763_ ;
wire _5343_ ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _10966_ ;
wire _10546_ ;
wire _10126_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _7086_ ;
wire _11084_ ;
wire _5819_ ;
wire _9652_ ;
wire _9232_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _7711__bF$buf0 ;
wire _7711__bF$buf1 ;
wire _7711__bF$buf2 ;
wire _7711__bF$buf3 ;
wire _10775_ ;
wire _10355_ ;
wire _2697_ ;
wire _2277_ ;
wire _8923_ ;
wire _8503_ ;
wire _9708_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _9881_ ;
wire _9461_ ;
wire _9041_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _10584_ ;
wire _10164_ ;
wire _2086_ ;
wire _8732_ ;
wire _8312_ ;
wire _11789_ ;
wire _11369_ ;
wire _9937_ ;
wire _9517_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _9690_ ;
wire _9270_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _10393_ ;
wire _4708_ ;
wire _8961_ ;
wire _8541_ ;
wire _8121_ ;
wire _11598_ ;
wire _11178_ ;
wire _9746_ ;
wire _9326_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _7812_ ;
wire _10869_ ;
wire _10449_ ;
wire _10029_ ;
wire _497_ ;
wire _11810_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _8770_ ;
wire _8350_ ;
wire _9975_ ;
wire _9555_ ;
wire _9135_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _7621_ ;
wire _7201_ ;
wire _10678_ ;
wire _10258_ ;
wire _8826_ ;
wire _8406_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _2465__bF$buf0 ;
wire _2465__bF$buf1 ;
wire _2465__bF$buf2 ;
wire _2465__bF$buf3 ;
wire _2465__bF$buf4 ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _9784_ ;
wire _9364_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7850_ ;
wire _7430_ ;
wire _7010_ ;
wire _10487_ ;
wire _10067_ ;
wire _8635_ ;
wire _8215_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _9593_ ;
wire _9173_ ;
wire _7906_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _11904_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _10296_ ;
wire _8864_ ;
wire _8444_ ;
wire _8024_ ;
wire _9649_ ;
wire _9229_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _7715_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _11713_ ;
wire _3635_ ;
wire _3215_ ;
wire _8673_ ;
wire _8253_ ;
wire _1701_ ;
wire _9878_ ;
wire _9458_ ;
wire _9038_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _7944_ ;
wire _7524_ ;
wire _7104_ ;
wire _11522_ ;
wire _11102_ ;
wire _10869__bF$buf0 ;
wire _10869__bF$buf1 ;
wire _8729_ ;
wire _10869__bF$buf2 ;
wire _8309_ ;
wire _10869__bF$buf3 ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _8482_ ;
wire _8062_ ;
wire _1930_ ;
wire _1510_ ;
wire _9687_ ;
wire _9267_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire breg_12_bF$buf0 ;
wire breg_12_bF$buf1 ;
wire breg_12_bF$buf2 ;
wire breg_12_bF$buf3 ;
wire breg_12_bF$buf4 ;
wire _7753_ ;
wire _7333_ ;
wire _11751_ ;
wire _11331_ ;
wire _8958_ ;
wire _8538_ ;
wire _8118_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _8291_ ;
wire _6604_ ;
wire _9496_ ;
wire _9076_ ;
wire _10602_ ;
wire _650_ ;
wire _230_ ;
wire _7809_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _11807_ ;
wire _3729_ ;
wire _3309_ ;
wire _7982_ ;
wire _7562_ ;
wire _7142_ ;
wire _10199_ ;
wire _11560_ ;
wire _11140_ ;
wire _8767_ ;
wire _8347_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _10831_ ;
wire _10411_ ;
wire _7618_ ;
wire _2753_ ;
wire _2333_ ;
wire _11616_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _7791_ ;
wire _7371_ ;
wire _8996_ ;
wire _8576_ ;
wire _8156_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _10640_ ;
wire _10220_ ;
wire _7847_ ;
wire _7427_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _11845_ ;
wire _11425_ ;
wire _11005_ ;
wire _3767_ ;
wire _3347_ ;
wire _7180_ ;
wire _5913_ ;
wire _8385_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire _7656_ ;
wire _7236_ ;
wire _2791_ ;
wire _2371_ ;
wire _11654_ ;
wire _11234_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _9802_ ;
wire _5722_ ;
wire _5302_ ;
wire _8194_ ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _9399_ ;
wire _10925_ ;
wire _10505_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7885_ ;
wire _7465_ ;
wire _7045_ ;
wire _2180_ ;
wire _11883_ ;
wire _11463_ ;
wire _11043_ ;
wire _3385_ ;
wire _9611_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _10734_ ;
wire _10314_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _11519_ ;
wire _4802_ ;
wire _7694_ ;
wire _7274_ ;
wire _11692_ ;
wire _11272_ ;
wire _8899_ ;
wire _8479_ ;
wire _8059_ ;
wire _3194_ ;
wire _9840_ ;
wire _9420_ ;
wire _9000_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _10963_ ;
wire _10543_ ;
wire _10123_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _11748_ ;
wire _11328_ ;
wire _4611_ ;
wire _7083_ ;
wire _11081_ ;
wire _5816_ ;
wire _8288_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire _10772_ ;
wire _10352_ ;
wire _7979_ ;
wire _7559_ ;
wire _7139_ ;
wire _2694_ ;
wire _2274_ ;
wire _8920_ ;
wire _8500_ ;
wire _11557_ ;
wire _11137_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _9705_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _8097_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _10828_ ;
wire _10408_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _10581_ ;
wire _10161_ ;
wire _7788_ ;
wire _7368_ ;
wire _2083_ ;
wire _11786_ ;
wire _11366_ ;
wire _3288_ ;
wire _9934_ ;
wire _9514_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _10637_ ;
wire _10217_ ;
wire _2551__bF$buf0 ;
wire _2551__bF$buf1 ;
wire _2551__bF$buf2 ;
wire _2551__bF$buf3 ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _10390_ ;
wire _4705_ ;
wire _7597_ ;
wire _7177_ ;
wire _11595_ ;
wire _11175_ ;
wire _3097_ ;
wire _9743_ ;
wire _9323_ ;
wire _5663_ ;
wire _5243_ ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _10866_ ;
wire _10446_ ;
wire _10026_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _9972_ ;
wire _9552_ ;
wire _9132_ ;
wire _1639_ ;
wire _1219_ ;
wire areg_14_bF$buf0 ;
wire areg_14_bF$buf1 ;
wire areg_14_bF$buf2 ;
wire areg_14_bF$buf3 ;
wire areg_14_bF$buf4 ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _10675_ ;
wire _10255_ ;
wire _2597_ ;
wire _2177_ ;
wire _8823_ ;
wire _8403_ ;
wire _9608_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _9781_ ;
wire _9361_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;
wire _10484_ ;
wire _10064_ ;
wire _8632_ ;
wire _8212_ ;

BUFX2 BUFX2_insert536 (
    .A(areg[30]),
    .Y(areg_30_bF$buf0)
);

BUFX2 BUFX2_insert535 (
    .A(areg[30]),
    .Y(areg_30_bF$buf1)
);

BUFX2 BUFX2_insert534 (
    .A(areg[30]),
    .Y(areg_30_bF$buf2)
);

BUFX2 BUFX2_insert533 (
    .A(areg[30]),
    .Y(areg_30_bF$buf3)
);

BUFX2 BUFX2_insert532 (
    .A(areg[30]),
    .Y(areg_30_bF$buf4)
);

BUFX2 BUFX2_insert531 (
    .A(areg[30]),
    .Y(areg_30_bF$buf5)
);

BUFX2 BUFX2_insert530 (
    .A(_2465_),
    .Y(_2465__bF$buf0)
);

BUFX2 BUFX2_insert529 (
    .A(_2465_),
    .Y(_2465__bF$buf1)
);

BUFX2 BUFX2_insert528 (
    .A(_2465_),
    .Y(_2465__bF$buf2)
);

BUFX2 BUFX2_insert527 (
    .A(_2465_),
    .Y(_2465__bF$buf3)
);

BUFX2 BUFX2_insert526 (
    .A(_2465_),
    .Y(_2465__bF$buf4)
);

BUFX2 BUFX2_insert525 (
    .A(_2562_),
    .Y(_2562__bF$buf0)
);

BUFX2 BUFX2_insert524 (
    .A(_2562_),
    .Y(_2562__bF$buf1)
);

BUFX2 BUFX2_insert523 (
    .A(_2562_),
    .Y(_2562__bF$buf2)
);

BUFX2 BUFX2_insert522 (
    .A(_2562_),
    .Y(_2562__bF$buf3)
);

BUFX2 BUFX2_insert521 (
    .A(_2562_),
    .Y(_2562__bF$buf4)
);

BUFX2 BUFX2_insert520 (
    .A(_3958_),
    .Y(_3958__bF$buf0)
);

BUFX2 BUFX2_insert519 (
    .A(_3958_),
    .Y(_3958__bF$buf1)
);

BUFX2 BUFX2_insert518 (
    .A(_3958_),
    .Y(_3958__bF$buf2)
);

BUFX2 BUFX2_insert517 (
    .A(_3958_),
    .Y(_3958__bF$buf3)
);

BUFX2 BUFX2_insert516 (
    .A(_3253_),
    .Y(_3253__bF$buf0)
);

BUFX2 BUFX2_insert515 (
    .A(_3253_),
    .Y(_3253__bF$buf1)
);

BUFX2 BUFX2_insert514 (
    .A(_3253_),
    .Y(_3253__bF$buf2)
);

BUFX2 BUFX2_insert513 (
    .A(_3253_),
    .Y(_3253__bF$buf3)
);

BUFX2 BUFX2_insert512 (
    .A(_3961_),
    .Y(_3961__bF$buf0)
);

BUFX2 BUFX2_insert511 (
    .A(_3961_),
    .Y(_3961__bF$buf1)
);

BUFX2 BUFX2_insert510 (
    .A(_3961_),
    .Y(_3961__bF$buf2)
);

BUFX2 BUFX2_insert509 (
    .A(_3961_),
    .Y(_3961__bF$buf3)
);

BUFX2 BUFX2_insert508 (
    .A(_3961_),
    .Y(_3961__bF$buf4)
);

BUFX2 BUFX2_insert507 (
    .A(_10869_),
    .Y(_10869__bF$buf0)
);

BUFX2 BUFX2_insert506 (
    .A(_10869_),
    .Y(_10869__bF$buf1)
);

BUFX2 BUFX2_insert505 (
    .A(_10869_),
    .Y(_10869__bF$buf2)
);

BUFX2 BUFX2_insert504 (
    .A(_10869_),
    .Y(_10869__bF$buf3)
);

BUFX2 BUFX2_insert503 (
    .A(_5190_),
    .Y(_5190__bF$buf0)
);

BUFX2 BUFX2_insert502 (
    .A(_5190_),
    .Y(_5190__bF$buf1)
);

BUFX2 BUFX2_insert501 (
    .A(_5190_),
    .Y(_5190__bF$buf2)
);

BUFX2 BUFX2_insert500 (
    .A(_5190_),
    .Y(_5190__bF$buf3)
);

BUFX2 BUFX2_insert499 (
    .A(breg[11]),
    .Y(breg_11_bF$buf0)
);

BUFX2 BUFX2_insert498 (
    .A(breg[11]),
    .Y(breg_11_bF$buf1)
);

BUFX2 BUFX2_insert497 (
    .A(breg[11]),
    .Y(breg_11_bF$buf2)
);

BUFX2 BUFX2_insert496 (
    .A(breg[11]),
    .Y(breg_11_bF$buf3)
);

BUFX2 BUFX2_insert495 (
    .A(breg[11]),
    .Y(breg_11_bF$buf4)
);

BUFX2 BUFX2_insert494 (
    .A(_6686_),
    .Y(_6686__bF$buf0)
);

BUFX2 BUFX2_insert493 (
    .A(_6686_),
    .Y(_6686__bF$buf1)
);

BUFX2 BUFX2_insert492 (
    .A(_6686_),
    .Y(_6686__bF$buf2)
);

BUFX2 BUFX2_insert491 (
    .A(_6686_),
    .Y(_6686__bF$buf3)
);

BUFX2 BUFX2_insert490 (
    .A(breg[2]),
    .Y(breg_2_bF$buf0)
);

BUFX2 BUFX2_insert489 (
    .A(breg[2]),
    .Y(breg_2_bF$buf1)
);

BUFX2 BUFX2_insert488 (
    .A(breg[2]),
    .Y(breg_2_bF$buf2)
);

BUFX2 BUFX2_insert487 (
    .A(breg[2]),
    .Y(breg_2_bF$buf3)
);

BUFX2 BUFX2_insert486 (
    .A(breg[2]),
    .Y(breg_2_bF$buf4)
);

BUFX2 BUFX2_insert485 (
    .A(breg[14]),
    .Y(breg_14_bF$buf0)
);

BUFX2 BUFX2_insert484 (
    .A(breg[14]),
    .Y(breg_14_bF$buf1)
);

BUFX2 BUFX2_insert483 (
    .A(breg[14]),
    .Y(breg_14_bF$buf2)
);

BUFX2 BUFX2_insert482 (
    .A(breg[14]),
    .Y(breg_14_bF$buf3)
);

BUFX2 BUFX2_insert481 (
    .A(breg[5]),
    .Y(breg_5_bF$buf0)
);

BUFX2 BUFX2_insert480 (
    .A(breg[5]),
    .Y(breg_5_bF$buf1)
);

BUFX2 BUFX2_insert479 (
    .A(breg[5]),
    .Y(breg_5_bF$buf2)
);

BUFX2 BUFX2_insert478 (
    .A(breg[5]),
    .Y(breg_5_bF$buf3)
);

BUFX2 BUFX2_insert477 (
    .A(breg[17]),
    .Y(breg_17_bF$buf0)
);

BUFX2 BUFX2_insert476 (
    .A(breg[17]),
    .Y(breg_17_bF$buf1)
);

BUFX2 BUFX2_insert475 (
    .A(breg[17]),
    .Y(breg_17_bF$buf2)
);

BUFX2 BUFX2_insert474 (
    .A(breg[17]),
    .Y(breg_17_bF$buf3)
);

BUFX2 BUFX2_insert473 (
    .A(breg[17]),
    .Y(breg_17_bF$buf4)
);

BUFX2 BUFX2_insert472 (
    .A(breg[20]),
    .Y(breg_20_bF$buf0)
);

BUFX2 BUFX2_insert471 (
    .A(breg[20]),
    .Y(breg_20_bF$buf1)
);

BUFX2 BUFX2_insert470 (
    .A(breg[20]),
    .Y(breg_20_bF$buf2)
);

BUFX2 BUFX2_insert469 (
    .A(breg[20]),
    .Y(breg_20_bF$buf3)
);

BUFX2 BUFX2_insert468 (
    .A(breg[20]),
    .Y(breg_20_bF$buf4)
);

BUFX2 BUFX2_insert467 (
    .A(areg[10]),
    .Y(areg_10_bF$buf0)
);

BUFX2 BUFX2_insert466 (
    .A(areg[10]),
    .Y(areg_10_bF$buf1)
);

BUFX2 BUFX2_insert465 (
    .A(areg[10]),
    .Y(areg_10_bF$buf2)
);

BUFX2 BUFX2_insert464 (
    .A(areg[10]),
    .Y(areg_10_bF$buf3)
);

BUFX2 BUFX2_insert463 (
    .A(areg[10]),
    .Y(areg_10_bF$buf4)
);

BUFX2 BUFX2_insert462 (
    .A(breg[23]),
    .Y(breg_23_bF$buf0)
);

BUFX2 BUFX2_insert461 (
    .A(breg[23]),
    .Y(breg_23_bF$buf1)
);

BUFX2 BUFX2_insert460 (
    .A(breg[23]),
    .Y(breg_23_bF$buf2)
);

BUFX2 BUFX2_insert459 (
    .A(breg[23]),
    .Y(breg_23_bF$buf3)
);

BUFX2 BUFX2_insert458 (
    .A(areg[13]),
    .Y(areg_13_bF$buf0)
);

BUFX2 BUFX2_insert457 (
    .A(areg[13]),
    .Y(areg_13_bF$buf1)
);

BUFX2 BUFX2_insert456 (
    .A(areg[13]),
    .Y(areg_13_bF$buf2)
);

BUFX2 BUFX2_insert455 (
    .A(areg[13]),
    .Y(areg_13_bF$buf3)
);

BUFX2 BUFX2_insert454 (
    .A(areg[13]),
    .Y(areg_13_bF$buf4)
);

BUFX2 BUFX2_insert453 (
    .A(_5420_),
    .Y(_5420__bF$buf0)
);

BUFX2 BUFX2_insert452 (
    .A(_5420_),
    .Y(_5420__bF$buf1)
);

BUFX2 BUFX2_insert451 (
    .A(_5420_),
    .Y(_5420__bF$buf2)
);

BUFX2 BUFX2_insert450 (
    .A(_5420_),
    .Y(_5420__bF$buf3)
);

BUFX2 BUFX2_insert449 (
    .A(breg[26]),
    .Y(breg_26_bF$buf0)
);

BUFX2 BUFX2_insert448 (
    .A(breg[26]),
    .Y(breg_26_bF$buf1)
);

BUFX2 BUFX2_insert447 (
    .A(breg[26]),
    .Y(breg_26_bF$buf2)
);

BUFX2 BUFX2_insert446 (
    .A(breg[26]),
    .Y(breg_26_bF$buf3)
);

BUFX2 BUFX2_insert445 (
    .A(breg[26]),
    .Y(breg_26_bF$buf4)
);

BUFX2 BUFX2_insert444 (
    .A(areg[16]),
    .Y(areg_16_bF$buf0)
);

BUFX2 BUFX2_insert443 (
    .A(areg[16]),
    .Y(areg_16_bF$buf1)
);

BUFX2 BUFX2_insert442 (
    .A(areg[16]),
    .Y(areg_16_bF$buf2)
);

BUFX2 BUFX2_insert441 (
    .A(areg[16]),
    .Y(areg_16_bF$buf3)
);

BUFX2 BUFX2_insert440 (
    .A(areg[16]),
    .Y(areg_16_bF$buf4)
);

BUFX2 BUFX2_insert439 (
    .A(areg[16]),
    .Y(areg_16_bF$buf5)
);

BUFX2 BUFX2_insert438 (
    .A(_4541_),
    .Y(_4541__bF$buf0)
);

BUFX2 BUFX2_insert437 (
    .A(_4541_),
    .Y(_4541__bF$buf1)
);

BUFX2 BUFX2_insert436 (
    .A(_4541_),
    .Y(_4541__bF$buf2)
);

BUFX2 BUFX2_insert435 (
    .A(_4541_),
    .Y(_4541__bF$buf3)
);

BUFX2 BUFX2_insert434 (
    .A(_4541_),
    .Y(_4541__bF$buf4)
);

BUFX2 BUFX2_insert433 (
    .A(_2586_),
    .Y(_2586__bF$buf0)
);

BUFX2 BUFX2_insert432 (
    .A(_2586_),
    .Y(_2586__bF$buf1)
);

BUFX2 BUFX2_insert431 (
    .A(_2586_),
    .Y(_2586__bF$buf2)
);

BUFX2 BUFX2_insert430 (
    .A(_2586_),
    .Y(_2586__bF$buf3)
);

BUFX2 BUFX2_insert429 (
    .A(_2586_),
    .Y(_2586__bF$buf4)
);

BUFX2 BUFX2_insert428 (
    .A(breg[29]),
    .Y(breg_29_bF$buf0)
);

BUFX2 BUFX2_insert427 (
    .A(breg[29]),
    .Y(breg_29_bF$buf1)
);

BUFX2 BUFX2_insert426 (
    .A(breg[29]),
    .Y(breg_29_bF$buf2)
);

BUFX2 BUFX2_insert425 (
    .A(breg[29]),
    .Y(breg_29_bF$buf3)
);

BUFX2 BUFX2_insert424 (
    .A(breg[29]),
    .Y(breg_29_bF$buf4)
);

BUFX2 BUFX2_insert423 (
    .A(areg[2]),
    .Y(areg_2_bF$buf0)
);

BUFX2 BUFX2_insert422 (
    .A(areg[2]),
    .Y(areg_2_bF$buf1)
);

BUFX2 BUFX2_insert421 (
    .A(areg[2]),
    .Y(areg_2_bF$buf2)
);

BUFX2 BUFX2_insert420 (
    .A(areg[2]),
    .Y(areg_2_bF$buf3)
);

BUFX2 BUFX2_insert419 (
    .A(areg[2]),
    .Y(areg_2_bF$buf4)
);

BUFX2 BUFX2_insert418 (
    .A(_7225_),
    .Y(_7225__bF$buf0)
);

BUFX2 BUFX2_insert417 (
    .A(_7225_),
    .Y(_7225__bF$buf1)
);

BUFX2 BUFX2_insert416 (
    .A(_7225_),
    .Y(_7225__bF$buf2)
);

BUFX2 BUFX2_insert415 (
    .A(_7225_),
    .Y(_7225__bF$buf3)
);

BUFX2 BUFX2_insert414 (
    .A(_7225_),
    .Y(_7225__bF$buf4)
);

BUFX2 BUFX2_insert413 (
    .A(_2551_),
    .Y(_2551__bF$buf0)
);

BUFX2 BUFX2_insert412 (
    .A(_2551_),
    .Y(_2551__bF$buf1)
);

BUFX2 BUFX2_insert411 (
    .A(_2551_),
    .Y(_2551__bF$buf2)
);

BUFX2 BUFX2_insert410 (
    .A(_2551_),
    .Y(_2551__bF$buf3)
);

BUFX2 BUFX2_insert409 (
    .A(areg[19]),
    .Y(areg_19_bF$buf0)
);

BUFX2 BUFX2_insert408 (
    .A(areg[19]),
    .Y(areg_19_bF$buf1)
);

BUFX2 BUFX2_insert407 (
    .A(areg[19]),
    .Y(areg_19_bF$buf2)
);

BUFX2 BUFX2_insert406 (
    .A(areg[19]),
    .Y(areg_19_bF$buf3)
);

BUFX2 BUFX2_insert405 (
    .A(areg[19]),
    .Y(areg_19_bF$buf4)
);

BUFX2 BUFX2_insert404 (
    .A(areg[19]),
    .Y(areg_19_bF$buf5)
);

BUFX2 BUFX2_insert403 (
    .A(areg[22]),
    .Y(areg_22_bF$buf0)
);

BUFX2 BUFX2_insert402 (
    .A(areg[22]),
    .Y(areg_22_bF$buf1)
);

BUFX2 BUFX2_insert401 (
    .A(areg[22]),
    .Y(areg_22_bF$buf2)
);

BUFX2 BUFX2_insert400 (
    .A(areg[22]),
    .Y(areg_22_bF$buf3)
);

BUFX2 BUFX2_insert399 (
    .A(areg[22]),
    .Y(areg_22_bF$buf4)
);

BUFX2 BUFX2_insert398 (
    .A(areg[5]),
    .Y(areg_5_bF$buf0)
);

BUFX2 BUFX2_insert397 (
    .A(areg[5]),
    .Y(areg_5_bF$buf1)
);

BUFX2 BUFX2_insert396 (
    .A(areg[5]),
    .Y(areg_5_bF$buf2)
);

BUFX2 BUFX2_insert395 (
    .A(areg[5]),
    .Y(areg_5_bF$buf3)
);

BUFX2 BUFX2_insert394 (
    .A(areg[5]),
    .Y(areg_5_bF$buf4)
);

BUFX2 BUFX2_insert393 (
    .A(areg[25]),
    .Y(areg_25_bF$buf0)
);

BUFX2 BUFX2_insert392 (
    .A(areg[25]),
    .Y(areg_25_bF$buf1)
);

BUFX2 BUFX2_insert391 (
    .A(areg[25]),
    .Y(areg_25_bF$buf2)
);

BUFX2 BUFX2_insert390 (
    .A(areg[25]),
    .Y(areg_25_bF$buf3)
);

BUFX2 BUFX2_insert389 (
    .A(areg[25]),
    .Y(areg_25_bF$buf4)
);

BUFX2 BUFX2_insert388 (
    .A(areg[8]),
    .Y(areg_8_bF$buf0)
);

BUFX2 BUFX2_insert387 (
    .A(areg[8]),
    .Y(areg_8_bF$buf1)
);

BUFX2 BUFX2_insert386 (
    .A(areg[8]),
    .Y(areg_8_bF$buf2)
);

BUFX2 BUFX2_insert385 (
    .A(areg[8]),
    .Y(areg_8_bF$buf3)
);

BUFX2 BUFX2_insert384 (
    .A(areg[8]),
    .Y(areg_8_bF$buf4)
);

BUFX2 BUFX2_insert383 (
    .A(_2519_),
    .Y(_2519__bF$buf0)
);

BUFX2 BUFX2_insert382 (
    .A(_2519_),
    .Y(_2519__bF$buf1)
);

BUFX2 BUFX2_insert381 (
    .A(_2519_),
    .Y(_2519__bF$buf2)
);

BUFX2 BUFX2_insert380 (
    .A(_2519_),
    .Y(_2519__bF$buf3)
);

BUFX2 BUFX2_insert379 (
    .A(_2560_),
    .Y(_2560__bF$buf0)
);

BUFX2 BUFX2_insert378 (
    .A(_2560_),
    .Y(_2560__bF$buf1)
);

BUFX2 BUFX2_insert377 (
    .A(_2560_),
    .Y(_2560__bF$buf2)
);

BUFX2 BUFX2_insert376 (
    .A(_2560_),
    .Y(_2560__bF$buf3)
);

BUFX2 BUFX2_insert375 (
    .A(_2560_),
    .Y(_2560__bF$buf4)
);

BUFX2 BUFX2_insert374 (
    .A(areg[28]),
    .Y(areg_28_bF$buf0)
);

BUFX2 BUFX2_insert373 (
    .A(areg[28]),
    .Y(areg_28_bF$buf1)
);

BUFX2 BUFX2_insert372 (
    .A(areg[28]),
    .Y(areg_28_bF$buf2)
);

BUFX2 BUFX2_insert371 (
    .A(areg[28]),
    .Y(areg_28_bF$buf3)
);

BUFX2 BUFX2_insert370 (
    .A(areg[28]),
    .Y(areg_28_bF$buf4)
);

BUFX2 BUFX2_insert369 (
    .A(areg[28]),
    .Y(areg_28_bF$buf5)
);

BUFX2 BUFX2_insert368 (
    .A(areg[31]),
    .Y(areg_31_bF$buf0)
);

BUFX2 BUFX2_insert367 (
    .A(areg[31]),
    .Y(areg_31_bF$buf1)
);

BUFX2 BUFX2_insert366 (
    .A(areg[31]),
    .Y(areg_31_bF$buf2)
);

BUFX2 BUFX2_insert365 (
    .A(areg[31]),
    .Y(areg_31_bF$buf3)
);

BUFX2 BUFX2_insert364 (
    .A(areg[31]),
    .Y(areg_31_bF$buf4)
);

BUFX2 BUFX2_insert363 (
    .A(breg[0]),
    .Y(breg_0_bF$buf0)
);

BUFX2 BUFX2_insert362 (
    .A(breg[0]),
    .Y(breg_0_bF$buf1)
);

BUFX2 BUFX2_insert361 (
    .A(breg[0]),
    .Y(breg_0_bF$buf2)
);

BUFX2 BUFX2_insert360 (
    .A(breg[0]),
    .Y(breg_0_bF$buf3)
);

BUFX2 BUFX2_insert359 (
    .A(breg[0]),
    .Y(breg_0_bF$buf4)
);

BUFX2 BUFX2_insert358 (
    .A(breg[0]),
    .Y(breg_0_bF$buf5)
);

BUFX2 BUFX2_insert357 (
    .A(breg[0]),
    .Y(breg_0_bF$buf6)
);

BUFX2 BUFX2_insert356 (
    .A(breg[12]),
    .Y(breg_12_bF$buf0)
);

BUFX2 BUFX2_insert355 (
    .A(breg[12]),
    .Y(breg_12_bF$buf1)
);

BUFX2 BUFX2_insert354 (
    .A(breg[12]),
    .Y(breg_12_bF$buf2)
);

BUFX2 BUFX2_insert353 (
    .A(breg[12]),
    .Y(breg_12_bF$buf3)
);

BUFX2 BUFX2_insert352 (
    .A(breg[12]),
    .Y(breg_12_bF$buf4)
);

BUFX2 BUFX2_insert351 (
    .A(_9104_),
    .Y(_9104__bF$buf0)
);

BUFX2 BUFX2_insert350 (
    .A(_9104_),
    .Y(_9104__bF$buf1)
);

BUFX2 BUFX2_insert349 (
    .A(_9104_),
    .Y(_9104__bF$buf2)
);

BUFX2 BUFX2_insert348 (
    .A(_9104_),
    .Y(_9104__bF$buf3)
);

BUFX2 BUFX2_insert347 (
    .A(breg[3]),
    .Y(breg_3_bF$buf0)
);

BUFX2 BUFX2_insert346 (
    .A(breg[3]),
    .Y(breg_3_bF$buf1)
);

BUFX2 BUFX2_insert345 (
    .A(breg[3]),
    .Y(breg_3_bF$buf2)
);

BUFX2 BUFX2_insert344 (
    .A(breg[3]),
    .Y(breg_3_bF$buf3)
);

BUFX2 BUFX2_insert343 (
    .A(breg[3]),
    .Y(breg_3_bF$buf4)
);

BUFX2 BUFX2_insert342 (
    .A(breg[3]),
    .Y(breg_3_bF$buf5)
);

BUFX2 BUFX2_insert341 (
    .A(breg[15]),
    .Y(breg_15_bF$buf0)
);

BUFX2 BUFX2_insert340 (
    .A(breg[15]),
    .Y(breg_15_bF$buf1)
);

BUFX2 BUFX2_insert339 (
    .A(breg[15]),
    .Y(breg_15_bF$buf2)
);

BUFX2 BUFX2_insert338 (
    .A(breg[15]),
    .Y(breg_15_bF$buf3)
);

BUFX2 BUFX2_insert337 (
    .A(breg[15]),
    .Y(breg_15_bF$buf4)
);

BUFX2 BUFX2_insert336 (
    .A(breg[15]),
    .Y(breg_15_bF$buf5)
);

BUFX2 BUFX2_insert335 (
    .A(_2287_),
    .Y(_2287__bF$buf0)
);

BUFX2 BUFX2_insert334 (
    .A(_2287_),
    .Y(_2287__bF$buf1)
);

BUFX2 BUFX2_insert333 (
    .A(_2287_),
    .Y(_2287__bF$buf2)
);

BUFX2 BUFX2_insert332 (
    .A(_2287_),
    .Y(_2287__bF$buf3)
);

BUFX2 BUFX2_insert331 (
    .A(breg[6]),
    .Y(breg_6_bF$buf0)
);

BUFX2 BUFX2_insert330 (
    .A(breg[6]),
    .Y(breg_6_bF$buf1)
);

BUFX2 BUFX2_insert329 (
    .A(breg[6]),
    .Y(breg_6_bF$buf2)
);

BUFX2 BUFX2_insert328 (
    .A(breg[6]),
    .Y(breg_6_bF$buf3)
);

BUFX2 BUFX2_insert327 (
    .A(breg[6]),
    .Y(breg_6_bF$buf4)
);

BUFX2 BUFX2_insert326 (
    .A(breg[6]),
    .Y(breg_6_bF$buf5)
);

BUFX2 BUFX2_insert325 (
    .A(_2669_),
    .Y(_2669__bF$buf0)
);

BUFX2 BUFX2_insert324 (
    .A(_2669_),
    .Y(_2669__bF$buf1)
);

BUFX2 BUFX2_insert323 (
    .A(_2669_),
    .Y(_2669__bF$buf2)
);

BUFX2 BUFX2_insert322 (
    .A(_2669_),
    .Y(_2669__bF$buf3)
);

BUFX2 BUFX2_insert321 (
    .A(_5315_),
    .Y(_5315__bF$buf0)
);

BUFX2 BUFX2_insert320 (
    .A(_5315_),
    .Y(_5315__bF$buf1)
);

BUFX2 BUFX2_insert319 (
    .A(_5315_),
    .Y(_5315__bF$buf2)
);

BUFX2 BUFX2_insert318 (
    .A(_5315_),
    .Y(_5315__bF$buf3)
);

BUFX2 BUFX2_insert317 (
    .A(_5315_),
    .Y(_5315__bF$buf4)
);

BUFX2 BUFX2_insert316 (
    .A(_6044_),
    .Y(_6044__bF$buf0)
);

BUFX2 BUFX2_insert315 (
    .A(_6044_),
    .Y(_6044__bF$buf1)
);

BUFX2 BUFX2_insert314 (
    .A(_6044_),
    .Y(_6044__bF$buf2)
);

BUFX2 BUFX2_insert313 (
    .A(_6044_),
    .Y(_6044__bF$buf3)
);

BUFX2 BUFX2_insert312 (
    .A(_6044_),
    .Y(_6044__bF$buf4)
);

BUFX2 BUFX2_insert311 (
    .A(_6044_),
    .Y(_6044__bF$buf5)
);

BUFX2 BUFX2_insert310 (
    .A(breg[18]),
    .Y(breg_18_bF$buf0)
);

BUFX2 BUFX2_insert309 (
    .A(breg[18]),
    .Y(breg_18_bF$buf1)
);

BUFX2 BUFX2_insert308 (
    .A(breg[18]),
    .Y(breg_18_bF$buf2)
);

BUFX2 BUFX2_insert307 (
    .A(breg[18]),
    .Y(breg_18_bF$buf3)
);

BUFX2 BUFX2_insert306 (
    .A(breg[18]),
    .Y(breg_18_bF$buf4)
);

BUFX2 BUFX2_insert305 (
    .A(breg[18]),
    .Y(breg_18_bF$buf5)
);

BUFX2 BUFX2_insert304 (
    .A(_2825_),
    .Y(_2825__bF$buf0)
);

BUFX2 BUFX2_insert303 (
    .A(_2825_),
    .Y(_2825__bF$buf1)
);

BUFX2 BUFX2_insert302 (
    .A(_2825_),
    .Y(_2825__bF$buf2)
);

BUFX2 BUFX2_insert301 (
    .A(_2825_),
    .Y(_2825__bF$buf3)
);

BUFX2 BUFX2_insert300 (
    .A(_2825_),
    .Y(_2825__bF$buf4)
);

BUFX2 BUFX2_insert299 (
    .A(breg[21]),
    .Y(breg_21_bF$buf0)
);

BUFX2 BUFX2_insert298 (
    .A(breg[21]),
    .Y(breg_21_bF$buf1)
);

BUFX2 BUFX2_insert297 (
    .A(breg[21]),
    .Y(breg_21_bF$buf2)
);

BUFX2 BUFX2_insert296 (
    .A(breg[21]),
    .Y(breg_21_bF$buf3)
);

BUFX2 BUFX2_insert295 (
    .A(breg[21]),
    .Y(breg_21_bF$buf4)
);

BUFX2 BUFX2_insert294 (
    .A(breg[9]),
    .Y(breg_9_bF$buf0)
);

BUFX2 BUFX2_insert293 (
    .A(breg[9]),
    .Y(breg_9_bF$buf1)
);

BUFX2 BUFX2_insert292 (
    .A(breg[9]),
    .Y(breg_9_bF$buf2)
);

BUFX2 BUFX2_insert291 (
    .A(breg[9]),
    .Y(breg_9_bF$buf3)
);

BUFX2 BUFX2_insert290 (
    .A(breg[9]),
    .Y(breg_9_bF$buf4)
);

BUFX2 BUFX2_insert289 (
    .A(breg[9]),
    .Y(breg_9_bF$buf5)
);

BUFX2 BUFX2_insert288 (
    .A(_5453_),
    .Y(_5453__bF$buf0)
);

BUFX2 BUFX2_insert287 (
    .A(_5453_),
    .Y(_5453__bF$buf1)
);

BUFX2 BUFX2_insert286 (
    .A(_5453_),
    .Y(_5453__bF$buf2)
);

BUFX2 BUFX2_insert285 (
    .A(_5453_),
    .Y(_5453__bF$buf3)
);

BUFX2 BUFX2_insert284 (
    .A(_5453_),
    .Y(_5453__bF$buf4)
);

BUFX2 BUFX2_insert283 (
    .A(_5453_),
    .Y(_5453__bF$buf5)
);

BUFX2 BUFX2_insert282 (
    .A(areg[11]),
    .Y(areg_11_bF$buf0)
);

BUFX2 BUFX2_insert281 (
    .A(areg[11]),
    .Y(areg_11_bF$buf1)
);

BUFX2 BUFX2_insert280 (
    .A(areg[11]),
    .Y(areg_11_bF$buf2)
);

BUFX2 BUFX2_insert279 (
    .A(areg[11]),
    .Y(areg_11_bF$buf3)
);

BUFX2 BUFX2_insert278 (
    .A(areg[11]),
    .Y(areg_11_bF$buf4)
);

BUFX2 BUFX2_insert277 (
    .A(_6050_),
    .Y(_6050__bF$buf0)
);

BUFX2 BUFX2_insert276 (
    .A(_6050_),
    .Y(_6050__bF$buf1)
);

BUFX2 BUFX2_insert275 (
    .A(_6050_),
    .Y(_6050__bF$buf2)
);

BUFX2 BUFX2_insert274 (
    .A(_6050_),
    .Y(_6050__bF$buf3)
);

BUFX2 BUFX2_insert273 (
    .A(_7217_),
    .Y(_7217__bF$buf0)
);

BUFX2 BUFX2_insert272 (
    .A(_7217_),
    .Y(_7217__bF$buf1)
);

BUFX2 BUFX2_insert271 (
    .A(_7217_),
    .Y(_7217__bF$buf2)
);

BUFX2 BUFX2_insert270 (
    .A(_7217_),
    .Y(_7217__bF$buf3)
);

BUFX2 BUFX2_insert269 (
    .A(_7217_),
    .Y(_7217__bF$buf4)
);

BUFX2 BUFX2_insert268 (
    .A(breg[24]),
    .Y(breg_24_bF$buf0)
);

BUFX2 BUFX2_insert267 (
    .A(breg[24]),
    .Y(breg_24_bF$buf1)
);

BUFX2 BUFX2_insert266 (
    .A(breg[24]),
    .Y(breg_24_bF$buf2)
);

BUFX2 BUFX2_insert265 (
    .A(breg[24]),
    .Y(breg_24_bF$buf3)
);

BUFX2 BUFX2_insert264 (
    .A(breg[24]),
    .Y(breg_24_bF$buf4)
);

BUFX2 BUFX2_insert263 (
    .A(breg[24]),
    .Y(breg_24_bF$buf5)
);

BUFX2 BUFX2_insert262 (
    .A(_6300_),
    .Y(_6300__bF$buf0)
);

BUFX2 BUFX2_insert261 (
    .A(_6300_),
    .Y(_6300__bF$buf1)
);

BUFX2 BUFX2_insert260 (
    .A(_6300_),
    .Y(_6300__bF$buf2)
);

BUFX2 BUFX2_insert259 (
    .A(_6300_),
    .Y(_6300__bF$buf3)
);

BUFX2 BUFX2_insert258 (
    .A(_4116_),
    .Y(_4116__bF$buf0)
);

BUFX2 BUFX2_insert257 (
    .A(_4116_),
    .Y(_4116__bF$buf1)
);

BUFX2 BUFX2_insert256 (
    .A(_4116_),
    .Y(_4116__bF$buf2)
);

BUFX2 BUFX2_insert255 (
    .A(_4116_),
    .Y(_4116__bF$buf3)
);

BUFX2 BUFX2_insert254 (
    .A(_4116_),
    .Y(_4116__bF$buf4)
);

BUFX2 BUFX2_insert253 (
    .A(areg[14]),
    .Y(areg_14_bF$buf0)
);

BUFX2 BUFX2_insert252 (
    .A(areg[14]),
    .Y(areg_14_bF$buf1)
);

BUFX2 BUFX2_insert251 (
    .A(areg[14]),
    .Y(areg_14_bF$buf2)
);

BUFX2 BUFX2_insert250 (
    .A(areg[14]),
    .Y(areg_14_bF$buf3)
);

BUFX2 BUFX2_insert249 (
    .A(areg[14]),
    .Y(areg_14_bF$buf4)
);

BUFX2 BUFX2_insert248 (
    .A(breg[27]),
    .Y(breg_27_bF$buf0)
);

BUFX2 BUFX2_insert247 (
    .A(breg[27]),
    .Y(breg_27_bF$buf1)
);

BUFX2 BUFX2_insert246 (
    .A(breg[27]),
    .Y(breg_27_bF$buf2)
);

BUFX2 BUFX2_insert245 (
    .A(breg[27]),
    .Y(breg_27_bF$buf3)
);

BUFX2 BUFX2_insert244 (
    .A(breg[27]),
    .Y(breg_27_bF$buf4)
);

BUFX2 BUFX2_insert243 (
    .A(breg[27]),
    .Y(breg_27_bF$buf5)
);

BUFX2 BUFX2_insert242 (
    .A(areg[17]),
    .Y(areg_17_bF$buf0)
);

BUFX2 BUFX2_insert241 (
    .A(areg[17]),
    .Y(areg_17_bF$buf1)
);

BUFX2 BUFX2_insert240 (
    .A(areg[17]),
    .Y(areg_17_bF$buf2)
);

BUFX2 BUFX2_insert239 (
    .A(areg[17]),
    .Y(areg_17_bF$buf3)
);

BUFX2 BUFX2_insert238 (
    .A(areg[17]),
    .Y(areg_17_bF$buf4)
);

BUFX2 BUFX2_insert237 (
    .A(areg[17]),
    .Y(areg_17_bF$buf5)
);

BUFX2 BUFX2_insert236 (
    .A(areg[20]),
    .Y(areg_20_bF$buf0)
);

BUFX2 BUFX2_insert235 (
    .A(areg[20]),
    .Y(areg_20_bF$buf1)
);

BUFX2 BUFX2_insert234 (
    .A(areg[20]),
    .Y(areg_20_bF$buf2)
);

BUFX2 BUFX2_insert233 (
    .A(areg[20]),
    .Y(areg_20_bF$buf3)
);

BUFX2 BUFX2_insert232 (
    .A(areg[20]),
    .Y(areg_20_bF$buf4)
);

BUFX2 BUFX2_insert231 (
    .A(areg[3]),
    .Y(areg_3_bF$buf0)
);

BUFX2 BUFX2_insert230 (
    .A(areg[3]),
    .Y(areg_3_bF$buf1)
);

BUFX2 BUFX2_insert229 (
    .A(areg[3]),
    .Y(areg_3_bF$buf2)
);

BUFX2 BUFX2_insert228 (
    .A(areg[3]),
    .Y(areg_3_bF$buf3)
);

BUFX2 BUFX2_insert227 (
    .A(areg[3]),
    .Y(areg_3_bF$buf4)
);

BUFX2 BUFX2_insert226 (
    .A(_3146_),
    .Y(_3146__bF$buf0)
);

BUFX2 BUFX2_insert225 (
    .A(_3146_),
    .Y(_3146__bF$buf1)
);

BUFX2 BUFX2_insert224 (
    .A(_3146_),
    .Y(_3146__bF$buf2)
);

BUFX2 BUFX2_insert223 (
    .A(_3146_),
    .Y(_3146__bF$buf3)
);

BUFX2 BUFX2_insert222 (
    .A(areg[23]),
    .Y(areg_23_bF$buf0)
);

BUFX2 BUFX2_insert221 (
    .A(areg[23]),
    .Y(areg_23_bF$buf1)
);

BUFX2 BUFX2_insert220 (
    .A(areg[23]),
    .Y(areg_23_bF$buf2)
);

BUFX2 BUFX2_insert219 (
    .A(areg[23]),
    .Y(areg_23_bF$buf3)
);

BUFX2 BUFX2_insert218 (
    .A(areg[23]),
    .Y(areg_23_bF$buf4)
);

BUFX2 BUFX2_insert217 (
    .A(areg[6]),
    .Y(areg_6_bF$buf0)
);

BUFX2 BUFX2_insert216 (
    .A(areg[6]),
    .Y(areg_6_bF$buf1)
);

BUFX2 BUFX2_insert215 (
    .A(areg[6]),
    .Y(areg_6_bF$buf2)
);

BUFX2 BUFX2_insert214 (
    .A(areg[6]),
    .Y(areg_6_bF$buf3)
);

BUFX2 BUFX2_insert213 (
    .A(areg[6]),
    .Y(areg_6_bF$buf4)
);

BUFX2 BUFX2_insert212 (
    .A(areg[26]),
    .Y(areg_26_bF$buf0)
);

BUFX2 BUFX2_insert211 (
    .A(areg[26]),
    .Y(areg_26_bF$buf1)
);

BUFX2 BUFX2_insert210 (
    .A(areg[26]),
    .Y(areg_26_bF$buf2)
);

BUFX2 BUFX2_insert209 (
    .A(areg[26]),
    .Y(areg_26_bF$buf3)
);

BUFX2 BUFX2_insert208 (
    .A(areg[26]),
    .Y(areg_26_bF$buf4)
);

BUFX2 BUFX2_insert207 (
    .A(_7100_),
    .Y(_7100__bF$buf0)
);

BUFX2 BUFX2_insert206 (
    .A(_7100_),
    .Y(_7100__bF$buf1)
);

BUFX2 BUFX2_insert205 (
    .A(_7100_),
    .Y(_7100__bF$buf2)
);

BUFX2 BUFX2_insert204 (
    .A(_7100_),
    .Y(_7100__bF$buf3)
);

BUFX2 BUFX2_insert203 (
    .A(_7520_),
    .Y(_7520__bF$buf0)
);

BUFX2 BUFX2_insert202 (
    .A(_7520_),
    .Y(_7520__bF$buf1)
);

BUFX2 BUFX2_insert201 (
    .A(_7520_),
    .Y(_7520__bF$buf2)
);

BUFX2 BUFX2_insert200 (
    .A(_7520_),
    .Y(_7520__bF$buf3)
);

BUFX2 BUFX2_insert199 (
    .A(_7711_),
    .Y(_7711__bF$buf0)
);

BUFX2 BUFX2_insert198 (
    .A(_7711_),
    .Y(_7711__bF$buf1)
);

BUFX2 BUFX2_insert197 (
    .A(_7711_),
    .Y(_7711__bF$buf2)
);

BUFX2 BUFX2_insert196 (
    .A(_7711_),
    .Y(_7711__bF$buf3)
);

BUFX2 BUFX2_insert195 (
    .A(_3402_),
    .Y(_3402__bF$buf0)
);

BUFX2 BUFX2_insert194 (
    .A(_3402_),
    .Y(_3402__bF$buf1)
);

BUFX2 BUFX2_insert193 (
    .A(_3402_),
    .Y(_3402__bF$buf2)
);

BUFX2 BUFX2_insert192 (
    .A(_3402_),
    .Y(_3402__bF$buf3)
);

BUFX2 BUFX2_insert191 (
    .A(_4551_),
    .Y(_4551__bF$buf0)
);

BUFX2 BUFX2_insert190 (
    .A(_4551_),
    .Y(_4551__bF$buf1)
);

BUFX2 BUFX2_insert189 (
    .A(_4551_),
    .Y(_4551__bF$buf2)
);

BUFX2 BUFX2_insert188 (
    .A(_4551_),
    .Y(_4551__bF$buf3)
);

BUFX2 BUFX2_insert187 (
    .A(_4551_),
    .Y(_4551__bF$buf4)
);

BUFX2 BUFX2_insert186 (
    .A(areg[9]),
    .Y(areg_9_bF$buf0)
);

BUFX2 BUFX2_insert185 (
    .A(areg[9]),
    .Y(areg_9_bF$buf1)
);

BUFX2 BUFX2_insert184 (
    .A(areg[9]),
    .Y(areg_9_bF$buf2)
);

BUFX2 BUFX2_insert183 (
    .A(areg[9]),
    .Y(areg_9_bF$buf3)
);

BUFX2 BUFX2_insert182 (
    .A(areg[9]),
    .Y(areg_9_bF$buf4)
);

BUFX2 BUFX2_insert181 (
    .A(_549_),
    .Y(_549__bF$buf0)
);

BUFX2 BUFX2_insert180 (
    .A(_549_),
    .Y(_549__bF$buf1)
);

BUFX2 BUFX2_insert179 (
    .A(_549_),
    .Y(_549__bF$buf2)
);

BUFX2 BUFX2_insert178 (
    .A(_549_),
    .Y(_549__bF$buf3)
);

BUFX2 BUFX2_insert177 (
    .A(_549_),
    .Y(_549__bF$buf4)
);

BUFX2 BUFX2_insert176 (
    .A(_6582_),
    .Y(_6582__bF$buf0)
);

BUFX2 BUFX2_insert175 (
    .A(_6582_),
    .Y(_6582__bF$buf1)
);

BUFX2 BUFX2_insert174 (
    .A(_6582_),
    .Y(_6582__bF$buf2)
);

BUFX2 BUFX2_insert173 (
    .A(_6582_),
    .Y(_6582__bF$buf3)
);

BUFX2 BUFX2_insert172 (
    .A(_2884_),
    .Y(_2884__bF$buf0)
);

BUFX2 BUFX2_insert171 (
    .A(_2884_),
    .Y(_2884__bF$buf1)
);

BUFX2 BUFX2_insert170 (
    .A(_2884_),
    .Y(_2884__bF$buf2)
);

BUFX2 BUFX2_insert169 (
    .A(_2884_),
    .Y(_2884__bF$buf3)
);

BUFX2 BUFX2_insert168 (
    .A(areg[29]),
    .Y(areg_29_bF$buf0)
);

BUFX2 BUFX2_insert167 (
    .A(areg[29]),
    .Y(areg_29_bF$buf1)
);

BUFX2 BUFX2_insert166 (
    .A(areg[29]),
    .Y(areg_29_bF$buf2)
);

BUFX2 BUFX2_insert165 (
    .A(areg[29]),
    .Y(areg_29_bF$buf3)
);

BUFX2 BUFX2_insert164 (
    .A(areg[29]),
    .Y(areg_29_bF$buf4)
);

BUFX2 BUFX2_insert163 (
    .A(areg[29]),
    .Y(areg_29_bF$buf5)
);

BUFX2 BUFX2_insert162 (
    .A(_5668_),
    .Y(_5668__bF$buf0)
);

BUFX2 BUFX2_insert161 (
    .A(_5668_),
    .Y(_5668__bF$buf1)
);

BUFX2 BUFX2_insert160 (
    .A(_5668_),
    .Y(_5668__bF$buf2)
);

BUFX2 BUFX2_insert159 (
    .A(_5668_),
    .Y(_5668__bF$buf3)
);

BUFX2 BUFX2_insert158 (
    .A(_5668_),
    .Y(_5668__bF$buf4)
);

BUFX2 BUFX2_insert157 (
    .A(_5668_),
    .Y(_5668__bF$buf5)
);

BUFX2 BUFX2_insert156 (
    .A(breg[10]),
    .Y(breg_10_bF$buf0)
);

BUFX2 BUFX2_insert155 (
    .A(breg[10]),
    .Y(breg_10_bF$buf1)
);

BUFX2 BUFX2_insert154 (
    .A(breg[10]),
    .Y(breg_10_bF$buf2)
);

BUFX2 BUFX2_insert153 (
    .A(breg[10]),
    .Y(breg_10_bF$buf3)
);

BUFX2 BUFX2_insert152 (
    .A(breg[10]),
    .Y(breg_10_bF$buf4)
);

BUFX2 BUFX2_insert151 (
    .A(breg[10]),
    .Y(breg_10_bF$buf5)
);

BUFX2 BUFX2_insert150 (
    .A(_2376_),
    .Y(_2376__bF$buf0)
);

BUFX2 BUFX2_insert149 (
    .A(_2376_),
    .Y(_2376__bF$buf1)
);

BUFX2 BUFX2_insert148 (
    .A(_2376_),
    .Y(_2376__bF$buf2)
);

BUFX2 BUFX2_insert147 (
    .A(_2376_),
    .Y(_2376__bF$buf3)
);

BUFX2 BUFX2_insert146 (
    .A(breg[1]),
    .Y(breg_1_bF$buf0)
);

BUFX2 BUFX2_insert145 (
    .A(breg[1]),
    .Y(breg_1_bF$buf1)
);

BUFX2 BUFX2_insert144 (
    .A(breg[1]),
    .Y(breg_1_bF$buf2)
);

BUFX2 BUFX2_insert143 (
    .A(breg[1]),
    .Y(breg_1_bF$buf3)
);

BUFX2 BUFX2_insert142 (
    .A(breg[1]),
    .Y(breg_1_bF$buf4)
);

BUFX2 BUFX2_insert141 (
    .A(breg[1]),
    .Y(breg_1_bF$buf5)
);

BUFX2 BUFX2_insert140 (
    .A(breg[1]),
    .Y(breg_1_bF$buf6)
);

BUFX2 BUFX2_insert139 (
    .A(_5921_),
    .Y(_5921__bF$buf0)
);

BUFX2 BUFX2_insert138 (
    .A(_5921_),
    .Y(_5921__bF$buf1)
);

BUFX2 BUFX2_insert137 (
    .A(_5921_),
    .Y(_5921__bF$buf2)
);

BUFX2 BUFX2_insert136 (
    .A(_5921_),
    .Y(_5921__bF$buf3)
);

BUFX2 BUFX2_insert135 (
    .A(breg[13]),
    .Y(breg_13_bF$buf0)
);

BUFX2 BUFX2_insert134 (
    .A(breg[13]),
    .Y(breg_13_bF$buf1)
);

BUFX2 BUFX2_insert133 (
    .A(breg[13]),
    .Y(breg_13_bF$buf2)
);

BUFX2 BUFX2_insert132 (
    .A(breg[13]),
    .Y(breg_13_bF$buf3)
);

BUFX2 BUFX2_insert131 (
    .A(breg[13]),
    .Y(breg_13_bF$buf4)
);

BUFX2 BUFX2_insert130 (
    .A(breg[4]),
    .Y(breg_4_bF$buf0)
);

BUFX2 BUFX2_insert129 (
    .A(breg[4]),
    .Y(breg_4_bF$buf1)
);

BUFX2 BUFX2_insert128 (
    .A(breg[4]),
    .Y(breg_4_bF$buf2)
);

BUFX2 BUFX2_insert127 (
    .A(breg[4]),
    .Y(breg_4_bF$buf3)
);

BUFX2 BUFX2_insert126 (
    .A(breg[4]),
    .Y(breg_4_bF$buf4)
);

BUFX2 BUFX2_insert125 (
    .A(breg[4]),
    .Y(breg_4_bF$buf5)
);

BUFX2 BUFX2_insert124 (
    .A(_3646_),
    .Y(_3646__bF$buf0)
);

BUFX2 BUFX2_insert123 (
    .A(_3646_),
    .Y(_3646__bF$buf1)
);

BUFX2 BUFX2_insert122 (
    .A(_3646_),
    .Y(_3646__bF$buf2)
);

BUFX2 BUFX2_insert121 (
    .A(_3646_),
    .Y(_3646__bF$buf3)
);

BUFX2 BUFX2_insert120 (
    .A(breg[16]),
    .Y(breg_16_bF$buf0)
);

BUFX2 BUFX2_insert119 (
    .A(breg[16]),
    .Y(breg_16_bF$buf1)
);

BUFX2 BUFX2_insert118 (
    .A(breg[16]),
    .Y(breg_16_bF$buf2)
);

BUFX2 BUFX2_insert117 (
    .A(breg[16]),
    .Y(breg_16_bF$buf3)
);

BUFX2 BUFX2_insert116 (
    .A(breg[16]),
    .Y(breg_16_bF$buf4)
);

BUFX2 BUFX2_insert115 (
    .A(breg[16]),
    .Y(breg_16_bF$buf5)
);

BUFX2 BUFX2_insert114 (
    .A(_3781_),
    .Y(_3781__bF$buf0)
);

BUFX2 BUFX2_insert113 (
    .A(_3781_),
    .Y(_3781__bF$buf1)
);

BUFX2 BUFX2_insert112 (
    .A(_3781_),
    .Y(_3781__bF$buf2)
);

BUFX2 BUFX2_insert111 (
    .A(_3781_),
    .Y(_3781__bF$buf3)
);

BUFX2 BUFX2_insert110 (
    .A(_4434_),
    .Y(_4434__bF$buf0)
);

BUFX2 BUFX2_insert109 (
    .A(_4434_),
    .Y(_4434__bF$buf1)
);

BUFX2 BUFX2_insert108 (
    .A(_4434_),
    .Y(_4434__bF$buf2)
);

BUFX2 BUFX2_insert107 (
    .A(_4434_),
    .Y(_4434__bF$buf3)
);

BUFX2 BUFX2_insert106 (
    .A(breg[7]),
    .Y(breg_7_bF$buf0)
);

BUFX2 BUFX2_insert105 (
    .A(breg[7]),
    .Y(breg_7_bF$buf1)
);

BUFX2 BUFX2_insert104 (
    .A(breg[7]),
    .Y(breg_7_bF$buf2)
);

BUFX2 BUFX2_insert103 (
    .A(breg[7]),
    .Y(breg_7_bF$buf3)
);

BUFX2 BUFX2_insert102 (
    .A(breg[7]),
    .Y(breg_7_bF$buf4)
);

BUFX2 BUFX2_insert101 (
    .A(breg[7]),
    .Y(breg_7_bF$buf5)
);

BUFX2 BUFX2_insert100 (
    .A(breg[19]),
    .Y(breg_19_bF$buf0)
);

BUFX2 BUFX2_insert99 (
    .A(breg[19]),
    .Y(breg_19_bF$buf1)
);

BUFX2 BUFX2_insert98 (
    .A(breg[19]),
    .Y(breg_19_bF$buf2)
);

BUFX2 BUFX2_insert97 (
    .A(breg[19]),
    .Y(breg_19_bF$buf3)
);

BUFX2 BUFX2_insert96 (
    .A(breg[19]),
    .Y(breg_19_bF$buf4)
);

BUFX2 BUFX2_insert95 (
    .A(breg[19]),
    .Y(breg_19_bF$buf5)
);

CLKBUF1 CLKBUF1_insert94 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert93 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert92 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert91 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert90 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert89 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert88 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert87 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert86 (
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert85 (
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert84 (
    .A(clk),
    .Y(clk_bF$buf10)
);

BUFX2 BUFX2_insert83 (
    .A(breg[22]),
    .Y(breg_22_bF$buf0)
);

BUFX2 BUFX2_insert82 (
    .A(breg[22]),
    .Y(breg_22_bF$buf1)
);

BUFX2 BUFX2_insert81 (
    .A(breg[22]),
    .Y(breg_22_bF$buf2)
);

BUFX2 BUFX2_insert80 (
    .A(breg[22]),
    .Y(breg_22_bF$buf3)
);

BUFX2 BUFX2_insert79 (
    .A(breg[22]),
    .Y(breg_22_bF$buf4)
);

BUFX2 BUFX2_insert78 (
    .A(areg[12]),
    .Y(areg_12_bF$buf0)
);

BUFX2 BUFX2_insert77 (
    .A(areg[12]),
    .Y(areg_12_bF$buf1)
);

BUFX2 BUFX2_insert76 (
    .A(areg[12]),
    .Y(areg_12_bF$buf2)
);

BUFX2 BUFX2_insert75 (
    .A(areg[12]),
    .Y(areg_12_bF$buf3)
);

BUFX2 BUFX2_insert74 (
    .A(areg[12]),
    .Y(areg_12_bF$buf4)
);

BUFX2 BUFX2_insert73 (
    .A(_6815_),
    .Y(_6815__bF$buf0)
);

BUFX2 BUFX2_insert72 (
    .A(_6815_),
    .Y(_6815__bF$buf1)
);

BUFX2 BUFX2_insert71 (
    .A(_6815_),
    .Y(_6815__bF$buf2)
);

BUFX2 BUFX2_insert70 (
    .A(_6815_),
    .Y(_6815__bF$buf3)
);

BUFX2 BUFX2_insert69 (
    .A(_6815_),
    .Y(_6815__bF$buf4)
);

BUFX2 BUFX2_insert68 (
    .A(breg[25]),
    .Y(breg_25_bF$buf0)
);

BUFX2 BUFX2_insert67 (
    .A(breg[25]),
    .Y(breg_25_bF$buf1)
);

BUFX2 BUFX2_insert66 (
    .A(breg[25]),
    .Y(breg_25_bF$buf2)
);

BUFX2 BUFX2_insert65 (
    .A(breg[25]),
    .Y(breg_25_bF$buf3)
);

BUFX2 BUFX2_insert64 (
    .A(breg[25]),
    .Y(breg_25_bF$buf4)
);

BUFX2 BUFX2_insert63 (
    .A(breg[25]),
    .Y(breg_25_bF$buf5)
);

BUFX2 BUFX2_insert62 (
    .A(areg[15]),
    .Y(areg_15_bF$buf0)
);

BUFX2 BUFX2_insert61 (
    .A(areg[15]),
    .Y(areg_15_bF$buf1)
);

BUFX2 BUFX2_insert60 (
    .A(areg[15]),
    .Y(areg_15_bF$buf2)
);

BUFX2 BUFX2_insert59 (
    .A(areg[15]),
    .Y(areg_15_bF$buf3)
);

BUFX2 BUFX2_insert58 (
    .A(areg[15]),
    .Y(areg_15_bF$buf4)
);

BUFX2 BUFX2_insert57 (
    .A(breg[28]),
    .Y(breg_28_bF$buf0)
);

BUFX2 BUFX2_insert56 (
    .A(breg[28]),
    .Y(breg_28_bF$buf1)
);

BUFX2 BUFX2_insert55 (
    .A(breg[28]),
    .Y(breg_28_bF$buf2)
);

BUFX2 BUFX2_insert54 (
    .A(breg[28]),
    .Y(breg_28_bF$buf3)
);

BUFX2 BUFX2_insert53 (
    .A(breg[28]),
    .Y(breg_28_bF$buf4)
);

BUFX2 BUFX2_insert52 (
    .A(breg[28]),
    .Y(breg_28_bF$buf5)
);

BUFX2 BUFX2_insert51 (
    .A(areg[1]),
    .Y(areg_1_bF$buf0)
);

BUFX2 BUFX2_insert50 (
    .A(areg[1]),
    .Y(areg_1_bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .A(areg[1]),
    .Y(areg_1_bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .A(areg[1]),
    .Y(areg_1_bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .A(areg[1]),
    .Y(areg_1_bF$buf4)
);

BUFX2 BUFX2_insert46 (
    .A(areg[18]),
    .Y(areg_18_bF$buf0)
);

BUFX2 BUFX2_insert45 (
    .A(areg[18]),
    .Y(areg_18_bF$buf1)
);

BUFX2 BUFX2_insert44 (
    .A(areg[18]),
    .Y(areg_18_bF$buf2)
);

BUFX2 BUFX2_insert43 (
    .A(areg[18]),
    .Y(areg_18_bF$buf3)
);

BUFX2 BUFX2_insert42 (
    .A(areg[18]),
    .Y(areg_18_bF$buf4)
);

BUFX2 BUFX2_insert41 (
    .A(areg[18]),
    .Y(areg_18_bF$buf5)
);

BUFX2 BUFX2_insert40 (
    .A(areg[21]),
    .Y(areg_21_bF$buf0)
);

BUFX2 BUFX2_insert39 (
    .A(areg[21]),
    .Y(areg_21_bF$buf1)
);

BUFX2 BUFX2_insert38 (
    .A(areg[21]),
    .Y(areg_21_bF$buf2)
);

BUFX2 BUFX2_insert37 (
    .A(areg[21]),
    .Y(areg_21_bF$buf3)
);

BUFX2 BUFX2_insert36 (
    .A(areg[21]),
    .Y(areg_21_bF$buf4)
);

BUFX2 BUFX2_insert35 (
    .A(areg[4]),
    .Y(areg_4_bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .A(areg[4]),
    .Y(areg_4_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .A(areg[4]),
    .Y(areg_4_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .A(areg[4]),
    .Y(areg_4_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .A(areg[4]),
    .Y(areg_4_bF$buf4)
);

BUFX2 BUFX2_insert30 (
    .A(_2362_),
    .Y(_2362__bF$buf0)
);

BUFX2 BUFX2_insert29 (
    .A(_2362_),
    .Y(_2362__bF$buf1)
);

BUFX2 BUFX2_insert28 (
    .A(_2362_),
    .Y(_2362__bF$buf2)
);

BUFX2 BUFX2_insert27 (
    .A(_2362_),
    .Y(_2362__bF$buf3)
);

BUFX2 BUFX2_insert26 (
    .A(_2362_),
    .Y(_2362__bF$buf4)
);

BUFX2 BUFX2_insert25 (
    .A(_2362_),
    .Y(_2362__bF$buf5)
);

BUFX2 BUFX2_insert24 (
    .A(_3529_),
    .Y(_3529__bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(_3529_),
    .Y(_3529__bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(_3529_),
    .Y(_3529__bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(_3529_),
    .Y(_3529__bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(_3529_),
    .Y(_3529__bF$buf4)
);

BUFX2 BUFX2_insert19 (
    .A(_4258_),
    .Y(_4258__bF$buf0)
);

BUFX2 BUFX2_insert18 (
    .A(_4258_),
    .Y(_4258__bF$buf1)
);

BUFX2 BUFX2_insert17 (
    .A(_4258_),
    .Y(_4258__bF$buf2)
);

BUFX2 BUFX2_insert16 (
    .A(_4258_),
    .Y(_4258__bF$buf3)
);

BUFX2 BUFX2_insert15 (
    .A(areg[24]),
    .Y(areg_24_bF$buf0)
);

BUFX2 BUFX2_insert14 (
    .A(areg[24]),
    .Y(areg_24_bF$buf1)
);

BUFX2 BUFX2_insert13 (
    .A(areg[24]),
    .Y(areg_24_bF$buf2)
);

BUFX2 BUFX2_insert12 (
    .A(areg[24]),
    .Y(areg_24_bF$buf3)
);

BUFX2 BUFX2_insert11 (
    .A(areg[24]),
    .Y(areg_24_bF$buf4)
);

BUFX2 BUFX2_insert10 (
    .A(areg[7]),
    .Y(areg_7_bF$buf0)
);

BUFX2 BUFX2_insert9 (
    .A(areg[7]),
    .Y(areg_7_bF$buf1)
);

BUFX2 BUFX2_insert8 (
    .A(areg[7]),
    .Y(areg_7_bF$buf2)
);

BUFX2 BUFX2_insert7 (
    .A(areg[7]),
    .Y(areg_7_bF$buf3)
);

BUFX2 BUFX2_insert6 (
    .A(areg[7]),
    .Y(areg_7_bF$buf4)
);

BUFX2 BUFX2_insert5 (
    .A(areg[27]),
    .Y(areg_27_bF$buf0)
);

BUFX2 BUFX2_insert4 (
    .A(areg[27]),
    .Y(areg_27_bF$buf1)
);

BUFX2 BUFX2_insert3 (
    .A(areg[27]),
    .Y(areg_27_bF$buf2)
);

BUFX2 BUFX2_insert2 (
    .A(areg[27]),
    .Y(areg_27_bF$buf3)
);

BUFX2 BUFX2_insert1 (
    .A(areg[27]),
    .Y(areg_27_bF$buf4)
);

BUFX2 BUFX2_insert0 (
    .A(areg[27]),
    .Y(areg_27_bF$buf5)
);

INVX8 _11910_ (
    .A(breg_3_bF$buf5),
    .Y(_2365_)
);

INVX8 _11911_ (
    .A(areg[0]),
    .Y(_2376_)
);

NOR2X1 _11912_ (
    .A(_2365_),
    .B(_2376__bF$buf3),
    .Y(_2387_)
);

INVX1 _11913_ (
    .A(_2387_),
    .Y(_2398_)
);

NAND2X1 _11914_ (
    .A(breg_4_bF$buf5),
    .B(areg_1_bF$buf4),
    .Y(_2419_)
);

OR2X2 _11915_ (
    .A(_2398_),
    .B(_2419_),
    .Y(_2420_)
);

INVX1 _11916_ (
    .A(_2420_),
    .Y(_2431_)
);

NAND2X1 _11917_ (
    .A(breg_1_bF$buf6),
    .B(areg_2_bF$buf4),
    .Y(_2442_)
);

NAND2X1 _11918_ (
    .A(breg_0_bF$buf6),
    .B(areg_3_bF$buf4),
    .Y(_2453_)
);

NAND2X1 _11919_ (
    .A(breg_2_bF$buf4),
    .B(areg_1_bF$buf3),
    .Y(_2464_)
);

XNOR2X1 _11920_ (
    .A(_2442_),
    .B(_2453_),
    .Y(_2475_)
);

OR2X2 _11921_ (
    .A(_2475_),
    .B(_2464_),
    .Y(_2486_)
);

OAI21X1 _11922_ (
    .A(_2442_),
    .B(_2453_),
    .C(_2486_),
    .Y(_2497_)
);

INVX4 _11923_ (
    .A(breg_2_bF$buf3),
    .Y(_2508_)
);

INVX8 _11924_ (
    .A(areg_2_bF$buf3),
    .Y(_2519_)
);

NOR2X1 _11925_ (
    .A(_2508_),
    .B(_2519__bF$buf3),
    .Y(_2530_)
);

NAND2X1 _11926_ (
    .A(breg_1_bF$buf5),
    .B(areg_4_bF$buf4),
    .Y(_2540_)
);

INVX8 _11927_ (
    .A(breg_0_bF$buf5),
    .Y(_2551_)
);

INVX8 _11928_ (
    .A(areg_4_bF$buf3),
    .Y(_2562_)
);

NAND2X1 _11929_ (
    .A(breg_1_bF$buf4),
    .B(areg_3_bF$buf3),
    .Y(_2573_)
);

OAI21X1 _11930_ (
    .A(_2551__bF$buf3),
    .B(_2562__bF$buf4),
    .C(_2573_),
    .Y(_2584_)
);

OAI21X1 _11931_ (
    .A(_2453_),
    .B(_2540_),
    .C(_2584_),
    .Y(_2605_)
);

XNOR2X1 _11932_ (
    .A(_2605_),
    .B(_2530_),
    .Y(_2616_)
);

NAND2X1 _11933_ (
    .A(_2616_),
    .B(_2497_),
    .Y(_2617_)
);

INVX1 _11934_ (
    .A(_2617_),
    .Y(_2628_)
);

OR2X2 _11935_ (
    .A(_2497_),
    .B(_2616_),
    .Y(_2639_)
);

INVX1 _11936_ (
    .A(breg_4_bF$buf4),
    .Y(_2650_)
);

INVX8 _11937_ (
    .A(areg_1_bF$buf2),
    .Y(_2661_)
);

OAI22X1 _11938_ (
    .A(_2365_),
    .B(_2661_),
    .C(_2650_),
    .D(_2376__bF$buf2),
    .Y(_2672_)
);

OAI21X1 _11939_ (
    .A(_2398_),
    .B(_2419_),
    .C(_2672_),
    .Y(_2683_)
);

INVX1 _11940_ (
    .A(_2683_),
    .Y(_2694_)
);

AOI21X1 _11941_ (
    .A(_2639_),
    .B(_2694_),
    .C(_2628_),
    .Y(_2705_)
);

NAND2X1 _11942_ (
    .A(breg_5_bF$buf3),
    .B(areg[0]),
    .Y(_2716_)
);

NAND2X1 _11943_ (
    .A(areg_2_bF$buf2),
    .B(breg_3_bF$buf4),
    .Y(_2727_)
);

XOR2X1 _11944_ (
    .A(_2419_),
    .B(_2727_),
    .Y(_2738_)
);

XNOR2X1 _11945_ (
    .A(_2738_),
    .B(_2716_),
    .Y(_2749_)
);

NAND2X1 _11946_ (
    .A(breg_0_bF$buf4),
    .B(areg_4_bF$buf2),
    .Y(_2759_)
);

NOR2X1 _11947_ (
    .A(_2573_),
    .B(_2759_),
    .Y(_2770_)
);

AOI21X1 _11948_ (
    .A(_2530_),
    .B(_2584_),
    .C(_2770_),
    .Y(_2781_)
);

INVX8 _11949_ (
    .A(areg_3_bF$buf2),
    .Y(_2792_)
);

NOR2X1 _11950_ (
    .A(_2508_),
    .B(_2792_),
    .Y(_2803_)
);

NAND2X1 _11951_ (
    .A(areg_5_bF$buf4),
    .B(breg_1_bF$buf3),
    .Y(_2814_)
);

INVX8 _11952_ (
    .A(areg_5_bF$buf3),
    .Y(_2825_)
);

OAI21X1 _11953_ (
    .A(_2551__bF$buf2),
    .B(_2825__bF$buf4),
    .C(_2540_),
    .Y(_2836_)
);

OAI21X1 _11954_ (
    .A(_2759_),
    .B(_2814_),
    .C(_2836_),
    .Y(_2847_)
);

XNOR2X1 _11955_ (
    .A(_2847_),
    .B(_2803_),
    .Y(_2858_)
);

XNOR2X1 _11956_ (
    .A(_2858_),
    .B(_2781_),
    .Y(_2869_)
);

NAND2X1 _11957_ (
    .A(_2749_),
    .B(_2869_),
    .Y(_2880_)
);

INVX1 _11958_ (
    .A(_2749_),
    .Y(_2901_)
);

INVX1 _11959_ (
    .A(_2803_),
    .Y(_2902_)
);

XNOR2X1 _11960_ (
    .A(_2847_),
    .B(_2902_),
    .Y(_2913_)
);

NOR2X1 _11961_ (
    .A(_2781_),
    .B(_2913_),
    .Y(_2924_)
);

INVX1 _11962_ (
    .A(_2781_),
    .Y(_2935_)
);

NOR2X1 _11963_ (
    .A(_2935_),
    .B(_2858_),
    .Y(_2946_)
);

OAI21X1 _11964_ (
    .A(_2924_),
    .B(_2946_),
    .C(_2901_),
    .Y(_2957_)
);

NAND2X1 _11965_ (
    .A(_2957_),
    .B(_2880_),
    .Y(_2968_)
);

OR2X2 _11966_ (
    .A(_2968_),
    .B(_2705_),
    .Y(_2978_)
);

NAND2X1 _11967_ (
    .A(_2705_),
    .B(_2968_),
    .Y(_2989_)
);

NAND3X1 _11968_ (
    .A(_2431_),
    .B(_2989_),
    .C(_2978_),
    .Y(_3000_)
);

NOR2X1 _11969_ (
    .A(_2705_),
    .B(_2968_),
    .Y(_3011_)
);

AND2X2 _11970_ (
    .A(_2968_),
    .B(_2705_),
    .Y(_3022_)
);

OAI21X1 _11971_ (
    .A(_3022_),
    .B(_3011_),
    .C(_2420_),
    .Y(_3033_)
);

NAND2X1 _11972_ (
    .A(_3033_),
    .B(_3000_),
    .Y(_3044_)
);

NAND2X1 _11973_ (
    .A(breg_0_bF$buf3),
    .B(areg_1_bF$buf1),
    .Y(_3055_)
);

NOR2X1 _11974_ (
    .A(_2442_),
    .B(_3055_),
    .Y(_3066_)
);

AOI22X1 _11975_ (
    .A(breg_0_bF$buf2),
    .B(areg_2_bF$buf1),
    .C(breg_1_bF$buf2),
    .D(areg_1_bF$buf0),
    .Y(_3077_)
);

NOR2X1 _11976_ (
    .A(_3077_),
    .B(_3066_),
    .Y(_3088_)
);

NOR2X1 _11977_ (
    .A(_2508_),
    .B(_2376__bF$buf1),
    .Y(_3099_)
);

AOI21X1 _11978_ (
    .A(_3099_),
    .B(_3088_),
    .C(_3066_),
    .Y(_3110_)
);

OAI21X1 _11979_ (
    .A(_2508_),
    .B(_2661_),
    .C(_2475_),
    .Y(_3131_)
);

NAND2X1 _11980_ (
    .A(_3131_),
    .B(_2486_),
    .Y(_3142_)
);

NOR2X1 _11981_ (
    .A(_3110_),
    .B(_3142_),
    .Y(_3143_)
);

INVX2 _11982_ (
    .A(_3099_),
    .Y(_3154_)
);

OAI22X1 _11983_ (
    .A(_2442_),
    .B(_3055_),
    .C(_3154_),
    .D(_3077_),
    .Y(_3165_)
);

XNOR2X1 _11984_ (
    .A(_3142_),
    .B(_3165_),
    .Y(_3176_)
);

AOI21X1 _11985_ (
    .A(_2387_),
    .B(_3176_),
    .C(_3143_),
    .Y(_3187_)
);

XNOR2X1 _11986_ (
    .A(_2497_),
    .B(_2616_),
    .Y(_3198_)
);

XNOR2X1 _11987_ (
    .A(_3198_),
    .B(_2683_),
    .Y(_3209_)
);

INVX4 _11988_ (
    .A(breg_1_bF$buf1),
    .Y(_3220_)
);

NOR2X1 _11989_ (
    .A(_3220_),
    .B(_2376__bF$buf0),
    .Y(_3231_)
);

INVX1 _11990_ (
    .A(_3231_),
    .Y(_3241_)
);

NOR2X1 _11991_ (
    .A(_3055_),
    .B(_3241_),
    .Y(_3252_)
);

XNOR2X1 _11992_ (
    .A(_3088_),
    .B(_3154_),
    .Y(_3263_)
);

NAND2X1 _11993_ (
    .A(_3252_),
    .B(_3263_),
    .Y(_3274_)
);

XNOR2X1 _11994_ (
    .A(_3176_),
    .B(_2387_),
    .Y(_3285_)
);

NOR2X1 _11995_ (
    .A(_3274_),
    .B(_3285_),
    .Y(_3296_)
);

XOR2X1 _11996_ (
    .A(_3209_),
    .B(_3187_),
    .Y(_3307_)
);

NAND2X1 _11997_ (
    .A(_3296_),
    .B(_3307_),
    .Y(_3318_)
);

OAI21X1 _11998_ (
    .A(_3187_),
    .B(_3209_),
    .C(_3318_),
    .Y(_3329_)
);

XNOR2X1 _11999_ (
    .A(_3329_),
    .B(_3044_),
    .Y(_0_[5])
);

NOR2X1 _12000_ (
    .A(_3044_),
    .B(_3318_),
    .Y(_3350_)
);

NOR2X1 _12001_ (
    .A(_3187_),
    .B(_3209_),
    .Y(_3361_)
);

NAND3X1 _12002_ (
    .A(_3361_),
    .B(_3033_),
    .C(_3000_),
    .Y(_3372_)
);

OAI21X1 _12003_ (
    .A(_3022_),
    .B(_2420_),
    .C(_2978_),
    .Y(_3383_)
);

NAND2X1 _12004_ (
    .A(areg[0]),
    .B(breg_6_bF$buf5),
    .Y(_3394_)
);

INVX1 _12005_ (
    .A(_3394_),
    .Y(_3405_)
);

NAND3X1 _12006_ (
    .A(breg_5_bF$buf2),
    .B(areg[0]),
    .C(_2738_),
    .Y(_3416_)
);

OAI21X1 _12007_ (
    .A(_2419_),
    .B(_2727_),
    .C(_3416_),
    .Y(_3427_)
);

NOR2X1 _12008_ (
    .A(_3405_),
    .B(_3427_),
    .Y(_3438_)
);

NAND2X1 _12009_ (
    .A(_3405_),
    .B(_3427_),
    .Y(_3449_)
);

INVX2 _12010_ (
    .A(_3449_),
    .Y(_3460_)
);

OR2X2 _12011_ (
    .A(_3460_),
    .B(_3438_),
    .Y(_3471_)
);

NAND2X1 _12012_ (
    .A(_2935_),
    .B(_2858_),
    .Y(_3482_)
);

OAI21X1 _12013_ (
    .A(_2946_),
    .B(_2901_),
    .C(_3482_),
    .Y(_3493_)
);

NAND2X1 _12014_ (
    .A(areg_1_bF$buf4),
    .B(breg_5_bF$buf1),
    .Y(_3503_)
);

NAND2X1 _12015_ (
    .A(areg_2_bF$buf0),
    .B(breg_4_bF$buf3),
    .Y(_3514_)
);

NAND2X1 _12016_ (
    .A(areg_3_bF$buf1),
    .B(breg_3_bF$buf3),
    .Y(_3525_)
);

XOR2X1 _12017_ (
    .A(_3514_),
    .B(_3525_),
    .Y(_3536_)
);

XNOR2X1 _12018_ (
    .A(_3536_),
    .B(_3503_),
    .Y(_3547_)
);

INVX2 _12019_ (
    .A(_3547_),
    .Y(_3558_)
);

NAND2X1 _12020_ (
    .A(breg_0_bF$buf1),
    .B(areg_5_bF$buf2),
    .Y(_3569_)
);

NOR2X1 _12021_ (
    .A(_2540_),
    .B(_3569_),
    .Y(_3580_)
);

AOI21X1 _12022_ (
    .A(_2803_),
    .B(_2836_),
    .C(_3580_),
    .Y(_3591_)
);

INVX1 _12023_ (
    .A(_3591_),
    .Y(_3612_)
);

NOR2X1 _12024_ (
    .A(_2562__bF$buf3),
    .B(_2508_),
    .Y(_3613_)
);

INVX1 _12025_ (
    .A(_3613_),
    .Y(_3624_)
);

NAND2X1 _12026_ (
    .A(breg_1_bF$buf0),
    .B(areg_6_bF$buf4),
    .Y(_3635_)
);

INVX8 _12027_ (
    .A(areg_6_bF$buf3),
    .Y(_3646_)
);

OAI21X1 _12028_ (
    .A(_2551__bF$buf1),
    .B(_3646__bF$buf3),
    .C(_2814_),
    .Y(_3657_)
);

OAI21X1 _12029_ (
    .A(_3569_),
    .B(_3635_),
    .C(_3657_),
    .Y(_3668_)
);

XNOR2X1 _12030_ (
    .A(_3668_),
    .B(_3624_),
    .Y(_3679_)
);

NAND2X1 _12031_ (
    .A(_3612_),
    .B(_3679_),
    .Y(_3690_)
);

XNOR2X1 _12032_ (
    .A(_3668_),
    .B(_3613_),
    .Y(_3701_)
);

NAND2X1 _12033_ (
    .A(_3591_),
    .B(_3701_),
    .Y(_3712_)
);

AOI21X1 _12034_ (
    .A(_3712_),
    .B(_3690_),
    .C(_3558_),
    .Y(_3723_)
);

NAND2X1 _12035_ (
    .A(_3612_),
    .B(_3701_),
    .Y(_3734_)
);

NAND2X1 _12036_ (
    .A(_3591_),
    .B(_3679_),
    .Y(_3745_)
);

AOI21X1 _12037_ (
    .A(_3734_),
    .B(_3745_),
    .C(_3547_),
    .Y(_3756_)
);

OAI21X1 _12038_ (
    .A(_3723_),
    .B(_3756_),
    .C(_3493_),
    .Y(_3776_)
);

NAND2X1 _12039_ (
    .A(_2781_),
    .B(_2913_),
    .Y(_3787_)
);

AOI21X1 _12040_ (
    .A(_2749_),
    .B(_3787_),
    .C(_2924_),
    .Y(_3788_)
);

NAND3X1 _12041_ (
    .A(_3547_),
    .B(_3734_),
    .C(_3745_),
    .Y(_3799_)
);

NOR2X1 _12042_ (
    .A(_3591_),
    .B(_3679_),
    .Y(_3810_)
);

NOR2X1 _12043_ (
    .A(_3612_),
    .B(_3701_),
    .Y(_3821_)
);

OAI21X1 _12044_ (
    .A(_3810_),
    .B(_3821_),
    .C(_3558_),
    .Y(_3832_)
);

NAND3X1 _12045_ (
    .A(_3788_),
    .B(_3799_),
    .C(_3832_),
    .Y(_3843_)
);

AOI21X1 _12046_ (
    .A(_3776_),
    .B(_3843_),
    .C(_3471_),
    .Y(_3854_)
);

NOR3X1 _12047_ (
    .A(_3723_),
    .B(_3756_),
    .C(_3788_),
    .Y(_3865_)
);

AOI21X1 _12048_ (
    .A(_3799_),
    .B(_3832_),
    .C(_3493_),
    .Y(_3876_)
);

OAI21X1 _12049_ (
    .A(_3865_),
    .B(_3876_),
    .C(_3471_),
    .Y(_3887_)
);

INVX1 _12050_ (
    .A(_3887_),
    .Y(_3898_)
);

OAI21X1 _12051_ (
    .A(_3898_),
    .B(_3854_),
    .C(_3383_),
    .Y(_3909_)
);

AOI21X1 _12052_ (
    .A(_2431_),
    .B(_2989_),
    .C(_3011_),
    .Y(_3920_)
);

INVX1 _12053_ (
    .A(_3854_),
    .Y(_3931_)
);

NAND3X1 _12054_ (
    .A(_3931_),
    .B(_3887_),
    .C(_3920_),
    .Y(_3942_)
);

AOI21X1 _12055_ (
    .A(_3909_),
    .B(_3942_),
    .C(_3372_),
    .Y(_3953_)
);

INVX1 _12056_ (
    .A(_3953_),
    .Y(_3964_)
);

NAND2X1 _12057_ (
    .A(_3942_),
    .B(_3909_),
    .Y(_3975_)
);

INVX1 _12058_ (
    .A(_3975_),
    .Y(_3986_)
);

NAND2X1 _12059_ (
    .A(_3372_),
    .B(_3986_),
    .Y(_3997_)
);

NAND3X1 _12060_ (
    .A(_3350_),
    .B(_3964_),
    .C(_3997_),
    .Y(_4008_)
);

INVX1 _12061_ (
    .A(_4008_),
    .Y(_4019_)
);

AOI21X1 _12062_ (
    .A(_3964_),
    .B(_3997_),
    .C(_3350_),
    .Y(_4030_)
);

NOR2X1 _12063_ (
    .A(_4030_),
    .B(_4019_),
    .Y(_0_[6])
);

NAND3X1 _12064_ (
    .A(_3931_),
    .B(_3887_),
    .C(_3383_),
    .Y(_4051_)
);

NAND3X1 _12065_ (
    .A(_3799_),
    .B(_3493_),
    .C(_3832_),
    .Y(_4061_)
);

OAI21X1 _12066_ (
    .A(_3876_),
    .B(_3471_),
    .C(_4061_),
    .Y(_4072_)
);

NAND2X1 _12067_ (
    .A(areg_1_bF$buf3),
    .B(breg_7_bF$buf5),
    .Y(_4083_)
);

NOR2X1 _12068_ (
    .A(_3394_),
    .B(_4083_),
    .Y(_4094_)
);

INVX2 _12069_ (
    .A(_4094_),
    .Y(_4105_)
);

INVX8 _12070_ (
    .A(breg_7_bF$buf4),
    .Y(_4116_)
);

NAND2X1 _12071_ (
    .A(areg_1_bF$buf2),
    .B(breg_6_bF$buf4),
    .Y(_4127_)
);

OAI21X1 _12072_ (
    .A(_2376__bF$buf3),
    .B(_4116__bF$buf4),
    .C(_4127_),
    .Y(_4138_)
);

AND2X2 _12073_ (
    .A(_4105_),
    .B(_4138_),
    .Y(_4149_)
);

NAND2X1 _12074_ (
    .A(areg_3_bF$buf0),
    .B(breg_4_bF$buf2),
    .Y(_4160_)
);

NAND3X1 _12075_ (
    .A(areg_1_bF$buf1),
    .B(breg_5_bF$buf0),
    .C(_3536_),
    .Y(_4171_)
);

OAI21X1 _12076_ (
    .A(_2727_),
    .B(_4160_),
    .C(_4171_),
    .Y(_4182_)
);

NOR2X1 _12077_ (
    .A(_4149_),
    .B(_4182_),
    .Y(_4193_)
);

NAND2X1 _12078_ (
    .A(_4149_),
    .B(_4182_),
    .Y(_4204_)
);

INVX2 _12079_ (
    .A(_4204_),
    .Y(_4215_)
);

NOR2X1 _12080_ (
    .A(_4193_),
    .B(_4215_),
    .Y(_4226_)
);

OAI21X1 _12081_ (
    .A(_3821_),
    .B(_3558_),
    .C(_3734_),
    .Y(_4237_)
);

INVX8 _12082_ (
    .A(breg_5_bF$buf3),
    .Y(_4258_)
);

NOR2X1 _12083_ (
    .A(_2519__bF$buf2),
    .B(_4258__bF$buf3),
    .Y(_4259_)
);

INVX2 _12084_ (
    .A(_4259_),
    .Y(_4270_)
);

NAND2X1 _12085_ (
    .A(areg_4_bF$buf1),
    .B(breg_3_bF$buf2),
    .Y(_4281_)
);

NOR2X1 _12086_ (
    .A(_4160_),
    .B(_4281_),
    .Y(_4292_)
);

AND2X2 _12087_ (
    .A(_4160_),
    .B(_4281_),
    .Y(_4303_)
);

NOR2X1 _12088_ (
    .A(_4292_),
    .B(_4303_),
    .Y(_4314_)
);

XNOR2X1 _12089_ (
    .A(_4314_),
    .B(_4270_),
    .Y(_4325_)
);

NAND2X1 _12090_ (
    .A(breg_0_bF$buf0),
    .B(areg_6_bF$buf2),
    .Y(_4336_)
);

NOR2X1 _12091_ (
    .A(_2814_),
    .B(_4336_),
    .Y(_4346_)
);

AOI21X1 _12092_ (
    .A(_3613_),
    .B(_3657_),
    .C(_4346_),
    .Y(_4357_)
);

INVX1 _12093_ (
    .A(_4357_),
    .Y(_4368_)
);

NOR2X1 _12094_ (
    .A(_2825__bF$buf3),
    .B(_2508_),
    .Y(_4379_)
);

NAND2X1 _12095_ (
    .A(breg_0_bF$buf6),
    .B(areg_7_bF$buf4),
    .Y(_4390_)
);

XOR2X1 _12096_ (
    .A(_3635_),
    .B(_4390_),
    .Y(_4401_)
);

NAND2X1 _12097_ (
    .A(_4379_),
    .B(_4401_),
    .Y(_4412_)
);

NAND2X1 _12098_ (
    .A(breg_1_bF$buf6),
    .B(areg_7_bF$buf3),
    .Y(_4423_)
);

INVX8 _12099_ (
    .A(areg_7_bF$buf2),
    .Y(_4434_)
);

OAI21X1 _12100_ (
    .A(_2551__bF$buf0),
    .B(_4434__bF$buf3),
    .C(_3635_),
    .Y(_4445_)
);

OAI21X1 _12101_ (
    .A(_4336_),
    .B(_4423_),
    .C(_4445_),
    .Y(_4466_)
);

OAI21X1 _12102_ (
    .A(_2825__bF$buf2),
    .B(_2508_),
    .C(_4466_),
    .Y(_4477_)
);

NAND3X1 _12103_ (
    .A(_4477_),
    .B(_4368_),
    .C(_4412_),
    .Y(_4478_)
);

INVX1 _12104_ (
    .A(_4379_),
    .Y(_4489_)
);

NOR2X1 _12105_ (
    .A(_4489_),
    .B(_4466_),
    .Y(_4500_)
);

NOR2X1 _12106_ (
    .A(_4379_),
    .B(_4401_),
    .Y(_4511_)
);

OAI21X1 _12107_ (
    .A(_4511_),
    .B(_4500_),
    .C(_4357_),
    .Y(_4522_)
);

NAND3X1 _12108_ (
    .A(_4325_),
    .B(_4478_),
    .C(_4522_),
    .Y(_4533_)
);

XNOR2X1 _12109_ (
    .A(_4314_),
    .B(_4259_),
    .Y(_4544_)
);

NOR3X1 _12110_ (
    .A(_4500_),
    .B(_4357_),
    .C(_4511_),
    .Y(_4555_)
);

AOI21X1 _12111_ (
    .A(_4477_),
    .B(_4412_),
    .C(_4368_),
    .Y(_4566_)
);

OAI21X1 _12112_ (
    .A(_4555_),
    .B(_4566_),
    .C(_4544_),
    .Y(_4577_)
);

NAND3X1 _12113_ (
    .A(_4533_),
    .B(_4577_),
    .C(_4237_),
    .Y(_4588_)
);

AOI21X1 _12114_ (
    .A(_3547_),
    .B(_3745_),
    .C(_3810_),
    .Y(_4599_)
);

NOR3X1 _12115_ (
    .A(_4544_),
    .B(_4566_),
    .C(_4555_),
    .Y(_4610_)
);

AOI21X1 _12116_ (
    .A(_4478_),
    .B(_4522_),
    .C(_4325_),
    .Y(_4621_)
);

OAI21X1 _12117_ (
    .A(_4610_),
    .B(_4621_),
    .C(_4599_),
    .Y(_4632_)
);

NAND3X1 _12118_ (
    .A(_4226_),
    .B(_4632_),
    .C(_4588_),
    .Y(_4642_)
);

OR2X2 _12119_ (
    .A(_4215_),
    .B(_4193_),
    .Y(_4653_)
);

NOR3X1 _12120_ (
    .A(_4610_),
    .B(_4621_),
    .C(_4599_),
    .Y(_4664_)
);

AOI21X1 _12121_ (
    .A(_4533_),
    .B(_4577_),
    .C(_4237_),
    .Y(_4675_)
);

OAI21X1 _12122_ (
    .A(_4664_),
    .B(_4675_),
    .C(_4653_),
    .Y(_4686_)
);

NAND3X1 _12123_ (
    .A(_4642_),
    .B(_4072_),
    .C(_4686_),
    .Y(_4697_)
);

NOR2X1 _12124_ (
    .A(_3438_),
    .B(_3460_),
    .Y(_4708_)
);

OAI21X1 _12125_ (
    .A(_3723_),
    .B(_3756_),
    .C(_3788_),
    .Y(_4719_)
);

AOI21X1 _12126_ (
    .A(_4708_),
    .B(_4719_),
    .C(_3865_),
    .Y(_4730_)
);

OAI21X1 _12127_ (
    .A(_4610_),
    .B(_4621_),
    .C(_4237_),
    .Y(_4741_)
);

NAND3X1 _12128_ (
    .A(_4533_),
    .B(_4577_),
    .C(_4599_),
    .Y(_4752_)
);

AOI21X1 _12129_ (
    .A(_4752_),
    .B(_4741_),
    .C(_4653_),
    .Y(_4763_)
);

AOI21X1 _12130_ (
    .A(_4632_),
    .B(_4588_),
    .C(_4226_),
    .Y(_4774_)
);

OAI21X1 _12131_ (
    .A(_4774_),
    .B(_4763_),
    .C(_4730_),
    .Y(_4785_)
);

NAND3X1 _12132_ (
    .A(_3460_),
    .B(_4785_),
    .C(_4697_),
    .Y(_4796_)
);

NOR3X1 _12133_ (
    .A(_4774_),
    .B(_4763_),
    .C(_4730_),
    .Y(_4807_)
);

AOI21X1 _12134_ (
    .A(_4642_),
    .B(_4686_),
    .C(_4072_),
    .Y(_4818_)
);

OAI21X1 _12135_ (
    .A(_4807_),
    .B(_4818_),
    .C(_3449_),
    .Y(_4829_)
);

NAND3X1 _12136_ (
    .A(_4051_),
    .B(_4796_),
    .C(_4829_),
    .Y(_4840_)
);

NOR3X1 _12137_ (
    .A(_3898_),
    .B(_3854_),
    .C(_3920_),
    .Y(_4851_)
);

NAND3X1 _12138_ (
    .A(_3449_),
    .B(_4785_),
    .C(_4697_),
    .Y(_4862_)
);

OAI21X1 _12139_ (
    .A(_4807_),
    .B(_4818_),
    .C(_3460_),
    .Y(_4873_)
);

NAND3X1 _12140_ (
    .A(_4862_),
    .B(_4851_),
    .C(_4873_),
    .Y(_4884_)
);

NAND2X1 _12141_ (
    .A(_4840_),
    .B(_4884_),
    .Y(_4895_)
);

OAI21X1 _12142_ (
    .A(_3372_),
    .B(_3986_),
    .C(_4895_),
    .Y(_4906_)
);

NAND3X1 _12143_ (
    .A(_3953_),
    .B(_4840_),
    .C(_4884_),
    .Y(_4917_)
);

AOI21X1 _12144_ (
    .A(_4917_),
    .B(_4906_),
    .C(_4008_),
    .Y(_4928_)
);

NAND2X1 _12145_ (
    .A(_4917_),
    .B(_4906_),
    .Y(_4939_)
);

NOR2X1 _12146_ (
    .A(_4939_),
    .B(_4019_),
    .Y(_4950_)
);

NOR2X1 _12147_ (
    .A(_4928_),
    .B(_4950_),
    .Y(_0_[7])
);

AOI21X1 _12148_ (
    .A(_4862_),
    .B(_4873_),
    .C(_4051_),
    .Y(_4970_)
);

OAI21X1 _12149_ (
    .A(_4818_),
    .B(_3449_),
    .C(_4697_),
    .Y(_4981_)
);

OAI21X1 _12150_ (
    .A(_4653_),
    .B(_4675_),
    .C(_4588_),
    .Y(_4992_)
);

OAI21X1 _12151_ (
    .A(_4566_),
    .B(_4544_),
    .C(_4478_),
    .Y(_5003_)
);

NOR2X1 _12152_ (
    .A(_2792_),
    .B(_4258__bF$buf2),
    .Y(_5014_)
);

INVX2 _12153_ (
    .A(_5014_),
    .Y(_5025_)
);

NAND2X1 _12154_ (
    .A(areg_4_bF$buf0),
    .B(breg_4_bF$buf1),
    .Y(_5036_)
);

NAND2X1 _12155_ (
    .A(areg_5_bF$buf1),
    .B(breg_3_bF$buf1),
    .Y(_5047_)
);

NOR2X1 _12156_ (
    .A(_5036_),
    .B(_5047_),
    .Y(_5058_)
);

AND2X2 _12157_ (
    .A(_5036_),
    .B(_5047_),
    .Y(_5069_)
);

NOR2X1 _12158_ (
    .A(_5058_),
    .B(_5069_),
    .Y(_5080_)
);

XNOR2X1 _12159_ (
    .A(_5080_),
    .B(_5025_),
    .Y(_5091_)
);

NOR2X1 _12160_ (
    .A(_3635_),
    .B(_4390_),
    .Y(_5102_)
);

AOI21X1 _12161_ (
    .A(_4379_),
    .B(_4445_),
    .C(_5102_),
    .Y(_5113_)
);

INVX2 _12162_ (
    .A(_5113_),
    .Y(_5124_)
);

NOR2X1 _12163_ (
    .A(_2508_),
    .B(_3646__bF$buf2),
    .Y(_5135_)
);

NAND2X1 _12164_ (
    .A(breg_0_bF$buf5),
    .B(areg_8_bF$buf4),
    .Y(_5146_)
);

XOR2X1 _12165_ (
    .A(_4423_),
    .B(_5146_),
    .Y(_5157_)
);

NAND2X1 _12166_ (
    .A(_5135_),
    .B(_5157_),
    .Y(_5168_)
);

NAND2X1 _12167_ (
    .A(breg_1_bF$buf5),
    .B(areg_8_bF$buf3),
    .Y(_5179_)
);

INVX8 _12168_ (
    .A(areg_8_bF$buf2),
    .Y(_5190_)
);

OAI21X1 _12169_ (
    .A(_2551__bF$buf3),
    .B(_5190__bF$buf3),
    .C(_4423_),
    .Y(_5201_)
);

OAI21X1 _12170_ (
    .A(_4390_),
    .B(_5179_),
    .C(_5201_),
    .Y(_5212_)
);

OAI21X1 _12171_ (
    .A(_2508_),
    .B(_3646__bF$buf1),
    .C(_5212_),
    .Y(_5233_)
);

NAND3X1 _12172_ (
    .A(_5233_),
    .B(_5124_),
    .C(_5168_),
    .Y(_5244_)
);

INVX1 _12173_ (
    .A(_5135_),
    .Y(_5245_)
);

NOR2X1 _12174_ (
    .A(_5245_),
    .B(_5212_),
    .Y(_5256_)
);

NOR2X1 _12175_ (
    .A(_5135_),
    .B(_5157_),
    .Y(_5267_)
);

OAI21X1 _12176_ (
    .A(_5267_),
    .B(_5256_),
    .C(_5113_),
    .Y(_5278_)
);

NAND3X1 _12177_ (
    .A(_5091_),
    .B(_5244_),
    .C(_5278_),
    .Y(_5289_)
);

XNOR2X1 _12178_ (
    .A(_5080_),
    .B(_5014_),
    .Y(_5299_)
);

NOR3X1 _12179_ (
    .A(_5256_),
    .B(_5113_),
    .C(_5267_),
    .Y(_5310_)
);

AOI21X1 _12180_ (
    .A(_5233_),
    .B(_5168_),
    .C(_5124_),
    .Y(_5321_)
);

OAI21X1 _12181_ (
    .A(_5310_),
    .B(_5321_),
    .C(_5299_),
    .Y(_5332_)
);

AOI21X1 _12182_ (
    .A(_5289_),
    .B(_5332_),
    .C(_5003_),
    .Y(_5343_)
);

AOI21X1 _12183_ (
    .A(_4325_),
    .B(_4522_),
    .C(_4555_),
    .Y(_5354_)
);

OAI21X1 _12184_ (
    .A(_5267_),
    .B(_5256_),
    .C(_5124_),
    .Y(_5365_)
);

NAND3X1 _12185_ (
    .A(_5113_),
    .B(_5233_),
    .C(_5168_),
    .Y(_5376_)
);

AOI21X1 _12186_ (
    .A(_5376_),
    .B(_5365_),
    .C(_5299_),
    .Y(_5387_)
);

AOI21X1 _12187_ (
    .A(_5244_),
    .B(_5278_),
    .C(_5091_),
    .Y(_5398_)
);

NOR3X1 _12188_ (
    .A(_5387_),
    .B(_5398_),
    .C(_5354_),
    .Y(_5409_)
);

INVX8 _12189_ (
    .A(breg[8]),
    .Y(_5420_)
);

NOR2X1 _12190_ (
    .A(_2376__bF$buf2),
    .B(_5420__bF$buf3),
    .Y(_5431_)
);

NAND2X1 _12191_ (
    .A(areg_2_bF$buf4),
    .B(breg_7_bF$buf3),
    .Y(_5442_)
);

INVX8 _12192_ (
    .A(breg_6_bF$buf3),
    .Y(_5453_)
);

OAI21X1 _12193_ (
    .A(_2519__bF$buf1),
    .B(_5453__bF$buf5),
    .C(_4083_),
    .Y(_5464_)
);

OAI21X1 _12194_ (
    .A(_4127_),
    .B(_5442_),
    .C(_5464_),
    .Y(_5475_)
);

XNOR2X1 _12195_ (
    .A(_5475_),
    .B(_5431_),
    .Y(_5486_)
);

OAI22X1 _12196_ (
    .A(_3525_),
    .B(_5036_),
    .C(_4270_),
    .D(_4303_),
    .Y(_5497_)
);

NAND2X1 _12197_ (
    .A(_5497_),
    .B(_5486_),
    .Y(_5508_)
);

OAI21X1 _12198_ (
    .A(_2376__bF$buf1),
    .B(_5420__bF$buf2),
    .C(_5475_),
    .Y(_5519_)
);

NAND2X1 _12199_ (
    .A(areg_2_bF$buf3),
    .B(breg_6_bF$buf2),
    .Y(_5530_)
);

OR2X2 _12200_ (
    .A(_4083_),
    .B(_5530_),
    .Y(_5541_)
);

NAND3X1 _12201_ (
    .A(_5431_),
    .B(_5464_),
    .C(_5541_),
    .Y(_5552_)
);

NAND2X1 _12202_ (
    .A(_5552_),
    .B(_5519_),
    .Y(_5563_)
);

INVX1 _12203_ (
    .A(_5497_),
    .Y(_5574_)
);

NAND2X1 _12204_ (
    .A(_5574_),
    .B(_5563_),
    .Y(_5585_)
);

NAND3X1 _12205_ (
    .A(_4105_),
    .B(_5508_),
    .C(_5585_),
    .Y(_5596_)
);

NAND2X1 _12206_ (
    .A(_5574_),
    .B(_5486_),
    .Y(_5607_)
);

NAND2X1 _12207_ (
    .A(_5497_),
    .B(_5563_),
    .Y(_5618_)
);

NAND3X1 _12208_ (
    .A(_4094_),
    .B(_5607_),
    .C(_5618_),
    .Y(_5629_)
);

AND2X2 _12209_ (
    .A(_5596_),
    .B(_5629_),
    .Y(_5640_)
);

OAI21X1 _12210_ (
    .A(_5409_),
    .B(_5343_),
    .C(_5640_),
    .Y(_5651_)
);

OAI21X1 _12211_ (
    .A(_5387_),
    .B(_5398_),
    .C(_5354_),
    .Y(_5661_)
);

NAND3X1 _12212_ (
    .A(_5003_),
    .B(_5289_),
    .C(_5332_),
    .Y(_5672_)
);

NAND2X1 _12213_ (
    .A(_5596_),
    .B(_5629_),
    .Y(_5683_)
);

NAND3X1 _12214_ (
    .A(_5683_),
    .B(_5661_),
    .C(_5672_),
    .Y(_5694_)
);

AOI21X1 _12215_ (
    .A(_5694_),
    .B(_5651_),
    .C(_4992_),
    .Y(_5705_)
);

AOI21X1 _12216_ (
    .A(_4226_),
    .B(_4632_),
    .C(_4664_),
    .Y(_5716_)
);

AOI21X1 _12217_ (
    .A(_5661_),
    .B(_5672_),
    .C(_5683_),
    .Y(_5727_)
);

NOR3X1 _12218_ (
    .A(_5409_),
    .B(_5343_),
    .C(_5640_),
    .Y(_5738_)
);

NOR3X1 _12219_ (
    .A(_5716_),
    .B(_5727_),
    .C(_5738_),
    .Y(_5749_)
);

OAI21X1 _12220_ (
    .A(_5749_),
    .B(_5705_),
    .C(_4204_),
    .Y(_5760_)
);

OAI21X1 _12221_ (
    .A(_5738_),
    .B(_5727_),
    .C(_5716_),
    .Y(_5771_)
);

NAND3X1 _12222_ (
    .A(_5694_),
    .B(_5651_),
    .C(_4992_),
    .Y(_5792_)
);

NAND3X1 _12223_ (
    .A(_4215_),
    .B(_5792_),
    .C(_5771_),
    .Y(_5793_)
);

NAND3X1 _12224_ (
    .A(_4981_),
    .B(_5793_),
    .C(_5760_),
    .Y(_5804_)
);

AOI21X1 _12225_ (
    .A(_3460_),
    .B(_4785_),
    .C(_4807_),
    .Y(_5815_)
);

AOI21X1 _12226_ (
    .A(_5792_),
    .B(_5771_),
    .C(_4215_),
    .Y(_5826_)
);

NOR3X1 _12227_ (
    .A(_4204_),
    .B(_5705_),
    .C(_5749_),
    .Y(_5837_)
);

OAI21X1 _12228_ (
    .A(_5837_),
    .B(_5826_),
    .C(_5815_),
    .Y(_5848_)
);

NAND3X1 _12229_ (
    .A(_4970_),
    .B(_5804_),
    .C(_5848_),
    .Y(_5859_)
);

NAND3X1 _12230_ (
    .A(_4796_),
    .B(_4851_),
    .C(_4829_),
    .Y(_5870_)
);

NAND3X1 _12231_ (
    .A(_4051_),
    .B(_4862_),
    .C(_4873_),
    .Y(_5881_)
);

NAND3X1 _12232_ (
    .A(_3953_),
    .B(_5881_),
    .C(_5870_),
    .Y(_5892_)
);

NAND2X1 _12233_ (
    .A(_5804_),
    .B(_5848_),
    .Y(_5903_)
);

NOR2X1 _12234_ (
    .A(_5892_),
    .B(_5903_),
    .Y(_5914_)
);

AOI22X1 _12235_ (
    .A(_5804_),
    .B(_5848_),
    .C(_4895_),
    .D(_3953_),
    .Y(_5925_)
);

OAI21X1 _12236_ (
    .A(_5914_),
    .B(_5925_),
    .C(_5870_),
    .Y(_5936_)
);

NAND3X1 _12237_ (
    .A(_4928_),
    .B(_5859_),
    .C(_5936_),
    .Y(_5947_)
);

INVX1 _12238_ (
    .A(_5947_),
    .Y(_5958_)
);

AOI21X1 _12239_ (
    .A(_5859_),
    .B(_5936_),
    .C(_4928_),
    .Y(_5969_)
);

NOR2X1 _12240_ (
    .A(_5969_),
    .B(_5958_),
    .Y(_0_[8])
);

OAI21X1 _12241_ (
    .A(_5837_),
    .B(_5826_),
    .C(_4981_),
    .Y(_5990_)
);

NAND3X1 _12242_ (
    .A(_5815_),
    .B(_5793_),
    .C(_5760_),
    .Y(_6001_)
);

AOI21X1 _12243_ (
    .A(_6001_),
    .B(_5990_),
    .C(_5870_),
    .Y(_6012_)
);

NOR3X1 _12244_ (
    .A(_5815_),
    .B(_5826_),
    .C(_5837_),
    .Y(_6023_)
);

OAI21X1 _12245_ (
    .A(_5705_),
    .B(_4204_),
    .C(_5792_),
    .Y(_6034_)
);

INVX8 _12246_ (
    .A(breg_9_bF$buf5),
    .Y(_6044_)
);

NOR2X1 _12247_ (
    .A(_2376__bF$buf0),
    .B(_6044__bF$buf5),
    .Y(_6055_)
);

INVX1 _12248_ (
    .A(_5585_),
    .Y(_6076_)
);

OAI21X1 _12249_ (
    .A(_6076_),
    .B(_4105_),
    .C(_5508_),
    .Y(_6087_)
);

XNOR2X1 _12250_ (
    .A(_6087_),
    .B(_6055_),
    .Y(_6088_)
);

INVX2 _12251_ (
    .A(_6088_),
    .Y(_6099_)
);

OAI21X1 _12252_ (
    .A(_5640_),
    .B(_5343_),
    .C(_5672_),
    .Y(_6110_)
);

OAI21X1 _12253_ (
    .A(_4127_),
    .B(_5442_),
    .C(_5552_),
    .Y(_6121_)
);

NOR2X1 _12254_ (
    .A(_2661_),
    .B(_5420__bF$buf1),
    .Y(_6132_)
);

NAND2X1 _12255_ (
    .A(areg_3_bF$buf4),
    .B(breg_7_bF$buf2),
    .Y(_6143_)
);

OAI21X1 _12256_ (
    .A(_2792_),
    .B(_5453__bF$buf4),
    .C(_5442_),
    .Y(_6154_)
);

OAI21X1 _12257_ (
    .A(_5530_),
    .B(_6143_),
    .C(_6154_),
    .Y(_6165_)
);

XNOR2X1 _12258_ (
    .A(_6165_),
    .B(_6132_),
    .Y(_6176_)
);

NAND2X1 _12259_ (
    .A(areg_5_bF$buf0),
    .B(breg_4_bF$buf0),
    .Y(_6187_)
);

OAI22X1 _12260_ (
    .A(_4281_),
    .B(_6187_),
    .C(_5025_),
    .D(_5069_),
    .Y(_6198_)
);

NAND2X1 _12261_ (
    .A(_6198_),
    .B(_6176_),
    .Y(_6209_)
);

NAND2X1 _12262_ (
    .A(areg_3_bF$buf3),
    .B(breg_6_bF$buf1),
    .Y(_6220_)
);

XOR2X1 _12263_ (
    .A(_5442_),
    .B(_6220_),
    .Y(_6231_)
);

NOR2X1 _12264_ (
    .A(_6132_),
    .B(_6231_),
    .Y(_6242_)
);

AND2X2 _12265_ (
    .A(_6231_),
    .B(_6132_),
    .Y(_6253_)
);

INVX1 _12266_ (
    .A(_6198_),
    .Y(_6264_)
);

OAI21X1 _12267_ (
    .A(_6253_),
    .B(_6242_),
    .C(_6264_),
    .Y(_6275_)
);

NAND3X1 _12268_ (
    .A(_6121_),
    .B(_6275_),
    .C(_6209_),
    .Y(_6286_)
);

INVX1 _12269_ (
    .A(_6121_),
    .Y(_6297_)
);

NAND2X1 _12270_ (
    .A(_6264_),
    .B(_6176_),
    .Y(_6308_)
);

OAI21X1 _12271_ (
    .A(_6253_),
    .B(_6242_),
    .C(_6198_),
    .Y(_6319_)
);

NAND3X1 _12272_ (
    .A(_6297_),
    .B(_6319_),
    .C(_6308_),
    .Y(_6330_)
);

AND2X2 _12273_ (
    .A(_6286_),
    .B(_6330_),
    .Y(_6341_)
);

OAI21X1 _12274_ (
    .A(_5321_),
    .B(_5299_),
    .C(_5244_),
    .Y(_6352_)
);

NOR2X1 _12275_ (
    .A(_2562__bF$buf2),
    .B(_4258__bF$buf1),
    .Y(_6363_)
);

INVX2 _12276_ (
    .A(_6363_),
    .Y(_6374_)
);

NAND2X1 _12277_ (
    .A(breg_3_bF$buf0),
    .B(areg_6_bF$buf1),
    .Y(_6385_)
);

NOR2X1 _12278_ (
    .A(_6187_),
    .B(_6385_),
    .Y(_6396_)
);

AND2X2 _12279_ (
    .A(_6187_),
    .B(_6385_),
    .Y(_6407_)
);

NOR2X1 _12280_ (
    .A(_6396_),
    .B(_6407_),
    .Y(_6417_)
);

XNOR2X1 _12281_ (
    .A(_6417_),
    .B(_6374_),
    .Y(_6428_)
);

NOR2X1 _12282_ (
    .A(_4423_),
    .B(_5146_),
    .Y(_6439_)
);

AOI21X1 _12283_ (
    .A(_5135_),
    .B(_5201_),
    .C(_6439_),
    .Y(_6450_)
);

INVX2 _12284_ (
    .A(_6450_),
    .Y(_6461_)
);

NOR2X1 _12285_ (
    .A(_2508_),
    .B(_4434__bF$buf2),
    .Y(_6472_)
);

NAND2X1 _12286_ (
    .A(breg_0_bF$buf4),
    .B(areg_9_bF$buf4),
    .Y(_6483_)
);

XOR2X1 _12287_ (
    .A(_5179_),
    .B(_6483_),
    .Y(_6494_)
);

NAND2X1 _12288_ (
    .A(_6472_),
    .B(_6494_),
    .Y(_6505_)
);

INVX1 _12289_ (
    .A(_6472_),
    .Y(_6516_)
);

NOR2X1 _12290_ (
    .A(_5179_),
    .B(_6483_),
    .Y(_6527_)
);

AND2X2 _12291_ (
    .A(_5179_),
    .B(_6483_),
    .Y(_6538_)
);

OAI21X1 _12292_ (
    .A(_6538_),
    .B(_6527_),
    .C(_6516_),
    .Y(_6549_)
);

NAND3X1 _12293_ (
    .A(_6549_),
    .B(_6461_),
    .C(_6505_),
    .Y(_6560_)
);

NAND2X1 _12294_ (
    .A(breg_1_bF$buf4),
    .B(areg_9_bF$buf3),
    .Y(_6571_)
);

INVX8 _12295_ (
    .A(areg_9_bF$buf2),
    .Y(_6582_)
);

OAI21X1 _12296_ (
    .A(_2551__bF$buf2),
    .B(_6582__bF$buf3),
    .C(_5179_),
    .Y(_6593_)
);

OAI21X1 _12297_ (
    .A(_5146_),
    .B(_6571_),
    .C(_6593_),
    .Y(_6604_)
);

NOR2X1 _12298_ (
    .A(_6516_),
    .B(_6604_),
    .Y(_6615_)
);

NOR2X1 _12299_ (
    .A(_6472_),
    .B(_6494_),
    .Y(_6626_)
);

OAI21X1 _12300_ (
    .A(_6626_),
    .B(_6615_),
    .C(_6450_),
    .Y(_6637_)
);

NAND3X1 _12301_ (
    .A(_6428_),
    .B(_6560_),
    .C(_6637_),
    .Y(_6658_)
);

XNOR2X1 _12302_ (
    .A(_6417_),
    .B(_6363_),
    .Y(_6659_)
);

NOR3X1 _12303_ (
    .A(_6615_),
    .B(_6450_),
    .C(_6626_),
    .Y(_6670_)
);

AOI21X1 _12304_ (
    .A(_6549_),
    .B(_6505_),
    .C(_6461_),
    .Y(_6681_)
);

OAI21X1 _12305_ (
    .A(_6670_),
    .B(_6681_),
    .C(_6659_),
    .Y(_6692_)
);

NAND3X1 _12306_ (
    .A(_6352_),
    .B(_6658_),
    .C(_6692_),
    .Y(_6703_)
);

AOI21X1 _12307_ (
    .A(_5091_),
    .B(_5278_),
    .C(_5310_),
    .Y(_6714_)
);

OAI21X1 _12308_ (
    .A(_6626_),
    .B(_6615_),
    .C(_6461_),
    .Y(_6725_)
);

NAND3X1 _12309_ (
    .A(_6450_),
    .B(_6549_),
    .C(_6505_),
    .Y(_6736_)
);

AOI21X1 _12310_ (
    .A(_6736_),
    .B(_6725_),
    .C(_6659_),
    .Y(_6747_)
);

AOI21X1 _12311_ (
    .A(_6560_),
    .B(_6637_),
    .C(_6428_),
    .Y(_6758_)
);

OAI21X1 _12312_ (
    .A(_6747_),
    .B(_6758_),
    .C(_6714_),
    .Y(_6769_)
);

NAND3X1 _12313_ (
    .A(_6703_),
    .B(_6769_),
    .C(_6341_),
    .Y(_6780_)
);

NAND2X1 _12314_ (
    .A(_6286_),
    .B(_6330_),
    .Y(_6791_)
);

NOR3X1 _12315_ (
    .A(_6747_),
    .B(_6758_),
    .C(_6714_),
    .Y(_6802_)
);

AOI21X1 _12316_ (
    .A(_6658_),
    .B(_6692_),
    .C(_6352_),
    .Y(_6812_)
);

OAI21X1 _12317_ (
    .A(_6802_),
    .B(_6812_),
    .C(_6791_),
    .Y(_6823_)
);

NAND3X1 _12318_ (
    .A(_6780_),
    .B(_6823_),
    .C(_6110_),
    .Y(_6834_)
);

AOI21X1 _12319_ (
    .A(_5661_),
    .B(_5683_),
    .C(_5409_),
    .Y(_6845_)
);

OAI21X1 _12320_ (
    .A(_6747_),
    .B(_6758_),
    .C(_6352_),
    .Y(_6856_)
);

NAND3X1 _12321_ (
    .A(_6714_),
    .B(_6658_),
    .C(_6692_),
    .Y(_6867_)
);

AOI21X1 _12322_ (
    .A(_6856_),
    .B(_6867_),
    .C(_6791_),
    .Y(_6878_)
);

AOI21X1 _12323_ (
    .A(_6703_),
    .B(_6769_),
    .C(_6341_),
    .Y(_6889_)
);

OAI21X1 _12324_ (
    .A(_6889_),
    .B(_6878_),
    .C(_6845_),
    .Y(_6900_)
);

NAND3X1 _12325_ (
    .A(_6099_),
    .B(_6900_),
    .C(_6834_),
    .Y(_6911_)
);

NOR3X1 _12326_ (
    .A(_6889_),
    .B(_6878_),
    .C(_6845_),
    .Y(_6922_)
);

AOI21X1 _12327_ (
    .A(_6780_),
    .B(_6823_),
    .C(_6110_),
    .Y(_6933_)
);

OAI21X1 _12328_ (
    .A(_6922_),
    .B(_6933_),
    .C(_6088_),
    .Y(_6944_)
);

NAND3X1 _12329_ (
    .A(_6911_),
    .B(_6034_),
    .C(_6944_),
    .Y(_6955_)
);

AOI21X1 _12330_ (
    .A(_4215_),
    .B(_5771_),
    .C(_5749_),
    .Y(_6966_)
);

NOR3X1 _12331_ (
    .A(_6933_),
    .B(_6088_),
    .C(_6922_),
    .Y(_6977_)
);

AOI21X1 _12332_ (
    .A(_6900_),
    .B(_6834_),
    .C(_6099_),
    .Y(_6988_)
);

OAI21X1 _12333_ (
    .A(_6977_),
    .B(_6988_),
    .C(_6966_),
    .Y(_6999_)
);

NAND3X1 _12334_ (
    .A(_6955_),
    .B(_6999_),
    .C(_6023_),
    .Y(_7020_)
);

OAI21X1 _12335_ (
    .A(_6977_),
    .B(_6988_),
    .C(_6034_),
    .Y(_7031_)
);

NAND3X1 _12336_ (
    .A(_6911_),
    .B(_6944_),
    .C(_6966_),
    .Y(_7032_)
);

NAND3X1 _12337_ (
    .A(_7032_),
    .B(_7031_),
    .C(_5804_),
    .Y(_7043_)
);

NAND3X1 _12338_ (
    .A(_7043_),
    .B(_6012_),
    .C(_7020_),
    .Y(_7054_)
);

AOI21X1 _12339_ (
    .A(_7032_),
    .B(_7031_),
    .C(_5804_),
    .Y(_7065_)
);

NOR2X1 _12340_ (
    .A(_5826_),
    .B(_5837_),
    .Y(_7076_)
);

AOI22X1 _12341_ (
    .A(_6955_),
    .B(_6999_),
    .C(_7076_),
    .D(_4981_),
    .Y(_7087_)
);

OAI21X1 _12342_ (
    .A(_7087_),
    .B(_7065_),
    .C(_5859_),
    .Y(_7098_)
);

NAND3X1 _12343_ (
    .A(_5914_),
    .B(_7098_),
    .C(_7054_),
    .Y(_7109_)
);

OR2X2 _12344_ (
    .A(_5903_),
    .B(_5892_),
    .Y(_7120_)
);

NAND3X1 _12345_ (
    .A(_7043_),
    .B(_5859_),
    .C(_7020_),
    .Y(_7131_)
);

OAI21X1 _12346_ (
    .A(_7087_),
    .B(_7065_),
    .C(_6012_),
    .Y(_7142_)
);

NAND3X1 _12347_ (
    .A(_7120_),
    .B(_7142_),
    .C(_7131_),
    .Y(_7153_)
);

NAND2X1 _12348_ (
    .A(_7109_),
    .B(_7153_),
    .Y(_7164_)
);

XOR2X1 _12349_ (
    .A(_7164_),
    .B(_5947_),
    .Y(_0_[9])
);

NAND2X1 _12350_ (
    .A(_6055_),
    .B(_6087_),
    .Y(_7185_)
);

OAI21X1 _12351_ (
    .A(_6933_),
    .B(_6088_),
    .C(_6834_),
    .Y(_7196_)
);

NAND3X1 _12352_ (
    .A(areg_1_bF$buf0),
    .B(breg_10_bF$buf5),
    .C(_6055_),
    .Y(_7207_)
);

INVX8 _12353_ (
    .A(breg_10_bF$buf4),
    .Y(_7217_)
);

NAND2X1 _12354_ (
    .A(areg_1_bF$buf4),
    .B(breg_9_bF$buf4),
    .Y(_7228_)
);

OAI21X1 _12355_ (
    .A(_2376__bF$buf3),
    .B(_7217__bF$buf4),
    .C(_7228_),
    .Y(_7239_)
);

AND2X2 _12356_ (
    .A(_7207_),
    .B(_7239_),
    .Y(_7250_)
);

NAND2X1 _12357_ (
    .A(_6209_),
    .B(_6286_),
    .Y(_7261_)
);

XNOR2X1 _12358_ (
    .A(_7261_),
    .B(_7250_),
    .Y(_7272_)
);

INVX2 _12359_ (
    .A(_7272_),
    .Y(_7283_)
);

OAI21X1 _12360_ (
    .A(_6812_),
    .B(_6791_),
    .C(_6703_),
    .Y(_7294_)
);

NOR2X1 _12361_ (
    .A(_5442_),
    .B(_6220_),
    .Y(_7305_)
);

NOR2X1 _12362_ (
    .A(_7305_),
    .B(_6253_),
    .Y(_7316_)
);

NOR2X1 _12363_ (
    .A(_2519__bF$buf0),
    .B(_5420__bF$buf0),
    .Y(_7327_)
);

NAND2X1 _12364_ (
    .A(areg_4_bF$buf4),
    .B(breg_7_bF$buf1),
    .Y(_7338_)
);

OAI21X1 _12365_ (
    .A(_2562__bF$buf1),
    .B(_5453__bF$buf3),
    .C(_6143_),
    .Y(_7349_)
);

OAI21X1 _12366_ (
    .A(_6220_),
    .B(_7338_),
    .C(_7349_),
    .Y(_7360_)
);

XNOR2X1 _12367_ (
    .A(_7360_),
    .B(_7327_),
    .Y(_7371_)
);

NAND2X1 _12368_ (
    .A(breg_4_bF$buf5),
    .B(areg_6_bF$buf0),
    .Y(_7382_)
);

OAI22X1 _12369_ (
    .A(_5047_),
    .B(_7382_),
    .C(_6374_),
    .D(_6407_),
    .Y(_7393_)
);

NAND2X1 _12370_ (
    .A(_7393_),
    .B(_7371_),
    .Y(_7404_)
);

OAI21X1 _12371_ (
    .A(_2519__bF$buf3),
    .B(_5420__bF$buf3),
    .C(_7360_),
    .Y(_7415_)
);

NAND2X1 _12372_ (
    .A(areg_4_bF$buf3),
    .B(breg_6_bF$buf0),
    .Y(_7426_)
);

OR2X2 _12373_ (
    .A(_6143_),
    .B(_7426_),
    .Y(_7437_)
);

NAND3X1 _12374_ (
    .A(_7327_),
    .B(_7349_),
    .C(_7437_),
    .Y(_7448_)
);

NAND2X1 _12375_ (
    .A(_7448_),
    .B(_7415_),
    .Y(_7459_)
);

INVX2 _12376_ (
    .A(_7393_),
    .Y(_7470_)
);

NAND2X1 _12377_ (
    .A(_7470_),
    .B(_7459_),
    .Y(_7481_)
);

NAND3X1 _12378_ (
    .A(_7316_),
    .B(_7404_),
    .C(_7481_),
    .Y(_7492_)
);

OR2X2 _12379_ (
    .A(_6253_),
    .B(_7305_),
    .Y(_7503_)
);

NAND2X1 _12380_ (
    .A(_7470_),
    .B(_7371_),
    .Y(_7514_)
);

NAND2X1 _12381_ (
    .A(_7393_),
    .B(_7459_),
    .Y(_7525_)
);

NAND3X1 _12382_ (
    .A(_7503_),
    .B(_7514_),
    .C(_7525_),
    .Y(_7536_)
);

NAND2X1 _12383_ (
    .A(_7492_),
    .B(_7536_),
    .Y(_7547_)
);

OAI21X1 _12384_ (
    .A(_6681_),
    .B(_6659_),
    .C(_6560_),
    .Y(_7558_)
);

NOR2X1 _12385_ (
    .A(_2825__bF$buf1),
    .B(_4258__bF$buf0),
    .Y(_7569_)
);

INVX2 _12386_ (
    .A(_7569_),
    .Y(_7580_)
);

NAND2X1 _12387_ (
    .A(breg_4_bF$buf4),
    .B(areg_7_bF$buf1),
    .Y(_7591_)
);

NOR2X1 _12388_ (
    .A(_6385_),
    .B(_7591_),
    .Y(_7602_)
);

AOI22X1 _12389_ (
    .A(breg_3_bF$buf5),
    .B(areg_7_bF$buf0),
    .C(breg_4_bF$buf3),
    .D(areg_6_bF$buf4),
    .Y(_7623_)
);

NOR2X1 _12390_ (
    .A(_7623_),
    .B(_7602_),
    .Y(_7624_)
);

XNOR2X1 _12391_ (
    .A(_7624_),
    .B(_7580_),
    .Y(_7635_)
);

AOI21X1 _12392_ (
    .A(_6472_),
    .B(_6593_),
    .C(_6527_),
    .Y(_7645_)
);

INVX1 _12393_ (
    .A(_7645_),
    .Y(_7656_)
);

NAND2X1 _12394_ (
    .A(breg_2_bF$buf2),
    .B(areg_8_bF$buf1),
    .Y(_7667_)
);

INVX2 _12395_ (
    .A(_7667_),
    .Y(_7678_)
);

NAND2X1 _12396_ (
    .A(breg_0_bF$buf3),
    .B(areg_10_bF$buf4),
    .Y(_7689_)
);

OR2X2 _12397_ (
    .A(_6571_),
    .B(_7689_),
    .Y(_7700_)
);

INVX8 _12398_ (
    .A(areg_10_bF$buf3),
    .Y(_7711_)
);

OAI21X1 _12399_ (
    .A(_2551__bF$buf1),
    .B(_7711__bF$buf3),
    .C(_6571_),
    .Y(_7722_)
);

NAND3X1 _12400_ (
    .A(_7678_),
    .B(_7722_),
    .C(_7700_),
    .Y(_7733_)
);

NOR2X1 _12401_ (
    .A(_6571_),
    .B(_7689_),
    .Y(_7744_)
);

AND2X2 _12402_ (
    .A(_6571_),
    .B(_7689_),
    .Y(_7755_)
);

OAI21X1 _12403_ (
    .A(_7755_),
    .B(_7744_),
    .C(_7667_),
    .Y(_7766_)
);

NAND3X1 _12404_ (
    .A(_7766_),
    .B(_7733_),
    .C(_7656_),
    .Y(_7777_)
);

NOR3X1 _12405_ (
    .A(_7667_),
    .B(_7744_),
    .C(_7755_),
    .Y(_7788_)
);

AOI21X1 _12406_ (
    .A(_7722_),
    .B(_7700_),
    .C(_7678_),
    .Y(_7799_)
);

OAI21X1 _12407_ (
    .A(_7788_),
    .B(_7799_),
    .C(_7645_),
    .Y(_7810_)
);

NAND3X1 _12408_ (
    .A(_7635_),
    .B(_7810_),
    .C(_7777_),
    .Y(_7821_)
);

XNOR2X1 _12409_ (
    .A(_7624_),
    .B(_7569_),
    .Y(_7832_)
);

NOR3X1 _12410_ (
    .A(_7799_),
    .B(_7645_),
    .C(_7788_),
    .Y(_7843_)
);

AOI21X1 _12411_ (
    .A(_7766_),
    .B(_7733_),
    .C(_7656_),
    .Y(_7854_)
);

OAI21X1 _12412_ (
    .A(_7854_),
    .B(_7843_),
    .C(_7832_),
    .Y(_7865_)
);

NAND3X1 _12413_ (
    .A(_7821_),
    .B(_7865_),
    .C(_7558_),
    .Y(_7876_)
);

AOI21X1 _12414_ (
    .A(_6428_),
    .B(_6637_),
    .C(_6670_),
    .Y(_7887_)
);

NOR3X1 _12415_ (
    .A(_7843_),
    .B(_7832_),
    .C(_7854_),
    .Y(_7898_)
);

AOI21X1 _12416_ (
    .A(_7810_),
    .B(_7777_),
    .C(_7635_),
    .Y(_7909_)
);

OAI21X1 _12417_ (
    .A(_7898_),
    .B(_7909_),
    .C(_7887_),
    .Y(_7920_)
);

NAND3X1 _12418_ (
    .A(_7876_),
    .B(_7920_),
    .C(_7547_),
    .Y(_7931_)
);

NAND3X1 _12419_ (
    .A(_7503_),
    .B(_7404_),
    .C(_7481_),
    .Y(_7942_)
);

NAND3X1 _12420_ (
    .A(_7316_),
    .B(_7514_),
    .C(_7525_),
    .Y(_7953_)
);

NAND2X1 _12421_ (
    .A(_7942_),
    .B(_7953_),
    .Y(_7964_)
);

NOR3X1 _12422_ (
    .A(_7898_),
    .B(_7909_),
    .C(_7887_),
    .Y(_7975_)
);

AOI21X1 _12423_ (
    .A(_7821_),
    .B(_7865_),
    .C(_7558_),
    .Y(_7986_)
);

OAI21X1 _12424_ (
    .A(_7975_),
    .B(_7986_),
    .C(_7964_),
    .Y(_7997_)
);

NAND3X1 _12425_ (
    .A(_7931_),
    .B(_7294_),
    .C(_7997_),
    .Y(_8008_)
);

AOI21X1 _12426_ (
    .A(_6769_),
    .B(_6341_),
    .C(_6802_),
    .Y(_8029_)
);

OAI21X1 _12427_ (
    .A(_7898_),
    .B(_7909_),
    .C(_7558_),
    .Y(_8040_)
);

NAND3X1 _12428_ (
    .A(_7821_),
    .B(_7865_),
    .C(_7887_),
    .Y(_8041_)
);

AOI21X1 _12429_ (
    .A(_8040_),
    .B(_8041_),
    .C(_7964_),
    .Y(_8052_)
);

AOI21X1 _12430_ (
    .A(_7876_),
    .B(_7920_),
    .C(_7547_),
    .Y(_8063_)
);

OAI21X1 _12431_ (
    .A(_8052_),
    .B(_8063_),
    .C(_8029_),
    .Y(_8073_)
);

NAND3X1 _12432_ (
    .A(_8073_),
    .B(_7283_),
    .C(_8008_),
    .Y(_8084_)
);

OAI21X1 _12433_ (
    .A(_8052_),
    .B(_8063_),
    .C(_7294_),
    .Y(_8095_)
);

NAND3X1 _12434_ (
    .A(_7931_),
    .B(_7997_),
    .C(_8029_),
    .Y(_8106_)
);

NAND3X1 _12435_ (
    .A(_7272_),
    .B(_8095_),
    .C(_8106_),
    .Y(_8117_)
);

NAND3X1 _12436_ (
    .A(_8084_),
    .B(_8117_),
    .C(_7196_),
    .Y(_8128_)
);

AOI21X1 _12437_ (
    .A(_6099_),
    .B(_6900_),
    .C(_6922_),
    .Y(_8139_)
);

AOI21X1 _12438_ (
    .A(_8095_),
    .B(_8106_),
    .C(_7272_),
    .Y(_8150_)
);

AOI21X1 _12439_ (
    .A(_8073_),
    .B(_8008_),
    .C(_7283_),
    .Y(_8161_)
);

OAI21X1 _12440_ (
    .A(_8150_),
    .B(_8161_),
    .C(_8139_),
    .Y(_8172_)
);

NAND3X1 _12441_ (
    .A(_7185_),
    .B(_8172_),
    .C(_8128_),
    .Y(_8183_)
);

INVX2 _12442_ (
    .A(_7185_),
    .Y(_8194_)
);

OAI21X1 _12443_ (
    .A(_8150_),
    .B(_8161_),
    .C(_7196_),
    .Y(_8205_)
);

NAND3X1 _12444_ (
    .A(_8084_),
    .B(_8117_),
    .C(_8139_),
    .Y(_8216_)
);

NAND3X1 _12445_ (
    .A(_8194_),
    .B(_8205_),
    .C(_8216_),
    .Y(_8227_)
);

AOI21X1 _12446_ (
    .A(_8183_),
    .B(_8227_),
    .C(_6955_),
    .Y(_8238_)
);

INVX2 _12447_ (
    .A(_6955_),
    .Y(_8249_)
);

NAND3X1 _12448_ (
    .A(_8194_),
    .B(_8172_),
    .C(_8128_),
    .Y(_8260_)
);

NAND3X1 _12449_ (
    .A(_7185_),
    .B(_8205_),
    .C(_8216_),
    .Y(_8271_)
);

AOI21X1 _12450_ (
    .A(_8260_),
    .B(_8271_),
    .C(_8249_),
    .Y(_8282_)
);

AOI21X1 _12451_ (
    .A(_7043_),
    .B(_6012_),
    .C(_7065_),
    .Y(_8293_)
);

OAI21X1 _12452_ (
    .A(_8238_),
    .B(_8282_),
    .C(_8293_),
    .Y(_8304_)
);

AOI21X1 _12453_ (
    .A(_8183_),
    .B(_8227_),
    .C(_8249_),
    .Y(_8315_)
);

AOI21X1 _12454_ (
    .A(_8260_),
    .B(_8271_),
    .C(_6955_),
    .Y(_8326_)
);

OAI21X1 _12455_ (
    .A(_5859_),
    .B(_7087_),
    .C(_7020_),
    .Y(_8337_)
);

OAI21X1 _12456_ (
    .A(_8315_),
    .B(_8326_),
    .C(_8337_),
    .Y(_8348_)
);

NAND2X1 _12457_ (
    .A(_8348_),
    .B(_8304_),
    .Y(_8359_)
);

OAI21X1 _12458_ (
    .A(_7164_),
    .B(_5947_),
    .C(_7109_),
    .Y(_8370_)
);

XNOR2X1 _12459_ (
    .A(_8370_),
    .B(_8359_),
    .Y(_0_[10])
);

NOR2X1 _12460_ (
    .A(_7109_),
    .B(_8359_),
    .Y(_8391_)
);

NOR3X1 _12461_ (
    .A(_5947_),
    .B(_8359_),
    .C(_7164_),
    .Y(_8402_)
);

NOR2X1 _12462_ (
    .A(_8391_),
    .B(_8402_),
    .Y(_8413_)
);

NOR2X1 _12463_ (
    .A(_7065_),
    .B(_7087_),
    .Y(_8424_)
);

NAND3X1 _12464_ (
    .A(_6955_),
    .B(_8260_),
    .C(_8271_),
    .Y(_8435_)
);

NAND3X1 _12465_ (
    .A(_8249_),
    .B(_8183_),
    .C(_8227_),
    .Y(_8446_)
);

NAND2X1 _12466_ (
    .A(_8435_),
    .B(_8446_),
    .Y(_8457_)
);

NAND3X1 _12467_ (
    .A(_6012_),
    .B(_8424_),
    .C(_8457_),
    .Y(_8467_)
);

AOI21X1 _12468_ (
    .A(_8435_),
    .B(_8446_),
    .C(_7020_),
    .Y(_8478_)
);

AOI21X1 _12469_ (
    .A(_8084_),
    .B(_8117_),
    .C(_7196_),
    .Y(_8489_)
);

OAI21X1 _12470_ (
    .A(_8489_),
    .B(_7185_),
    .C(_8128_),
    .Y(_8500_)
);

NAND2X1 _12471_ (
    .A(_7250_),
    .B(_7261_),
    .Y(_8511_)
);

INVX2 _12472_ (
    .A(_8511_),
    .Y(_8522_)
);

AOI21X1 _12473_ (
    .A(_7931_),
    .B(_7997_),
    .C(_7294_),
    .Y(_8533_)
);

OAI21X1 _12474_ (
    .A(_8533_),
    .B(_7272_),
    .C(_8008_),
    .Y(_8544_)
);

INVX4 _12475_ (
    .A(breg_11_bF$buf4),
    .Y(_8555_)
);

NOR2X1 _12476_ (
    .A(_2376__bF$buf2),
    .B(_8555_),
    .Y(_8566_)
);

INVX1 _12477_ (
    .A(_8566_),
    .Y(_8577_)
);

NAND2X1 _12478_ (
    .A(areg_2_bF$buf2),
    .B(breg_10_bF$buf3),
    .Y(_8588_)
);

NAND2X1 _12479_ (
    .A(areg_1_bF$buf3),
    .B(breg_10_bF$buf2),
    .Y(_8599_)
);

OAI21X1 _12480_ (
    .A(_2519__bF$buf2),
    .B(_6044__bF$buf4),
    .C(_8599_),
    .Y(_8610_)
);

OAI21X1 _12481_ (
    .A(_7228_),
    .B(_8588_),
    .C(_8610_),
    .Y(_8621_)
);

XNOR2X1 _12482_ (
    .A(_8621_),
    .B(_8577_),
    .Y(_8632_)
);

NAND2X1 _12483_ (
    .A(_7207_),
    .B(_8632_),
    .Y(_8643_)
);

NOR2X1 _12484_ (
    .A(_7207_),
    .B(_8632_),
    .Y(_8654_)
);

INVX2 _12485_ (
    .A(_8654_),
    .Y(_8665_)
);

NAND2X1 _12486_ (
    .A(_8643_),
    .B(_8665_),
    .Y(_8676_)
);

OAI21X1 _12487_ (
    .A(_7459_),
    .B(_7470_),
    .C(_7942_),
    .Y(_8687_)
);

XNOR2X1 _12488_ (
    .A(_8687_),
    .B(_8676_),
    .Y(_8698_)
);

OAI21X1 _12489_ (
    .A(_7964_),
    .B(_7986_),
    .C(_7876_),
    .Y(_8709_)
);

OAI21X1 _12490_ (
    .A(_6220_),
    .B(_7338_),
    .C(_7448_),
    .Y(_8720_)
);

INVX1 _12491_ (
    .A(_8720_),
    .Y(_8731_)
);

NAND2X1 _12492_ (
    .A(areg_3_bF$buf2),
    .B(breg[8]),
    .Y(_8742_)
);

NAND2X1 _12493_ (
    .A(areg_5_bF$buf4),
    .B(breg_6_bF$buf5),
    .Y(_8753_)
);

NOR2X1 _12494_ (
    .A(_7338_),
    .B(_8753_),
    .Y(_8764_)
);

AOI22X1 _12495_ (
    .A(areg_5_bF$buf3),
    .B(breg_6_bF$buf4),
    .C(areg_4_bF$buf2),
    .D(breg_7_bF$buf0),
    .Y(_8775_)
);

OAI21X1 _12496_ (
    .A(_8764_),
    .B(_8775_),
    .C(_8742_),
    .Y(_8786_)
);

INVX1 _12497_ (
    .A(_8742_),
    .Y(_8797_)
);

OR2X2 _12498_ (
    .A(_7338_),
    .B(_8753_),
    .Y(_8808_)
);

INVX1 _12499_ (
    .A(_8775_),
    .Y(_8819_)
);

NAND3X1 _12500_ (
    .A(_8797_),
    .B(_8819_),
    .C(_8808_),
    .Y(_8830_)
);

OAI22X1 _12501_ (
    .A(_6385_),
    .B(_7591_),
    .C(_7580_),
    .D(_7623_),
    .Y(_8851_)
);

AOI21X1 _12502_ (
    .A(_8786_),
    .B(_8830_),
    .C(_8851_),
    .Y(_8852_)
);

NAND2X1 _12503_ (
    .A(_8786_),
    .B(_8830_),
    .Y(_8863_)
);

AOI21X1 _12504_ (
    .A(_7569_),
    .B(_7624_),
    .C(_7602_),
    .Y(_8874_)
);

NOR2X1 _12505_ (
    .A(_8874_),
    .B(_8863_),
    .Y(_8884_)
);

OAI21X1 _12506_ (
    .A(_8884_),
    .B(_8852_),
    .C(_8731_),
    .Y(_8895_)
);

NAND2X1 _12507_ (
    .A(_8874_),
    .B(_8863_),
    .Y(_8906_)
);

NAND3X1 _12508_ (
    .A(_8786_),
    .B(_8830_),
    .C(_8851_),
    .Y(_8917_)
);

NAND3X1 _12509_ (
    .A(_8720_),
    .B(_8917_),
    .C(_8906_),
    .Y(_8928_)
);

NAND2X1 _12510_ (
    .A(_8928_),
    .B(_8895_),
    .Y(_8939_)
);

OAI21X1 _12511_ (
    .A(_7854_),
    .B(_7832_),
    .C(_7777_),
    .Y(_8950_)
);

NOR2X1 _12512_ (
    .A(_4258__bF$buf3),
    .B(_3646__bF$buf0),
    .Y(_8961_)
);

INVX2 _12513_ (
    .A(_8961_),
    .Y(_8972_)
);

NAND2X1 _12514_ (
    .A(breg_3_bF$buf4),
    .B(areg_8_bF$buf0),
    .Y(_8983_)
);

NOR2X1 _12515_ (
    .A(_7591_),
    .B(_8983_),
    .Y(_8994_)
);

AND2X2 _12516_ (
    .A(_7591_),
    .B(_8983_),
    .Y(_9005_)
);

NOR2X1 _12517_ (
    .A(_8994_),
    .B(_9005_),
    .Y(_9016_)
);

XNOR2X1 _12518_ (
    .A(_9016_),
    .B(_8972_),
    .Y(_9027_)
);

OAI21X1 _12519_ (
    .A(_7755_),
    .B(_7667_),
    .C(_7700_),
    .Y(_9038_)
);

NAND2X1 _12520_ (
    .A(breg_2_bF$buf1),
    .B(areg_9_bF$buf1),
    .Y(_9049_)
);

INVX2 _12521_ (
    .A(_9049_),
    .Y(_9060_)
);

AND2X2 _12522_ (
    .A(breg_1_bF$buf3),
    .B(areg_10_bF$buf2),
    .Y(_9071_)
);

AND2X2 _12523_ (
    .A(breg_0_bF$buf2),
    .B(areg_11_bF$buf4),
    .Y(_9092_)
);

NAND2X1 _12524_ (
    .A(_9071_),
    .B(_9092_),
    .Y(_9103_)
);

INVX8 _12525_ (
    .A(areg_11_bF$buf3),
    .Y(_9104_)
);

OAI22X1 _12526_ (
    .A(_2551__bF$buf0),
    .B(_9104__bF$buf3),
    .C(_3220_),
    .D(_7711__bF$buf2),
    .Y(_9115_)
);

NAND3X1 _12527_ (
    .A(_9060_),
    .B(_9115_),
    .C(_9103_),
    .Y(_9126_)
);

NAND2X1 _12528_ (
    .A(breg_1_bF$buf2),
    .B(areg_11_bF$buf2),
    .Y(_9137_)
);

NOR2X1 _12529_ (
    .A(_7689_),
    .B(_9137_),
    .Y(_9148_)
);

NOR2X1 _12530_ (
    .A(_9071_),
    .B(_9092_),
    .Y(_9159_)
);

OAI21X1 _12531_ (
    .A(_9159_),
    .B(_9148_),
    .C(_9049_),
    .Y(_9170_)
);

NAND3X1 _12532_ (
    .A(_9038_),
    .B(_9126_),
    .C(_9170_),
    .Y(_9181_)
);

AOI21X1 _12533_ (
    .A(_7678_),
    .B(_7722_),
    .C(_7744_),
    .Y(_9192_)
);

NOR3X1 _12534_ (
    .A(_9049_),
    .B(_9148_),
    .C(_9159_),
    .Y(_9203_)
);

AOI21X1 _12535_ (
    .A(_9115_),
    .B(_9103_),
    .C(_9060_),
    .Y(_9214_)
);

OAI21X1 _12536_ (
    .A(_9203_),
    .B(_9214_),
    .C(_9192_),
    .Y(_9225_)
);

NAND3X1 _12537_ (
    .A(_9181_),
    .B(_9225_),
    .C(_9027_),
    .Y(_9236_)
);

XNOR2X1 _12538_ (
    .A(_9016_),
    .B(_8961_),
    .Y(_9247_)
);

NOR3X1 _12539_ (
    .A(_9192_),
    .B(_9214_),
    .C(_9203_),
    .Y(_9257_)
);

AOI21X1 _12540_ (
    .A(_9126_),
    .B(_9170_),
    .C(_9038_),
    .Y(_9268_)
);

OAI21X1 _12541_ (
    .A(_9257_),
    .B(_9268_),
    .C(_9247_),
    .Y(_9279_)
);

AOI21X1 _12542_ (
    .A(_9236_),
    .B(_9279_),
    .C(_8950_),
    .Y(_9290_)
);

AOI21X1 _12543_ (
    .A(_7810_),
    .B(_7635_),
    .C(_7843_),
    .Y(_9301_)
);

OAI21X1 _12544_ (
    .A(_9203_),
    .B(_9214_),
    .C(_9038_),
    .Y(_9312_)
);

NAND3X1 _12545_ (
    .A(_9192_),
    .B(_9126_),
    .C(_9170_),
    .Y(_9323_)
);

AOI21X1 _12546_ (
    .A(_9312_),
    .B(_9323_),
    .C(_9247_),
    .Y(_9334_)
);

AOI21X1 _12547_ (
    .A(_9225_),
    .B(_9181_),
    .C(_9027_),
    .Y(_9345_)
);

NOR3X1 _12548_ (
    .A(_9334_),
    .B(_9301_),
    .C(_9345_),
    .Y(_9356_)
);

OAI21X1 _12549_ (
    .A(_9356_),
    .B(_9290_),
    .C(_8939_),
    .Y(_9367_)
);

AND2X2 _12550_ (
    .A(_8895_),
    .B(_8928_),
    .Y(_9378_)
);

OAI21X1 _12551_ (
    .A(_9334_),
    .B(_9345_),
    .C(_9301_),
    .Y(_9389_)
);

NAND3X1 _12552_ (
    .A(_9236_),
    .B(_8950_),
    .C(_9279_),
    .Y(_9400_)
);

NAND3X1 _12553_ (
    .A(_9389_),
    .B(_9400_),
    .C(_9378_),
    .Y(_9411_)
);

NAND3X1 _12554_ (
    .A(_9367_),
    .B(_9411_),
    .C(_8709_),
    .Y(_9422_)
);

AOI21X1 _12555_ (
    .A(_7920_),
    .B(_7547_),
    .C(_7975_),
    .Y(_9433_)
);

AOI21X1 _12556_ (
    .A(_9389_),
    .B(_9400_),
    .C(_9378_),
    .Y(_9444_)
);

NOR3X1 _12557_ (
    .A(_8939_),
    .B(_9290_),
    .C(_9356_),
    .Y(_9455_)
);

OAI21X1 _12558_ (
    .A(_9455_),
    .B(_9444_),
    .C(_9433_),
    .Y(_9466_)
);

NAND3X1 _12559_ (
    .A(_8698_),
    .B(_9422_),
    .C(_9466_),
    .Y(_9477_)
);

XOR2X1 _12560_ (
    .A(_8687_),
    .B(_8676_),
    .Y(_9488_)
);

OAI21X1 _12561_ (
    .A(_9455_),
    .B(_9444_),
    .C(_8709_),
    .Y(_9499_)
);

NAND3X1 _12562_ (
    .A(_9411_),
    .B(_9367_),
    .C(_9433_),
    .Y(_9510_)
);

NAND3X1 _12563_ (
    .A(_9488_),
    .B(_9510_),
    .C(_9499_),
    .Y(_9521_)
);

NAND3X1 _12564_ (
    .A(_9477_),
    .B(_9521_),
    .C(_8544_),
    .Y(_9532_)
);

NOR3X1 _12565_ (
    .A(_8052_),
    .B(_8063_),
    .C(_8029_),
    .Y(_9543_)
);

AOI21X1 _12566_ (
    .A(_7283_),
    .B(_8073_),
    .C(_9543_),
    .Y(_9554_)
);

AOI21X1 _12567_ (
    .A(_9510_),
    .B(_9499_),
    .C(_9488_),
    .Y(_9565_)
);

AOI21X1 _12568_ (
    .A(_9422_),
    .B(_9466_),
    .C(_8698_),
    .Y(_9576_)
);

OAI21X1 _12569_ (
    .A(_9565_),
    .B(_9576_),
    .C(_9554_),
    .Y(_9587_)
);

NAND3X1 _12570_ (
    .A(_8522_),
    .B(_9587_),
    .C(_9532_),
    .Y(_9598_)
);

OAI21X1 _12571_ (
    .A(_9565_),
    .B(_9576_),
    .C(_8544_),
    .Y(_9609_)
);

NAND3X1 _12572_ (
    .A(_9477_),
    .B(_9521_),
    .C(_9554_),
    .Y(_9620_)
);

NAND3X1 _12573_ (
    .A(_8511_),
    .B(_9609_),
    .C(_9620_),
    .Y(_9631_)
);

NAND3X1 _12574_ (
    .A(_9598_),
    .B(_9631_),
    .C(_8500_),
    .Y(_9641_)
);

NOR3X1 _12575_ (
    .A(_8150_),
    .B(_8161_),
    .C(_8139_),
    .Y(_9652_)
);

AOI21X1 _12576_ (
    .A(_8194_),
    .B(_8172_),
    .C(_9652_),
    .Y(_9663_)
);

AOI21X1 _12577_ (
    .A(_9609_),
    .B(_9620_),
    .C(_8511_),
    .Y(_9674_)
);

AOI21X1 _12578_ (
    .A(_9587_),
    .B(_9532_),
    .C(_8522_),
    .Y(_9685_)
);

OAI21X1 _12579_ (
    .A(_9674_),
    .B(_9685_),
    .C(_9663_),
    .Y(_9696_)
);

NAND3X1 _12580_ (
    .A(_9641_),
    .B(_8238_),
    .C(_9696_),
    .Y(_9707_)
);

NAND3X1 _12581_ (
    .A(_8249_),
    .B(_8260_),
    .C(_8271_),
    .Y(_9718_)
);

OAI21X1 _12582_ (
    .A(_9674_),
    .B(_9685_),
    .C(_8500_),
    .Y(_9729_)
);

NAND3X1 _12583_ (
    .A(_9598_),
    .B(_9631_),
    .C(_9663_),
    .Y(_9740_)
);

NAND3X1 _12584_ (
    .A(_9718_),
    .B(_9729_),
    .C(_9740_),
    .Y(_9751_)
);

NAND3X1 _12585_ (
    .A(_8478_),
    .B(_9707_),
    .C(_9751_),
    .Y(_9762_)
);

NAND3X1 _12586_ (
    .A(_6955_),
    .B(_8183_),
    .C(_8227_),
    .Y(_9773_)
);

NAND3X1 _12587_ (
    .A(_7065_),
    .B(_9718_),
    .C(_9773_),
    .Y(_9784_)
);

NAND3X1 _12588_ (
    .A(_9718_),
    .B(_9641_),
    .C(_9696_),
    .Y(_9795_)
);

NAND3X1 _12589_ (
    .A(_8238_),
    .B(_9729_),
    .C(_9740_),
    .Y(_9806_)
);

NAND3X1 _12590_ (
    .A(_9784_),
    .B(_9795_),
    .C(_9806_),
    .Y(_9817_)
);

NAND3X1 _12591_ (
    .A(_8467_),
    .B(_9817_),
    .C(_9762_),
    .Y(_9828_)
);

AOI21X1 _12592_ (
    .A(_8435_),
    .B(_8446_),
    .C(_7054_),
    .Y(_9839_)
);

NAND3X1 _12593_ (
    .A(_9784_),
    .B(_9707_),
    .C(_9751_),
    .Y(_9850_)
);

NAND3X1 _12594_ (
    .A(_8478_),
    .B(_9795_),
    .C(_9806_),
    .Y(_9861_)
);

NAND3X1 _12595_ (
    .A(_9839_),
    .B(_9850_),
    .C(_9861_),
    .Y(_9872_)
);

NAND2X1 _12596_ (
    .A(_9828_),
    .B(_9872_),
    .Y(_9883_)
);

XNOR2X1 _12597_ (
    .A(_8413_),
    .B(_9883_),
    .Y(_0_[11])
);

NAND3X1 _12598_ (
    .A(_8467_),
    .B(_9850_),
    .C(_9861_),
    .Y(_9904_)
);

NAND3X1 _12599_ (
    .A(_9839_),
    .B(_9817_),
    .C(_9762_),
    .Y(_9915_)
);

OAI21X1 _12600_ (
    .A(_7109_),
    .B(_8359_),
    .C(_9915_),
    .Y(_9926_)
);

AOI22X1 _12601_ (
    .A(_9883_),
    .B(_8402_),
    .C(_9904_),
    .D(_9926_),
    .Y(_9937_)
);

AOI21X1 _12602_ (
    .A(_9729_),
    .B(_9740_),
    .C(_9718_),
    .Y(_9948_)
);

INVX1 _12603_ (
    .A(_9641_),
    .Y(_9959_)
);

AOI21X1 _12604_ (
    .A(_9477_),
    .B(_9521_),
    .C(_8544_),
    .Y(_9970_)
);

OAI21X1 _12605_ (
    .A(_9970_),
    .B(_8511_),
    .C(_9532_),
    .Y(_9981_)
);

INVX1 _12606_ (
    .A(_8676_),
    .Y(_9991_)
);

NAND2X1 _12607_ (
    .A(_8687_),
    .B(_9991_),
    .Y(_10002_)
);

AOI21X1 _12608_ (
    .A(_9367_),
    .B(_9411_),
    .C(_8709_),
    .Y(_10013_)
);

OAI21X1 _12609_ (
    .A(_10013_),
    .B(_9488_),
    .C(_9422_),
    .Y(_10024_)
);

NAND2X1 _12610_ (
    .A(areg[0]),
    .B(breg_12_bF$buf4),
    .Y(_10035_)
);

NAND2X1 _12611_ (
    .A(areg_2_bF$buf1),
    .B(breg_9_bF$buf3),
    .Y(_10046_)
);

NOR2X1 _12612_ (
    .A(_8599_),
    .B(_10046_),
    .Y(_10057_)
);

AOI21X1 _12613_ (
    .A(_8566_),
    .B(_8610_),
    .C(_10057_),
    .Y(_10068_)
);

INVX1 _12614_ (
    .A(_10068_),
    .Y(_10079_)
);

NOR2X1 _12615_ (
    .A(_2661_),
    .B(_8555_),
    .Y(_10090_)
);

INVX1 _12616_ (
    .A(_10090_),
    .Y(_10101_)
);

NAND2X1 _12617_ (
    .A(areg_3_bF$buf1),
    .B(breg_9_bF$buf2),
    .Y(_10112_)
);

NOR2X1 _12618_ (
    .A(_8588_),
    .B(_10112_),
    .Y(_10123_)
);

AOI22X1 _12619_ (
    .A(areg_3_bF$buf0),
    .B(breg_9_bF$buf1),
    .C(areg_2_bF$buf0),
    .D(breg_10_bF$buf1),
    .Y(_10134_)
);

OAI21X1 _12620_ (
    .A(_10123_),
    .B(_10134_),
    .C(_10101_),
    .Y(_10145_)
);

NOR2X1 _12621_ (
    .A(_10134_),
    .B(_10123_),
    .Y(_10156_)
);

NAND2X1 _12622_ (
    .A(_10090_),
    .B(_10156_),
    .Y(_10167_)
);

AOI21X1 _12623_ (
    .A(_10145_),
    .B(_10167_),
    .C(_10079_),
    .Y(_10178_)
);

NOR2X1 _12624_ (
    .A(_10090_),
    .B(_10156_),
    .Y(_10189_)
);

NAND2X1 _12625_ (
    .A(areg_3_bF$buf4),
    .B(breg_10_bF$buf0),
    .Y(_10200_)
);

OAI21X1 _12626_ (
    .A(_2519__bF$buf1),
    .B(_7217__bF$buf3),
    .C(_10112_),
    .Y(_10221_)
);

OAI21X1 _12627_ (
    .A(_10046_),
    .B(_10200_),
    .C(_10221_),
    .Y(_10232_)
);

NOR2X1 _12628_ (
    .A(_10101_),
    .B(_10232_),
    .Y(_10233_)
);

NOR3X1 _12629_ (
    .A(_10233_),
    .B(_10068_),
    .C(_10189_),
    .Y(_10244_)
);

OAI21X1 _12630_ (
    .A(_10244_),
    .B(_10178_),
    .C(_10035_),
    .Y(_10255_)
);

INVX1 _12631_ (
    .A(_10035_),
    .Y(_10266_)
);

OAI21X1 _12632_ (
    .A(_10189_),
    .B(_10233_),
    .C(_10068_),
    .Y(_10277_)
);

NAND3X1 _12633_ (
    .A(_10145_),
    .B(_10079_),
    .C(_10167_),
    .Y(_10288_)
);

NAND3X1 _12634_ (
    .A(_10266_),
    .B(_10288_),
    .C(_10277_),
    .Y(_10299_)
);

OAI21X1 _12635_ (
    .A(_8731_),
    .B(_8852_),
    .C(_8917_),
    .Y(_10310_)
);

AOI21X1 _12636_ (
    .A(_10299_),
    .B(_10255_),
    .C(_10310_),
    .Y(_10321_)
);

AOI21X1 _12637_ (
    .A(_10288_),
    .B(_10277_),
    .C(_10266_),
    .Y(_10332_)
);

NOR3X1 _12638_ (
    .A(_10035_),
    .B(_10178_),
    .C(_10244_),
    .Y(_10342_)
);

AOI21X1 _12639_ (
    .A(_8720_),
    .B(_8906_),
    .C(_8884_),
    .Y(_10353_)
);

NOR3X1 _12640_ (
    .A(_10332_),
    .B(_10353_),
    .C(_10342_),
    .Y(_10364_)
);

OAI21X1 _12641_ (
    .A(_10364_),
    .B(_10321_),
    .C(_8665_),
    .Y(_10375_)
);

OAI21X1 _12642_ (
    .A(_10342_),
    .B(_10332_),
    .C(_10353_),
    .Y(_10386_)
);

NAND3X1 _12643_ (
    .A(_10299_),
    .B(_10310_),
    .C(_10255_),
    .Y(_10397_)
);

NAND3X1 _12644_ (
    .A(_8654_),
    .B(_10397_),
    .C(_10386_),
    .Y(_10408_)
);

NAND2X1 _12645_ (
    .A(_10408_),
    .B(_10375_),
    .Y(_10419_)
);

OAI21X1 _12646_ (
    .A(_8939_),
    .B(_9290_),
    .C(_9400_),
    .Y(_10430_)
);

OAI21X1 _12647_ (
    .A(_8742_),
    .B(_8775_),
    .C(_8808_),
    .Y(_10441_)
);

NAND2X1 _12648_ (
    .A(areg_6_bF$buf3),
    .B(breg_7_bF$buf5),
    .Y(_10452_)
);

NAND2X1 _12649_ (
    .A(areg_6_bF$buf2),
    .B(breg_6_bF$buf3),
    .Y(_10463_)
);

OAI21X1 _12650_ (
    .A(_2825__bF$buf0),
    .B(_4116__bF$buf3),
    .C(_10463_),
    .Y(_10474_)
);

OAI21X1 _12651_ (
    .A(_8753_),
    .B(_10452_),
    .C(_10474_),
    .Y(_10485_)
);

OAI21X1 _12652_ (
    .A(_2562__bF$buf0),
    .B(_5420__bF$buf2),
    .C(_10485_),
    .Y(_10496_)
);

NOR2X1 _12653_ (
    .A(_2562__bF$buf4),
    .B(_5420__bF$buf1),
    .Y(_10507_)
);

NAND2X1 _12654_ (
    .A(areg_5_bF$buf2),
    .B(breg_7_bF$buf4),
    .Y(_10518_)
);

XOR2X1 _12655_ (
    .A(_10518_),
    .B(_10463_),
    .Y(_10529_)
);

NAND2X1 _12656_ (
    .A(_10507_),
    .B(_10529_),
    .Y(_10540_)
);

INVX1 _12657_ (
    .A(_8994_),
    .Y(_10551_)
);

OAI21X1 _12658_ (
    .A(_8972_),
    .B(_9005_),
    .C(_10551_),
    .Y(_10562_)
);

NAND3X1 _12659_ (
    .A(_10562_),
    .B(_10496_),
    .C(_10540_),
    .Y(_10573_)
);

NOR2X1 _12660_ (
    .A(_10507_),
    .B(_10529_),
    .Y(_10584_)
);

AND2X2 _12661_ (
    .A(_10529_),
    .B(_10507_),
    .Y(_10595_)
);

INVX1 _12662_ (
    .A(_9005_),
    .Y(_10606_)
);

AOI21X1 _12663_ (
    .A(_8961_),
    .B(_10606_),
    .C(_8994_),
    .Y(_10617_)
);

OAI21X1 _12664_ (
    .A(_10595_),
    .B(_10584_),
    .C(_10617_),
    .Y(_10628_)
);

NAND3X1 _12665_ (
    .A(_10441_),
    .B(_10573_),
    .C(_10628_),
    .Y(_10639_)
);

INVX1 _12666_ (
    .A(_10441_),
    .Y(_10650_)
);

NAND3X1 _12667_ (
    .A(_10496_),
    .B(_10540_),
    .C(_10617_),
    .Y(_10661_)
);

OAI21X1 _12668_ (
    .A(_10595_),
    .B(_10584_),
    .C(_10562_),
    .Y(_10671_)
);

NAND3X1 _12669_ (
    .A(_10650_),
    .B(_10661_),
    .C(_10671_),
    .Y(_10682_)
);

NAND2X1 _12670_ (
    .A(_10639_),
    .B(_10682_),
    .Y(_10693_)
);

OAI21X1 _12671_ (
    .A(_9247_),
    .B(_9268_),
    .C(_9181_),
    .Y(_10704_)
);

NOR2X1 _12672_ (
    .A(_4258__bF$buf2),
    .B(_4434__bF$buf1),
    .Y(_10715_)
);

INVX2 _12673_ (
    .A(_10715_),
    .Y(_10726_)
);

NAND2X1 _12674_ (
    .A(breg_4_bF$buf2),
    .B(areg_8_bF$buf4),
    .Y(_10737_)
);

NAND2X1 _12675_ (
    .A(breg_3_bF$buf3),
    .B(areg_9_bF$buf0),
    .Y(_10748_)
);

NOR2X1 _12676_ (
    .A(_10737_),
    .B(_10748_),
    .Y(_10759_)
);

AND2X2 _12677_ (
    .A(_10737_),
    .B(_10748_),
    .Y(_10770_)
);

NOR2X1 _12678_ (
    .A(_10759_),
    .B(_10770_),
    .Y(_10781_)
);

XNOR2X1 _12679_ (
    .A(_10781_),
    .B(_10726_),
    .Y(_10792_)
);

OAI21X1 _12680_ (
    .A(_9159_),
    .B(_9049_),
    .C(_9103_),
    .Y(_10803_)
);

NAND2X1 _12681_ (
    .A(breg_2_bF$buf0),
    .B(areg_10_bF$buf1),
    .Y(_10814_)
);

INVX2 _12682_ (
    .A(_10814_),
    .Y(_10825_)
);

AND2X2 _12683_ (
    .A(breg_1_bF$buf1),
    .B(areg_11_bF$buf1),
    .Y(_10836_)
);

AND2X2 _12684_ (
    .A(breg_0_bF$buf1),
    .B(areg_12_bF$buf4),
    .Y(_10847_)
);

NAND2X1 _12685_ (
    .A(_10836_),
    .B(_10847_),
    .Y(_10858_)
);

INVX8 _12686_ (
    .A(areg_12_bF$buf3),
    .Y(_10869_)
);

OAI21X1 _12687_ (
    .A(_2551__bF$buf3),
    .B(_10869__bF$buf3),
    .C(_9137_),
    .Y(_10880_)
);

NAND3X1 _12688_ (
    .A(_10825_),
    .B(_10880_),
    .C(_10858_),
    .Y(_10891_)
);

NAND2X1 _12689_ (
    .A(breg_0_bF$buf0),
    .B(areg_12_bF$buf2),
    .Y(_10902_)
);

NOR2X1 _12690_ (
    .A(_9137_),
    .B(_10902_),
    .Y(_10913_)
);

NOR2X1 _12691_ (
    .A(_10836_),
    .B(_10847_),
    .Y(_10924_)
);

OAI21X1 _12692_ (
    .A(_10924_),
    .B(_10913_),
    .C(_10814_),
    .Y(_10935_)
);

NAND3X1 _12693_ (
    .A(_10891_),
    .B(_10803_),
    .C(_10935_),
    .Y(_10946_)
);

AOI21X1 _12694_ (
    .A(_9060_),
    .B(_9115_),
    .C(_9148_),
    .Y(_10957_)
);

NOR3X1 _12695_ (
    .A(_10814_),
    .B(_10913_),
    .C(_10924_),
    .Y(_10968_)
);

AOI21X1 _12696_ (
    .A(_10880_),
    .B(_10858_),
    .C(_10825_),
    .Y(_10979_)
);

OAI21X1 _12697_ (
    .A(_10968_),
    .B(_10979_),
    .C(_10957_),
    .Y(_10990_)
);

NAND3X1 _12698_ (
    .A(_10946_),
    .B(_10990_),
    .C(_10792_),
    .Y(_11000_)
);

XNOR2X1 _12699_ (
    .A(_10781_),
    .B(_10715_),
    .Y(_11011_)
);

NOR3X1 _12700_ (
    .A(_10957_),
    .B(_10979_),
    .C(_10968_),
    .Y(_11022_)
);

AOI21X1 _12701_ (
    .A(_10891_),
    .B(_10935_),
    .C(_10803_),
    .Y(_11043_)
);

OAI21X1 _12702_ (
    .A(_11022_),
    .B(_11043_),
    .C(_11011_),
    .Y(_11044_)
);

AOI21X1 _12703_ (
    .A(_11000_),
    .B(_11044_),
    .C(_10704_),
    .Y(_11055_)
);

AOI21X1 _12704_ (
    .A(_9225_),
    .B(_9027_),
    .C(_9257_),
    .Y(_11066_)
);

OAI21X1 _12705_ (
    .A(_10968_),
    .B(_10979_),
    .C(_10803_),
    .Y(_11077_)
);

NAND3X1 _12706_ (
    .A(_10957_),
    .B(_10891_),
    .C(_10935_),
    .Y(_11088_)
);

AOI21X1 _12707_ (
    .A(_11077_),
    .B(_11088_),
    .C(_11011_),
    .Y(_11099_)
);

AOI21X1 _12708_ (
    .A(_10990_),
    .B(_10946_),
    .C(_10792_),
    .Y(_11110_)
);

NOR3X1 _12709_ (
    .A(_11099_),
    .B(_11110_),
    .C(_11066_),
    .Y(_11121_)
);

OAI21X1 _12710_ (
    .A(_11121_),
    .B(_11055_),
    .C(_10693_),
    .Y(_11132_)
);

AND2X2 _12711_ (
    .A(_10639_),
    .B(_10682_),
    .Y(_11143_)
);

OAI21X1 _12712_ (
    .A(_11099_),
    .B(_11110_),
    .C(_11066_),
    .Y(_11154_)
);

NAND3X1 _12713_ (
    .A(_11000_),
    .B(_11044_),
    .C(_10704_),
    .Y(_11165_)
);

NAND3X1 _12714_ (
    .A(_11154_),
    .B(_11165_),
    .C(_11143_),
    .Y(_11176_)
);

AOI21X1 _12715_ (
    .A(_11132_),
    .B(_11176_),
    .C(_10430_),
    .Y(_11187_)
);

AOI21X1 _12716_ (
    .A(_9389_),
    .B(_9378_),
    .C(_9356_),
    .Y(_11198_)
);

AOI21X1 _12717_ (
    .A(_11154_),
    .B(_11165_),
    .C(_11143_),
    .Y(_11209_)
);

NOR3X1 _12718_ (
    .A(_10693_),
    .B(_11055_),
    .C(_11121_),
    .Y(_11220_)
);

NOR3X1 _12719_ (
    .A(_11198_),
    .B(_11209_),
    .C(_11220_),
    .Y(_11231_)
);

OAI21X1 _12720_ (
    .A(_11231_),
    .B(_11187_),
    .C(_10419_),
    .Y(_11242_)
);

AND2X2 _12721_ (
    .A(_10375_),
    .B(_10408_),
    .Y(_11253_)
);

OAI21X1 _12722_ (
    .A(_11220_),
    .B(_11209_),
    .C(_11198_),
    .Y(_11264_)
);

NAND3X1 _12723_ (
    .A(_10430_),
    .B(_11132_),
    .C(_11176_),
    .Y(_11275_)
);

NAND3X1 _12724_ (
    .A(_11264_),
    .B(_11275_),
    .C(_11253_),
    .Y(_11286_)
);

AOI21X1 _12725_ (
    .A(_11242_),
    .B(_11286_),
    .C(_10024_),
    .Y(_11297_)
);

NOR3X1 _12726_ (
    .A(_9455_),
    .B(_9444_),
    .C(_9433_),
    .Y(_11308_)
);

AOI21X1 _12727_ (
    .A(_8698_),
    .B(_9466_),
    .C(_11308_),
    .Y(_11318_)
);

AOI21X1 _12728_ (
    .A(_11264_),
    .B(_11275_),
    .C(_11253_),
    .Y(_11329_)
);

NOR3X1 _12729_ (
    .A(_10419_),
    .B(_11187_),
    .C(_11231_),
    .Y(_11350_)
);

NOR3X1 _12730_ (
    .A(_11329_),
    .B(_11318_),
    .C(_11350_),
    .Y(_11361_)
);

OAI21X1 _12731_ (
    .A(_11361_),
    .B(_11297_),
    .C(_10002_),
    .Y(_11362_)
);

INVX2 _12732_ (
    .A(_10002_),
    .Y(_11373_)
);

OAI21X1 _12733_ (
    .A(_11350_),
    .B(_11329_),
    .C(_11318_),
    .Y(_11384_)
);

NAND3X1 _12734_ (
    .A(_10024_),
    .B(_11242_),
    .C(_11286_),
    .Y(_11395_)
);

NAND3X1 _12735_ (
    .A(_11373_),
    .B(_11395_),
    .C(_11384_),
    .Y(_11406_)
);

NAND3X1 _12736_ (
    .A(_9981_),
    .B(_11406_),
    .C(_11362_),
    .Y(_11417_)
);

NAND2X1 _12737_ (
    .A(_9477_),
    .B(_9521_),
    .Y(_11428_)
);

NOR2X1 _12738_ (
    .A(_9554_),
    .B(_11428_),
    .Y(_11439_)
);

AOI21X1 _12739_ (
    .A(_8522_),
    .B(_9587_),
    .C(_11439_),
    .Y(_11450_)
);

AOI21X1 _12740_ (
    .A(_11395_),
    .B(_11384_),
    .C(_11373_),
    .Y(_11461_)
);

NOR3X1 _12741_ (
    .A(_10002_),
    .B(_11297_),
    .C(_11361_),
    .Y(_11472_)
);

OAI21X1 _12742_ (
    .A(_11472_),
    .B(_11461_),
    .C(_11450_),
    .Y(_11483_)
);

NAND3X1 _12743_ (
    .A(_11417_),
    .B(_11483_),
    .C(_9959_),
    .Y(_11494_)
);

OAI21X1 _12744_ (
    .A(_11472_),
    .B(_11461_),
    .C(_9981_),
    .Y(_11505_)
);

NAND3X1 _12745_ (
    .A(_11406_),
    .B(_11450_),
    .C(_11362_),
    .Y(_11516_)
);

NAND3X1 _12746_ (
    .A(_9641_),
    .B(_11516_),
    .C(_11505_),
    .Y(_11527_)
);

NAND3X1 _12747_ (
    .A(_9948_),
    .B(_11527_),
    .C(_11494_),
    .Y(_11538_)
);

AOI21X1 _12748_ (
    .A(_11516_),
    .B(_11505_),
    .C(_9641_),
    .Y(_11549_)
);

AOI21X1 _12749_ (
    .A(_11417_),
    .B(_11483_),
    .C(_9959_),
    .Y(_11560_)
);

OAI21X1 _12750_ (
    .A(_11549_),
    .B(_11560_),
    .C(_9707_),
    .Y(_11571_)
);

NAND3X1 _12751_ (
    .A(_9762_),
    .B(_11538_),
    .C(_11571_),
    .Y(_11582_)
);

INVX1 _12752_ (
    .A(_9762_),
    .Y(_11592_)
);

NAND3X1 _12753_ (
    .A(_9707_),
    .B(_11527_),
    .C(_11494_),
    .Y(_11603_)
);

OAI21X1 _12754_ (
    .A(_11549_),
    .B(_11560_),
    .C(_9948_),
    .Y(_11614_)
);

NAND3X1 _12755_ (
    .A(_11603_),
    .B(_11614_),
    .C(_11592_),
    .Y(_11625_)
);

NAND2X1 _12756_ (
    .A(_11582_),
    .B(_11625_),
    .Y(_11636_)
);

XNOR2X1 _12757_ (
    .A(_9937_),
    .B(_11636_),
    .Y(_0_[12])
);

OAI21X1 _12758_ (
    .A(_11297_),
    .B(_10002_),
    .C(_11395_),
    .Y(_11657_)
);

OAI21X1 _12759_ (
    .A(_10321_),
    .B(_8665_),
    .C(_10397_),
    .Y(_11668_)
);

OAI21X1 _12760_ (
    .A(_10419_),
    .B(_11187_),
    .C(_11275_),
    .Y(_11679_)
);

OAI21X1 _12761_ (
    .A(_10178_),
    .B(_10035_),
    .C(_10288_),
    .Y(_11690_)
);

INVX1 _12762_ (
    .A(_11690_),
    .Y(_11701_)
);

NAND2X1 _12763_ (
    .A(areg_1_bF$buf2),
    .B(breg_13_bF$buf4),
    .Y(_11712_)
);

NOR2X1 _12764_ (
    .A(_10035_),
    .B(_11712_),
    .Y(_11723_)
);

AOI22X1 _12765_ (
    .A(areg_1_bF$buf1),
    .B(breg_12_bF$buf3),
    .C(areg[0]),
    .D(breg_13_bF$buf3),
    .Y(_11734_)
);

NOR2X1 _12766_ (
    .A(_11734_),
    .B(_11723_),
    .Y(_11745_)
);

NOR2X1 _12767_ (
    .A(_2519__bF$buf0),
    .B(_8555_),
    .Y(_11756_)
);

NAND2X1 _12768_ (
    .A(areg_4_bF$buf1),
    .B(breg_10_bF$buf5),
    .Y(_11767_)
);

OAI21X1 _12769_ (
    .A(_2562__bF$buf3),
    .B(_6044__bF$buf3),
    .C(_10200_),
    .Y(_11778_)
);

OAI21X1 _12770_ (
    .A(_10112_),
    .B(_11767_),
    .C(_11778_),
    .Y(_11789_)
);

XNOR2X1 _12771_ (
    .A(_11789_),
    .B(_11756_),
    .Y(_11800_)
);

OAI21X1 _12772_ (
    .A(_10123_),
    .B(_10233_),
    .C(_11800_),
    .Y(_11811_)
);

AOI21X1 _12773_ (
    .A(_10090_),
    .B(_10221_),
    .C(_10123_),
    .Y(_11822_)
);

INVX1 _12774_ (
    .A(_11756_),
    .Y(_11833_)
);

XNOR2X1 _12775_ (
    .A(_11789_),
    .B(_11833_),
    .Y(_11844_)
);

NAND2X1 _12776_ (
    .A(_11822_),
    .B(_11844_),
    .Y(_11855_)
);

NAND3X1 _12777_ (
    .A(_11745_),
    .B(_11855_),
    .C(_11811_),
    .Y(_11866_)
);

INVX1 _12778_ (
    .A(_11745_),
    .Y(_11876_)
);

OAI21X1 _12779_ (
    .A(_10123_),
    .B(_10233_),
    .C(_11844_),
    .Y(_11887_)
);

NAND2X1 _12780_ (
    .A(_11822_),
    .B(_11800_),
    .Y(_11898_)
);

NAND3X1 _12781_ (
    .A(_11876_),
    .B(_11898_),
    .C(_11887_),
    .Y(_1_)
);

AOI21X1 _12782_ (
    .A(_10496_),
    .B(_10540_),
    .C(_10562_),
    .Y(_12_)
);

OAI21X1 _12783_ (
    .A(_12_),
    .B(_10650_),
    .C(_10573_),
    .Y(_23_)
);

NAND3X1 _12784_ (
    .A(_23_),
    .B(_11866_),
    .C(_1_),
    .Y(_34_)
);

AOI21X1 _12785_ (
    .A(_11898_),
    .B(_11887_),
    .C(_11876_),
    .Y(_45_)
);

AOI21X1 _12786_ (
    .A(_11855_),
    .B(_11811_),
    .C(_11745_),
    .Y(_56_)
);

INVX1 _12787_ (
    .A(_23_),
    .Y(_67_)
);

OAI21X1 _12788_ (
    .A(_45_),
    .B(_56_),
    .C(_67_),
    .Y(_78_)
);

NAND3X1 _12789_ (
    .A(_11701_),
    .B(_34_),
    .C(_78_),
    .Y(_89_)
);

NAND3X1 _12790_ (
    .A(_11866_),
    .B(_1_),
    .C(_67_),
    .Y(_100_)
);

OAI21X1 _12791_ (
    .A(_45_),
    .B(_56_),
    .C(_23_),
    .Y(_111_)
);

NAND3X1 _12792_ (
    .A(_11690_),
    .B(_111_),
    .C(_100_),
    .Y(_122_)
);

NAND2X1 _12793_ (
    .A(_89_),
    .B(_122_),
    .Y(_133_)
);

OAI21X1 _12794_ (
    .A(_10693_),
    .B(_11055_),
    .C(_11165_),
    .Y(_144_)
);

OAI21X1 _12795_ (
    .A(_10518_),
    .B(_10463_),
    .C(_10540_),
    .Y(_155_)
);

NOR2X1 _12796_ (
    .A(_2825__bF$buf4),
    .B(_5420__bF$buf0),
    .Y(_166_)
);

NAND2X1 _12797_ (
    .A(areg_7_bF$buf4),
    .B(breg_7_bF$buf3),
    .Y(_177_)
);

OAI21X1 _12798_ (
    .A(_5453__bF$buf2),
    .B(_4434__bF$buf0),
    .C(_10452_),
    .Y(_188_)
);

OAI21X1 _12799_ (
    .A(_10463_),
    .B(_177_),
    .C(_188_),
    .Y(_199_)
);

XNOR2X1 _12800_ (
    .A(_199_),
    .B(_166_),
    .Y(_210_)
);

NAND2X1 _12801_ (
    .A(breg_4_bF$buf1),
    .B(areg_9_bF$buf4),
    .Y(_221_)
);

OAI22X1 _12802_ (
    .A(_8983_),
    .B(_221_),
    .C(_10726_),
    .D(_10770_),
    .Y(_232_)
);

NAND2X1 _12803_ (
    .A(_232_),
    .B(_210_),
    .Y(_242_)
);

NAND2X1 _12804_ (
    .A(breg_6_bF$buf2),
    .B(areg_7_bF$buf3),
    .Y(_253_)
);

XOR2X1 _12805_ (
    .A(_10452_),
    .B(_253_),
    .Y(_264_)
);

NOR2X1 _12806_ (
    .A(_166_),
    .B(_264_),
    .Y(_275_)
);

AND2X2 _12807_ (
    .A(_264_),
    .B(_166_),
    .Y(_286_)
);

INVX1 _12808_ (
    .A(_232_),
    .Y(_297_)
);

OAI21X1 _12809_ (
    .A(_286_),
    .B(_275_),
    .C(_297_),
    .Y(_308_)
);

NAND3X1 _12810_ (
    .A(_155_),
    .B(_308_),
    .C(_242_),
    .Y(_319_)
);

NOR2X1 _12811_ (
    .A(_10518_),
    .B(_10463_),
    .Y(_330_)
);

NOR2X1 _12812_ (
    .A(_330_),
    .B(_10595_),
    .Y(_341_)
);

NAND2X1 _12813_ (
    .A(_297_),
    .B(_210_),
    .Y(_352_)
);

OAI21X1 _12814_ (
    .A(_286_),
    .B(_275_),
    .C(_232_),
    .Y(_373_)
);

NAND3X1 _12815_ (
    .A(_341_),
    .B(_373_),
    .C(_352_),
    .Y(_374_)
);

NAND2X1 _12816_ (
    .A(_319_),
    .B(_374_),
    .Y(_385_)
);

OAI21X1 _12817_ (
    .A(_11011_),
    .B(_11043_),
    .C(_10946_),
    .Y(_396_)
);

NOR2X1 _12818_ (
    .A(_4258__bF$buf1),
    .B(_5190__bF$buf2),
    .Y(_407_)
);

INVX2 _12819_ (
    .A(_407_),
    .Y(_418_)
);

NAND2X1 _12820_ (
    .A(breg_3_bF$buf2),
    .B(areg_10_bF$buf0),
    .Y(_429_)
);

NOR2X1 _12821_ (
    .A(_221_),
    .B(_429_),
    .Y(_440_)
);

AND2X2 _12822_ (
    .A(_221_),
    .B(_429_),
    .Y(_451_)
);

NOR2X1 _12823_ (
    .A(_440_),
    .B(_451_),
    .Y(_462_)
);

XNOR2X1 _12824_ (
    .A(_462_),
    .B(_418_),
    .Y(_473_)
);

AOI21X1 _12825_ (
    .A(_10825_),
    .B(_10880_),
    .C(_10913_),
    .Y(_484_)
);

INVX2 _12826_ (
    .A(_484_),
    .Y(_494_)
);

NOR2X1 _12827_ (
    .A(_2508_),
    .B(_9104__bF$buf2),
    .Y(_505_)
);

NAND2X1 _12828_ (
    .A(breg_1_bF$buf0),
    .B(areg_12_bF$buf1),
    .Y(_516_)
);

NAND2X1 _12829_ (
    .A(breg_0_bF$buf6),
    .B(areg_13_bF$buf4),
    .Y(_527_)
);

OR2X2 _12830_ (
    .A(_516_),
    .B(_527_),
    .Y(_538_)
);

INVX8 _12831_ (
    .A(areg_13_bF$buf3),
    .Y(_549_)
);

OAI21X1 _12832_ (
    .A(_2551__bF$buf2),
    .B(_549__bF$buf4),
    .C(_516_),
    .Y(_560_)
);

NAND3X1 _12833_ (
    .A(_505_),
    .B(_560_),
    .C(_538_),
    .Y(_571_)
);

NAND2X1 _12834_ (
    .A(breg_1_bF$buf6),
    .B(areg_13_bF$buf2),
    .Y(_582_)
);

OAI21X1 _12835_ (
    .A(_10902_),
    .B(_582_),
    .C(_560_),
    .Y(_593_)
);

OAI21X1 _12836_ (
    .A(_2508_),
    .B(_9104__bF$buf1),
    .C(_593_),
    .Y(_604_)
);

NAND3X1 _12837_ (
    .A(_571_),
    .B(_604_),
    .C(_494_),
    .Y(_615_)
);

INVX1 _12838_ (
    .A(_505_),
    .Y(_626_)
);

NOR2X1 _12839_ (
    .A(_626_),
    .B(_593_),
    .Y(_637_)
);

AOI21X1 _12840_ (
    .A(_560_),
    .B(_538_),
    .C(_505_),
    .Y(_648_)
);

OAI21X1 _12841_ (
    .A(_637_),
    .B(_648_),
    .C(_484_),
    .Y(_659_)
);

NAND3X1 _12842_ (
    .A(_473_),
    .B(_615_),
    .C(_659_),
    .Y(_680_)
);

XNOR2X1 _12843_ (
    .A(_462_),
    .B(_407_),
    .Y(_691_)
);

NOR3X1 _12844_ (
    .A(_648_),
    .B(_484_),
    .C(_637_),
    .Y(_692_)
);

AOI21X1 _12845_ (
    .A(_571_),
    .B(_604_),
    .C(_494_),
    .Y(_703_)
);

OAI21X1 _12846_ (
    .A(_692_),
    .B(_703_),
    .C(_691_),
    .Y(_713_)
);

AOI21X1 _12847_ (
    .A(_680_),
    .B(_713_),
    .C(_396_),
    .Y(_724_)
);

AOI21X1 _12848_ (
    .A(_10990_),
    .B(_10792_),
    .C(_11022_),
    .Y(_735_)
);

OAI21X1 _12849_ (
    .A(_637_),
    .B(_648_),
    .C(_494_),
    .Y(_746_)
);

NAND3X1 _12850_ (
    .A(_484_),
    .B(_571_),
    .C(_604_),
    .Y(_757_)
);

AOI21X1 _12851_ (
    .A(_757_),
    .B(_746_),
    .C(_691_),
    .Y(_768_)
);

AOI21X1 _12852_ (
    .A(_615_),
    .B(_659_),
    .C(_473_),
    .Y(_779_)
);

NOR3X1 _12853_ (
    .A(_768_),
    .B(_735_),
    .C(_779_),
    .Y(_790_)
);

OAI21X1 _12854_ (
    .A(_790_),
    .B(_724_),
    .C(_385_),
    .Y(_801_)
);

AND2X2 _12855_ (
    .A(_319_),
    .B(_374_),
    .Y(_812_)
);

OAI21X1 _12856_ (
    .A(_768_),
    .B(_779_),
    .C(_735_),
    .Y(_823_)
);

NAND3X1 _12857_ (
    .A(_396_),
    .B(_680_),
    .C(_713_),
    .Y(_834_)
);

NAND3X1 _12858_ (
    .A(_823_),
    .B(_834_),
    .C(_812_),
    .Y(_845_)
);

NAND3X1 _12859_ (
    .A(_144_),
    .B(_801_),
    .C(_845_),
    .Y(_856_)
);

AOI21X1 _12860_ (
    .A(_11154_),
    .B(_11143_),
    .C(_11121_),
    .Y(_867_)
);

AOI21X1 _12861_ (
    .A(_823_),
    .B(_834_),
    .C(_812_),
    .Y(_878_)
);

NOR3X1 _12862_ (
    .A(_724_),
    .B(_385_),
    .C(_790_),
    .Y(_889_)
);

OAI21X1 _12863_ (
    .A(_889_),
    .B(_878_),
    .C(_867_),
    .Y(_900_)
);

NAND3X1 _12864_ (
    .A(_133_),
    .B(_856_),
    .C(_900_),
    .Y(_911_)
);

AND2X2 _12865_ (
    .A(_122_),
    .B(_89_),
    .Y(_921_)
);

NOR3X1 _12866_ (
    .A(_878_),
    .B(_867_),
    .C(_889_),
    .Y(_932_)
);

AOI21X1 _12867_ (
    .A(_801_),
    .B(_845_),
    .C(_144_),
    .Y(_943_)
);

OAI21X1 _12868_ (
    .A(_932_),
    .B(_943_),
    .C(_921_),
    .Y(_954_)
);

NAND3X1 _12869_ (
    .A(_11679_),
    .B(_911_),
    .C(_954_),
    .Y(_965_)
);

AOI21X1 _12870_ (
    .A(_11264_),
    .B(_11253_),
    .C(_11231_),
    .Y(_976_)
);

OAI21X1 _12871_ (
    .A(_889_),
    .B(_878_),
    .C(_144_),
    .Y(_987_)
);

NAND3X1 _12872_ (
    .A(_867_),
    .B(_801_),
    .C(_845_),
    .Y(_998_)
);

AOI21X1 _12873_ (
    .A(_998_),
    .B(_987_),
    .C(_921_),
    .Y(_1009_)
);

AOI21X1 _12874_ (
    .A(_856_),
    .B(_900_),
    .C(_133_),
    .Y(_1020_)
);

OAI21X1 _12875_ (
    .A(_1009_),
    .B(_1020_),
    .C(_976_),
    .Y(_1031_)
);

NAND3X1 _12876_ (
    .A(_11668_),
    .B(_1031_),
    .C(_965_),
    .Y(_1042_)
);

INVX1 _12877_ (
    .A(_11668_),
    .Y(_1053_)
);

OAI21X1 _12878_ (
    .A(_1009_),
    .B(_1020_),
    .C(_11679_),
    .Y(_1064_)
);

NAND3X1 _12879_ (
    .A(_911_),
    .B(_954_),
    .C(_976_),
    .Y(_1075_)
);

NAND3X1 _12880_ (
    .A(_1053_),
    .B(_1064_),
    .C(_1075_),
    .Y(_1086_)
);

NAND3X1 _12881_ (
    .A(_1042_),
    .B(_1086_),
    .C(_11657_),
    .Y(_1096_)
);

AOI21X1 _12882_ (
    .A(_11373_),
    .B(_11384_),
    .C(_11361_),
    .Y(_1107_)
);

AOI21X1 _12883_ (
    .A(_1064_),
    .B(_1075_),
    .C(_1053_),
    .Y(_1118_)
);

AOI21X1 _12884_ (
    .A(_1031_),
    .B(_965_),
    .C(_11668_),
    .Y(_1129_)
);

OAI21X1 _12885_ (
    .A(_1118_),
    .B(_1129_),
    .C(_1107_),
    .Y(_1140_)
);

NAND3X1 _12886_ (
    .A(_1096_),
    .B(_1140_),
    .C(_11417_),
    .Y(_1151_)
);

NOR3X1 _12887_ (
    .A(_11450_),
    .B(_11461_),
    .C(_11472_),
    .Y(_1162_)
);

NOR3X1 _12888_ (
    .A(_1118_),
    .B(_1129_),
    .C(_1107_),
    .Y(_1173_)
);

AOI21X1 _12889_ (
    .A(_1042_),
    .B(_1086_),
    .C(_11657_),
    .Y(_1184_)
);

OAI21X1 _12890_ (
    .A(_1173_),
    .B(_1184_),
    .C(_1162_),
    .Y(_1195_)
);

NAND2X1 _12891_ (
    .A(_1151_),
    .B(_1195_),
    .Y(_1206_)
);

AOI21X1 _12892_ (
    .A(_9948_),
    .B(_11527_),
    .C(_11549_),
    .Y(_1217_)
);

XNOR2X1 _12893_ (
    .A(_1217_),
    .B(_1206_),
    .Y(_1228_)
);

AOI21X1 _12894_ (
    .A(_9850_),
    .B(_9861_),
    .C(_8467_),
    .Y(_1239_)
);

OAI21X1 _12895_ (
    .A(_8391_),
    .B(_1239_),
    .C(_9904_),
    .Y(_1250_)
);

NAND3X1 _12896_ (
    .A(_9915_),
    .B(_9904_),
    .C(_8402_),
    .Y(_1260_)
);

NAND2X1 _12897_ (
    .A(_1250_),
    .B(_1260_),
    .Y(_1271_)
);

AOI21X1 _12898_ (
    .A(_11603_),
    .B(_11614_),
    .C(_9762_),
    .Y(_1282_)
);

AOI21X1 _12899_ (
    .A(_11636_),
    .B(_1271_),
    .C(_1282_),
    .Y(_1293_)
);

XNOR2X1 _12900_ (
    .A(_1293_),
    .B(_1228_),
    .Y(_0_[13])
);

AOI21X1 _12901_ (
    .A(_11603_),
    .B(_11614_),
    .C(_11592_),
    .Y(_1314_)
);

AOI21X1 _12902_ (
    .A(_11538_),
    .B(_11571_),
    .C(_9762_),
    .Y(_1325_)
);

AND2X2 _12903_ (
    .A(_1195_),
    .B(_1151_),
    .Y(_1336_)
);

OAI21X1 _12904_ (
    .A(_11560_),
    .B(_9707_),
    .C(_11494_),
    .Y(_1347_)
);

NOR2X1 _12905_ (
    .A(_1336_),
    .B(_1347_),
    .Y(_1358_)
);

NOR2X1 _12906_ (
    .A(_1206_),
    .B(_1217_),
    .Y(_1369_)
);

OAI22X1 _12907_ (
    .A(_1369_),
    .B(_1358_),
    .C(_1314_),
    .D(_1325_),
    .Y(_1380_)
);

NOR2X1 _12908_ (
    .A(_11538_),
    .B(_1336_),
    .Y(_1391_)
);

AOI21X1 _12909_ (
    .A(_1282_),
    .B(_1228_),
    .C(_1391_),
    .Y(_1401_)
);

OAI21X1 _12910_ (
    .A(_9937_),
    .B(_1380_),
    .C(_1401_),
    .Y(_1412_)
);

NAND2X1 _12911_ (
    .A(_965_),
    .B(_1042_),
    .Y(_1423_)
);

NAND2X1 _12912_ (
    .A(_34_),
    .B(_78_),
    .Y(_1434_)
);

OAI21X1 _12913_ (
    .A(_1434_),
    .B(_11701_),
    .C(_34_),
    .Y(_1445_)
);

XNOR2X1 _12914_ (
    .A(_1445_),
    .B(_11723_),
    .Y(_1456_)
);

INVX2 _12915_ (
    .A(_1456_),
    .Y(_1467_)
);

OAI21X1 _12916_ (
    .A(_921_),
    .B(_943_),
    .C(_856_),
    .Y(_1478_)
);

AND2X2 _12917_ (
    .A(_11866_),
    .B(_11811_),
    .Y(_1489_)
);

NAND2X1 _12918_ (
    .A(areg[0]),
    .B(breg_14_bF$buf3),
    .Y(_1500_)
);

NAND2X1 _12919_ (
    .A(areg_2_bF$buf4),
    .B(breg_12_bF$buf2),
    .Y(_1511_)
);

XOR2X1 _12920_ (
    .A(_11712_),
    .B(_1511_),
    .Y(_1522_)
);

XNOR2X1 _12921_ (
    .A(_1522_),
    .B(_1500_),
    .Y(_1533_)
);

NOR2X1 _12922_ (
    .A(_10112_),
    .B(_11767_),
    .Y(_1543_)
);

AOI21X1 _12923_ (
    .A(_11756_),
    .B(_11778_),
    .C(_1543_),
    .Y(_1554_)
);

INVX2 _12924_ (
    .A(_1554_),
    .Y(_1565_)
);

NOR2X1 _12925_ (
    .A(_2792_),
    .B(_8555_),
    .Y(_1586_)
);

NAND2X1 _12926_ (
    .A(areg_4_bF$buf0),
    .B(breg_9_bF$buf0),
    .Y(_1587_)
);

NAND2X1 _12927_ (
    .A(areg_5_bF$buf1),
    .B(breg_10_bF$buf4),
    .Y(_1598_)
);

OAI21X1 _12928_ (
    .A(_2825__bF$buf3),
    .B(_6044__bF$buf2),
    .C(_11767_),
    .Y(_1609_)
);

OAI21X1 _12929_ (
    .A(_1587_),
    .B(_1598_),
    .C(_1609_),
    .Y(_1620_)
);

XNOR2X1 _12930_ (
    .A(_1620_),
    .B(_1586_),
    .Y(_1631_)
);

NAND2X1 _12931_ (
    .A(_1565_),
    .B(_1631_),
    .Y(_1642_)
);

INVX1 _12932_ (
    .A(_1586_),
    .Y(_1653_)
);

XNOR2X1 _12933_ (
    .A(_1620_),
    .B(_1653_),
    .Y(_1663_)
);

NAND2X1 _12934_ (
    .A(_1554_),
    .B(_1663_),
    .Y(_1674_)
);

NAND3X1 _12935_ (
    .A(_1533_),
    .B(_1642_),
    .C(_1674_),
    .Y(_1685_)
);

INVX1 _12936_ (
    .A(_1533_),
    .Y(_1696_)
);

NAND2X1 _12937_ (
    .A(_1565_),
    .B(_1663_),
    .Y(_1707_)
);

NAND2X1 _12938_ (
    .A(_1554_),
    .B(_1631_),
    .Y(_1718_)
);

NAND3X1 _12939_ (
    .A(_1696_),
    .B(_1707_),
    .C(_1718_),
    .Y(_1729_)
);

NOR2X1 _12940_ (
    .A(_232_),
    .B(_210_),
    .Y(_1740_)
);

OAI21X1 _12941_ (
    .A(_1740_),
    .B(_341_),
    .C(_242_),
    .Y(_1751_)
);

NAND3X1 _12942_ (
    .A(_1685_),
    .B(_1729_),
    .C(_1751_),
    .Y(_1762_)
);

AOI21X1 _12943_ (
    .A(_1718_),
    .B(_1707_),
    .C(_1696_),
    .Y(_1772_)
);

AOI21X1 _12944_ (
    .A(_1642_),
    .B(_1674_),
    .C(_1533_),
    .Y(_1783_)
);

AND2X2 _12945_ (
    .A(_210_),
    .B(_232_),
    .Y(_1794_)
);

AOI21X1 _12946_ (
    .A(_155_),
    .B(_308_),
    .C(_1794_),
    .Y(_1805_)
);

OAI21X1 _12947_ (
    .A(_1772_),
    .B(_1783_),
    .C(_1805_),
    .Y(_1816_)
);

NAND3X1 _12948_ (
    .A(_1489_),
    .B(_1816_),
    .C(_1762_),
    .Y(_1827_)
);

OAI21X1 _12949_ (
    .A(_11822_),
    .B(_11844_),
    .C(_11866_),
    .Y(_1838_)
);

NAND3X1 _12950_ (
    .A(_1685_),
    .B(_1729_),
    .C(_1805_),
    .Y(_1849_)
);

OAI21X1 _12951_ (
    .A(_1772_),
    .B(_1783_),
    .C(_1751_),
    .Y(_1860_)
);

NAND3X1 _12952_ (
    .A(_1838_),
    .B(_1860_),
    .C(_1849_),
    .Y(_1870_)
);

NAND2X1 _12953_ (
    .A(_1827_),
    .B(_1870_),
    .Y(_1881_)
);

OAI21X1 _12954_ (
    .A(_724_),
    .B(_385_),
    .C(_834_),
    .Y(_1902_)
);

NOR2X1 _12955_ (
    .A(_10463_),
    .B(_177_),
    .Y(_1913_)
);

OR2X2 _12956_ (
    .A(_286_),
    .B(_1913_),
    .Y(_1914_)
);

NOR2X1 _12957_ (
    .A(_3646__bF$buf3),
    .B(_5420__bF$buf3),
    .Y(_1925_)
);

NAND2X1 _12958_ (
    .A(breg_7_bF$buf2),
    .B(areg_8_bF$buf3),
    .Y(_1936_)
);

OAI21X1 _12959_ (
    .A(_5453__bF$buf1),
    .B(_5190__bF$buf1),
    .C(_177_),
    .Y(_1947_)
);

OAI21X1 _12960_ (
    .A(_253_),
    .B(_1936_),
    .C(_1947_),
    .Y(_1957_)
);

XNOR2X1 _12961_ (
    .A(_1957_),
    .B(_1925_),
    .Y(_1968_)
);

NAND2X1 _12962_ (
    .A(breg_4_bF$buf0),
    .B(areg_10_bF$buf4),
    .Y(_1979_)
);

OAI22X1 _12963_ (
    .A(_10748_),
    .B(_1979_),
    .C(_418_),
    .D(_451_),
    .Y(_1990_)
);

NAND2X1 _12964_ (
    .A(_1990_),
    .B(_1968_),
    .Y(_2001_)
);

NAND2X1 _12965_ (
    .A(breg_6_bF$buf1),
    .B(areg_8_bF$buf2),
    .Y(_2012_)
);

XOR2X1 _12966_ (
    .A(_177_),
    .B(_2012_),
    .Y(_2023_)
);

AND2X2 _12967_ (
    .A(_2023_),
    .B(_1925_),
    .Y(_2034_)
);

NOR2X1 _12968_ (
    .A(_1925_),
    .B(_2023_),
    .Y(_2045_)
);

INVX1 _12969_ (
    .A(_1990_),
    .Y(_2055_)
);

OAI21X1 _12970_ (
    .A(_2034_),
    .B(_2045_),
    .C(_2055_),
    .Y(_2066_)
);

NAND3X1 _12971_ (
    .A(_2066_),
    .B(_1914_),
    .C(_2001_),
    .Y(_2077_)
);

NOR2X1 _12972_ (
    .A(_1913_),
    .B(_286_),
    .Y(_2088_)
);

NAND2X1 _12973_ (
    .A(_2055_),
    .B(_1968_),
    .Y(_2099_)
);

OAI21X1 _12974_ (
    .A(_2034_),
    .B(_2045_),
    .C(_1990_),
    .Y(_2109_)
);

NAND3X1 _12975_ (
    .A(_2088_),
    .B(_2109_),
    .C(_2099_),
    .Y(_2120_)
);

NAND2X1 _12976_ (
    .A(_2077_),
    .B(_2120_),
    .Y(_2131_)
);

OAI21X1 _12977_ (
    .A(_703_),
    .B(_691_),
    .C(_615_),
    .Y(_2142_)
);

NOR2X1 _12978_ (
    .A(_4258__bF$buf0),
    .B(_6582__bF$buf2),
    .Y(_2153_)
);

INVX2 _12979_ (
    .A(_2153_),
    .Y(_2163_)
);

NAND2X1 _12980_ (
    .A(breg_3_bF$buf1),
    .B(areg_11_bF$buf0),
    .Y(_2174_)
);

NOR2X1 _12981_ (
    .A(_1979_),
    .B(_2174_),
    .Y(_2185_)
);

AND2X2 _12982_ (
    .A(_1979_),
    .B(_2174_),
    .Y(_2196_)
);

NOR2X1 _12983_ (
    .A(_2185_),
    .B(_2196_),
    .Y(_2207_)
);

XNOR2X1 _12984_ (
    .A(_2207_),
    .B(_2163_),
    .Y(_2217_)
);

NOR2X1 _12985_ (
    .A(_516_),
    .B(_527_),
    .Y(_2228_)
);

AOI21X1 _12986_ (
    .A(_505_),
    .B(_560_),
    .C(_2228_),
    .Y(_2238_)
);

INVX2 _12987_ (
    .A(_2238_),
    .Y(_2249_)
);

NAND2X1 _12988_ (
    .A(breg_2_bF$buf4),
    .B(areg_12_bF$buf0),
    .Y(_2259_)
);

INVX2 _12989_ (
    .A(_2259_),
    .Y(_2270_)
);

NAND2X1 _12990_ (
    .A(breg_0_bF$buf5),
    .B(areg_14_bF$buf4),
    .Y(_2280_)
);

OR2X2 _12991_ (
    .A(_582_),
    .B(_2280_),
    .Y(_2286_)
);

INVX8 _12992_ (
    .A(areg_14_bF$buf3),
    .Y(_2287_)
);

OAI21X1 _12993_ (
    .A(_2551__bF$buf1),
    .B(_2287__bF$buf3),
    .C(_582_),
    .Y(_2288_)
);

NAND3X1 _12994_ (
    .A(_2270_),
    .B(_2288_),
    .C(_2286_),
    .Y(_2289_)
);

NOR2X1 _12995_ (
    .A(_582_),
    .B(_2280_),
    .Y(_2290_)
);

AND2X2 _12996_ (
    .A(_582_),
    .B(_2280_),
    .Y(_2291_)
);

OAI21X1 _12997_ (
    .A(_2291_),
    .B(_2290_),
    .C(_2259_),
    .Y(_2292_)
);

NAND3X1 _12998_ (
    .A(_2289_),
    .B(_2292_),
    .C(_2249_),
    .Y(_2293_)
);

NAND2X1 _12999_ (
    .A(breg_1_bF$buf5),
    .B(areg_14_bF$buf2),
    .Y(_2294_)
);

OAI21X1 _13000_ (
    .A(_527_),
    .B(_2294_),
    .C(_2288_),
    .Y(_2295_)
);

NOR2X1 _13001_ (
    .A(_2259_),
    .B(_2295_),
    .Y(_2296_)
);

AOI21X1 _13002_ (
    .A(_2288_),
    .B(_2286_),
    .C(_2270_),
    .Y(_2297_)
);

OAI21X1 _13003_ (
    .A(_2296_),
    .B(_2297_),
    .C(_2238_),
    .Y(_2298_)
);

NAND3X1 _13004_ (
    .A(_2217_),
    .B(_2293_),
    .C(_2298_),
    .Y(_2299_)
);

XNOR2X1 _13005_ (
    .A(_2207_),
    .B(_2153_),
    .Y(_2300_)
);

NAND2X1 _13006_ (
    .A(_2292_),
    .B(_2289_),
    .Y(_2301_)
);

NOR2X1 _13007_ (
    .A(_2238_),
    .B(_2301_),
    .Y(_2302_)
);

AOI21X1 _13008_ (
    .A(_2292_),
    .B(_2289_),
    .C(_2249_),
    .Y(_2303_)
);

OAI21X1 _13009_ (
    .A(_2302_),
    .B(_2303_),
    .C(_2300_),
    .Y(_2304_)
);

AOI21X1 _13010_ (
    .A(_2299_),
    .B(_2304_),
    .C(_2142_),
    .Y(_2305_)
);

AOI21X1 _13011_ (
    .A(_473_),
    .B(_659_),
    .C(_692_),
    .Y(_2306_)
);

OAI21X1 _13012_ (
    .A(_2296_),
    .B(_2297_),
    .C(_2249_),
    .Y(_2307_)
);

NAND3X1 _13013_ (
    .A(_2238_),
    .B(_2292_),
    .C(_2289_),
    .Y(_2308_)
);

AOI21X1 _13014_ (
    .A(_2308_),
    .B(_2307_),
    .C(_2300_),
    .Y(_2309_)
);

AOI21X1 _13015_ (
    .A(_2293_),
    .B(_2298_),
    .C(_2217_),
    .Y(_2310_)
);

NOR3X1 _13016_ (
    .A(_2309_),
    .B(_2310_),
    .C(_2306_),
    .Y(_2311_)
);

OAI21X1 _13017_ (
    .A(_2311_),
    .B(_2305_),
    .C(_2131_),
    .Y(_2312_)
);

AND2X2 _13018_ (
    .A(_2077_),
    .B(_2120_),
    .Y(_2313_)
);

OAI21X1 _13019_ (
    .A(_2309_),
    .B(_2310_),
    .C(_2306_),
    .Y(_2314_)
);

NAND3X1 _13020_ (
    .A(_2299_),
    .B(_2142_),
    .C(_2304_),
    .Y(_2315_)
);

NAND3X1 _13021_ (
    .A(_2314_),
    .B(_2315_),
    .C(_2313_),
    .Y(_2316_)
);

NAND3X1 _13022_ (
    .A(_1902_),
    .B(_2312_),
    .C(_2316_),
    .Y(_2317_)
);

AOI21X1 _13023_ (
    .A(_823_),
    .B(_812_),
    .C(_790_),
    .Y(_2318_)
);

AOI21X1 _13024_ (
    .A(_2314_),
    .B(_2315_),
    .C(_2313_),
    .Y(_2319_)
);

NOR3X1 _13025_ (
    .A(_2305_),
    .B(_2131_),
    .C(_2311_),
    .Y(_2320_)
);

OAI21X1 _13026_ (
    .A(_2320_),
    .B(_2319_),
    .C(_2318_),
    .Y(_2321_)
);

NAND3X1 _13027_ (
    .A(_1881_),
    .B(_2317_),
    .C(_2321_),
    .Y(_2322_)
);

AND2X2 _13028_ (
    .A(_1827_),
    .B(_1870_),
    .Y(_2323_)
);

OAI21X1 _13029_ (
    .A(_2320_),
    .B(_2319_),
    .C(_1902_),
    .Y(_2324_)
);

NAND3X1 _13030_ (
    .A(_2312_),
    .B(_2316_),
    .C(_2318_),
    .Y(_2325_)
);

NAND3X1 _13031_ (
    .A(_2325_),
    .B(_2324_),
    .C(_2323_),
    .Y(_2326_)
);

NAND3X1 _13032_ (
    .A(_2322_),
    .B(_2326_),
    .C(_1478_),
    .Y(_2327_)
);

AOI21X1 _13033_ (
    .A(_133_),
    .B(_900_),
    .C(_932_),
    .Y(_2328_)
);

AOI21X1 _13034_ (
    .A(_2325_),
    .B(_2324_),
    .C(_2323_),
    .Y(_2329_)
);

AOI21X1 _13035_ (
    .A(_2317_),
    .B(_2321_),
    .C(_1881_),
    .Y(_2330_)
);

OAI21X1 _13036_ (
    .A(_2329_),
    .B(_2330_),
    .C(_2328_),
    .Y(_2331_)
);

NAND3X1 _13037_ (
    .A(_1467_),
    .B(_2327_),
    .C(_2331_),
    .Y(_2332_)
);

NOR3X1 _13038_ (
    .A(_2329_),
    .B(_2328_),
    .C(_2330_),
    .Y(_2333_)
);

AOI21X1 _13039_ (
    .A(_2322_),
    .B(_2326_),
    .C(_1478_),
    .Y(_2334_)
);

OAI21X1 _13040_ (
    .A(_2333_),
    .B(_2334_),
    .C(_1456_),
    .Y(_2335_)
);

NAND3X1 _13041_ (
    .A(_2332_),
    .B(_2335_),
    .C(_1423_),
    .Y(_2336_)
);

AND2X2 _13042_ (
    .A(_1042_),
    .B(_965_),
    .Y(_2337_)
);

INVX1 _13043_ (
    .A(_2332_),
    .Y(_2338_)
);

AOI21X1 _13044_ (
    .A(_2327_),
    .B(_2331_),
    .C(_1467_),
    .Y(_2339_)
);

OAI21X1 _13045_ (
    .A(_2338_),
    .B(_2339_),
    .C(_2337_),
    .Y(_2340_)
);

NAND3X1 _13046_ (
    .A(_1173_),
    .B(_2336_),
    .C(_2340_),
    .Y(_2341_)
);

OAI21X1 _13047_ (
    .A(_2338_),
    .B(_2339_),
    .C(_1423_),
    .Y(_2342_)
);

NAND3X1 _13048_ (
    .A(_2332_),
    .B(_2335_),
    .C(_2337_),
    .Y(_2343_)
);

NAND3X1 _13049_ (
    .A(_1096_),
    .B(_2342_),
    .C(_2343_),
    .Y(_2344_)
);

NAND2X1 _13050_ (
    .A(_2341_),
    .B(_2344_),
    .Y(_2345_)
);

NAND3X1 _13051_ (
    .A(_1096_),
    .B(_1140_),
    .C(_1162_),
    .Y(_2346_)
);

AOI21X1 _13052_ (
    .A(_1096_),
    .B(_1140_),
    .C(_1162_),
    .Y(_2347_)
);

OAI21X1 _13053_ (
    .A(_2347_),
    .B(_11494_),
    .C(_2346_),
    .Y(_2348_)
);

OR2X2 _13054_ (
    .A(_2345_),
    .B(_2348_),
    .Y(_2349_)
);

AOI21X1 _13055_ (
    .A(_2342_),
    .B(_2343_),
    .C(_1096_),
    .Y(_2350_)
);

AOI21X1 _13056_ (
    .A(_2336_),
    .B(_2340_),
    .C(_1173_),
    .Y(_2351_)
);

OAI21X1 _13057_ (
    .A(_2350_),
    .B(_2351_),
    .C(_2348_),
    .Y(_2352_)
);

NAND2X1 _13058_ (
    .A(_2352_),
    .B(_2349_),
    .Y(_2353_)
);

XOR2X1 _13059_ (
    .A(_1412_),
    .B(_2353_),
    .Y(_0_[14])
);

NAND2X1 _13060_ (
    .A(_11549_),
    .B(_1206_),
    .Y(_2354_)
);

NOR2X1 _13061_ (
    .A(_2345_),
    .B(_2354_),
    .Y(_2355_)
);

AOI21X1 _13062_ (
    .A(_2353_),
    .B(_1412_),
    .C(_2355_),
    .Y(_2356_)
);

NAND2X1 _13063_ (
    .A(_2332_),
    .B(_2335_),
    .Y(_2357_)
);

NOR2X1 _13064_ (
    .A(_2337_),
    .B(_2357_),
    .Y(_2358_)
);

NAND2X1 _13065_ (
    .A(_11723_),
    .B(_1445_),
    .Y(_2359_)
);

INVX2 _13066_ (
    .A(_2359_),
    .Y(_2360_)
);

OAI21X1 _13067_ (
    .A(_2334_),
    .B(_1456_),
    .C(_2327_),
    .Y(_2361_)
);

INVX8 _13068_ (
    .A(breg_15_bF$buf5),
    .Y(_2362_)
);

NOR2X1 _13069_ (
    .A(_2376__bF$buf1),
    .B(_2362__bF$buf5),
    .Y(_2363_)
);

NAND3X1 _13070_ (
    .A(areg[0]),
    .B(breg_14_bF$buf2),
    .C(_1522_),
    .Y(_2364_)
);

OAI21X1 _13071_ (
    .A(_11712_),
    .B(_1511_),
    .C(_2364_),
    .Y(_2366_)
);

NOR2X1 _13072_ (
    .A(_2363_),
    .B(_2366_),
    .Y(_2367_)
);

NAND2X1 _13073_ (
    .A(_2363_),
    .B(_2366_),
    .Y(_2368_)
);

INVX1 _13074_ (
    .A(_2368_),
    .Y(_2369_)
);

NOR2X1 _13075_ (
    .A(_2367_),
    .B(_2369_),
    .Y(_2370_)
);

NAND2X1 _13076_ (
    .A(_1816_),
    .B(_1762_),
    .Y(_2371_)
);

OAI21X1 _13077_ (
    .A(_2371_),
    .B(_1489_),
    .C(_1762_),
    .Y(_2372_)
);

XNOR2X1 _13078_ (
    .A(_2372_),
    .B(_2370_),
    .Y(_2373_)
);

INVX2 _13079_ (
    .A(_2373_),
    .Y(_2374_)
);

AOI21X1 _13080_ (
    .A(_2312_),
    .B(_2316_),
    .C(_1902_),
    .Y(_2375_)
);

OAI21X1 _13081_ (
    .A(_2323_),
    .B(_2375_),
    .C(_2317_),
    .Y(_2377_)
);

AOI21X1 _13082_ (
    .A(_1565_),
    .B(_1631_),
    .C(_1772_),
    .Y(_2378_)
);

INVX4 _13083_ (
    .A(breg_14_bF$buf1),
    .Y(_2379_)
);

AOI22X1 _13084_ (
    .A(areg_3_bF$buf3),
    .B(breg_12_bF$buf1),
    .C(areg_2_bF$buf3),
    .D(breg_13_bF$buf2),
    .Y(_2380_)
);

NAND2X1 _13085_ (
    .A(areg_3_bF$buf2),
    .B(breg_13_bF$buf1),
    .Y(_2381_)
);

NOR2X1 _13086_ (
    .A(_1511_),
    .B(_2381_),
    .Y(_2382_)
);

OAI22X1 _13087_ (
    .A(_2661_),
    .B(_2379_),
    .C(_2382_),
    .D(_2380_),
    .Y(_2383_)
);

NOR2X1 _13088_ (
    .A(_2380_),
    .B(_2382_),
    .Y(_2384_)
);

NAND3X1 _13089_ (
    .A(areg_1_bF$buf0),
    .B(breg_14_bF$buf0),
    .C(_2384_),
    .Y(_2385_)
);

AND2X2 _13090_ (
    .A(_2385_),
    .B(_2383_),
    .Y(_2386_)
);

NAND2X1 _13091_ (
    .A(areg_5_bF$buf0),
    .B(breg_9_bF$buf5),
    .Y(_2388_)
);

NOR2X1 _13092_ (
    .A(_11767_),
    .B(_2388_),
    .Y(_2389_)
);

AOI21X1 _13093_ (
    .A(_1586_),
    .B(_1609_),
    .C(_2389_),
    .Y(_2390_)
);

INVX2 _13094_ (
    .A(_2390_),
    .Y(_2391_)
);

NOR2X1 _13095_ (
    .A(_2562__bF$buf2),
    .B(_8555_),
    .Y(_2392_)
);

NAND2X1 _13096_ (
    .A(areg_6_bF$buf1),
    .B(breg_10_bF$buf3),
    .Y(_2393_)
);

OAI21X1 _13097_ (
    .A(_3646__bF$buf2),
    .B(_6044__bF$buf1),
    .C(_1598_),
    .Y(_2394_)
);

OAI21X1 _13098_ (
    .A(_2388_),
    .B(_2393_),
    .C(_2394_),
    .Y(_2395_)
);

XNOR2X1 _13099_ (
    .A(_2395_),
    .B(_2392_),
    .Y(_2396_)
);

NAND2X1 _13100_ (
    .A(_2391_),
    .B(_2396_),
    .Y(_2397_)
);

INVX1 _13101_ (
    .A(_2392_),
    .Y(_2399_)
);

XNOR2X1 _13102_ (
    .A(_2395_),
    .B(_2399_),
    .Y(_2400_)
);

NAND2X1 _13103_ (
    .A(_2390_),
    .B(_2400_),
    .Y(_2401_)
);

NAND3X1 _13104_ (
    .A(_2386_),
    .B(_2397_),
    .C(_2401_),
    .Y(_2402_)
);

NAND2X1 _13105_ (
    .A(_2383_),
    .B(_2385_),
    .Y(_2403_)
);

NAND2X1 _13106_ (
    .A(_2391_),
    .B(_2400_),
    .Y(_2404_)
);

NAND2X1 _13107_ (
    .A(_2390_),
    .B(_2396_),
    .Y(_2405_)
);

NAND3X1 _13108_ (
    .A(_2403_),
    .B(_2404_),
    .C(_2405_),
    .Y(_2406_)
);

NOR2X1 _13109_ (
    .A(_1990_),
    .B(_1968_),
    .Y(_2407_)
);

OAI21X1 _13110_ (
    .A(_2407_),
    .B(_2088_),
    .C(_2001_),
    .Y(_2408_)
);

NAND3X1 _13111_ (
    .A(_2402_),
    .B(_2406_),
    .C(_2408_),
    .Y(_2409_)
);

AOI21X1 _13112_ (
    .A(_2405_),
    .B(_2404_),
    .C(_2403_),
    .Y(_2410_)
);

AOI21X1 _13113_ (
    .A(_2397_),
    .B(_2401_),
    .C(_2386_),
    .Y(_2411_)
);

AND2X2 _13114_ (
    .A(_1968_),
    .B(_1990_),
    .Y(_2412_)
);

AOI21X1 _13115_ (
    .A(_1914_),
    .B(_2066_),
    .C(_2412_),
    .Y(_2413_)
);

OAI21X1 _13116_ (
    .A(_2410_),
    .B(_2411_),
    .C(_2413_),
    .Y(_2414_)
);

NAND3X1 _13117_ (
    .A(_2378_),
    .B(_2414_),
    .C(_2409_),
    .Y(_2415_)
);

OAI21X1 _13118_ (
    .A(_1554_),
    .B(_1663_),
    .C(_1685_),
    .Y(_2416_)
);

NAND3X1 _13119_ (
    .A(_2402_),
    .B(_2406_),
    .C(_2413_),
    .Y(_2417_)
);

OAI21X1 _13120_ (
    .A(_2410_),
    .B(_2411_),
    .C(_2408_),
    .Y(_2418_)
);

NAND3X1 _13121_ (
    .A(_2416_),
    .B(_2418_),
    .C(_2417_),
    .Y(_2421_)
);

NAND2X1 _13122_ (
    .A(_2415_),
    .B(_2421_),
    .Y(_2422_)
);

OAI21X1 _13123_ (
    .A(_2305_),
    .B(_2131_),
    .C(_2315_),
    .Y(_2423_)
);

NOR2X1 _13124_ (
    .A(_177_),
    .B(_2012_),
    .Y(_2424_)
);

OR2X2 _13125_ (
    .A(_2034_),
    .B(_2424_),
    .Y(_2425_)
);

NOR2X1 _13126_ (
    .A(_4434__bF$buf3),
    .B(_5420__bF$buf2),
    .Y(_2426_)
);

NAND2X1 _13127_ (
    .A(breg_7_bF$buf1),
    .B(areg_9_bF$buf3),
    .Y(_2427_)
);

OAI21X1 _13128_ (
    .A(_5453__bF$buf0),
    .B(_6582__bF$buf1),
    .C(_1936_),
    .Y(_2428_)
);

OAI21X1 _13129_ (
    .A(_2012_),
    .B(_2427_),
    .C(_2428_),
    .Y(_2429_)
);

XNOR2X1 _13130_ (
    .A(_2429_),
    .B(_2426_),
    .Y(_2430_)
);

NAND2X1 _13131_ (
    .A(breg_4_bF$buf5),
    .B(areg_11_bF$buf4),
    .Y(_2432_)
);

OAI22X1 _13132_ (
    .A(_429_),
    .B(_2432_),
    .C(_2163_),
    .D(_2196_),
    .Y(_2433_)
);

NAND2X1 _13133_ (
    .A(_2433_),
    .B(_2430_),
    .Y(_2434_)
);

NAND2X1 _13134_ (
    .A(breg_6_bF$buf0),
    .B(areg_9_bF$buf2),
    .Y(_2435_)
);

XOR2X1 _13135_ (
    .A(_1936_),
    .B(_2435_),
    .Y(_2436_)
);

AND2X2 _13136_ (
    .A(_2436_),
    .B(_2426_),
    .Y(_2437_)
);

NOR2X1 _13137_ (
    .A(_2426_),
    .B(_2436_),
    .Y(_2438_)
);

INVX1 _13138_ (
    .A(_2433_),
    .Y(_2439_)
);

OAI21X1 _13139_ (
    .A(_2437_),
    .B(_2438_),
    .C(_2439_),
    .Y(_2440_)
);

NAND3X1 _13140_ (
    .A(_2440_),
    .B(_2425_),
    .C(_2434_),
    .Y(_2441_)
);

NOR2X1 _13141_ (
    .A(_2424_),
    .B(_2034_),
    .Y(_2443_)
);

NAND2X1 _13142_ (
    .A(_2439_),
    .B(_2430_),
    .Y(_2444_)
);

OAI21X1 _13143_ (
    .A(_2437_),
    .B(_2438_),
    .C(_2433_),
    .Y(_2445_)
);

NAND3X1 _13144_ (
    .A(_2443_),
    .B(_2445_),
    .C(_2444_),
    .Y(_2446_)
);

NAND2X1 _13145_ (
    .A(_2441_),
    .B(_2446_),
    .Y(_2447_)
);

OAI21X1 _13146_ (
    .A(_2300_),
    .B(_2303_),
    .C(_2293_),
    .Y(_2448_)
);

NOR2X1 _13147_ (
    .A(_4258__bF$buf3),
    .B(_7711__bF$buf1),
    .Y(_2449_)
);

INVX2 _13148_ (
    .A(_2449_),
    .Y(_2450_)
);

NAND2X1 _13149_ (
    .A(breg_3_bF$buf0),
    .B(areg_12_bF$buf4),
    .Y(_2451_)
);

NOR2X1 _13150_ (
    .A(_2432_),
    .B(_2451_),
    .Y(_2452_)
);

AND2X2 _13151_ (
    .A(_2432_),
    .B(_2451_),
    .Y(_2454_)
);

NOR2X1 _13152_ (
    .A(_2452_),
    .B(_2454_),
    .Y(_2455_)
);

XNOR2X1 _13153_ (
    .A(_2455_),
    .B(_2450_),
    .Y(_2456_)
);

AOI21X1 _13154_ (
    .A(_2270_),
    .B(_2288_),
    .C(_2290_),
    .Y(_2457_)
);

INVX2 _13155_ (
    .A(_2457_),
    .Y(_2458_)
);

NAND2X1 _13156_ (
    .A(breg_2_bF$buf3),
    .B(areg_13_bF$buf1),
    .Y(_2459_)
);

INVX2 _13157_ (
    .A(_2459_),
    .Y(_2460_)
);

NAND2X1 _13158_ (
    .A(breg_0_bF$buf4),
    .B(areg_15_bF$buf4),
    .Y(_2461_)
);

NOR2X1 _13159_ (
    .A(_2294_),
    .B(_2461_),
    .Y(_2462_)
);

INVX1 _13160_ (
    .A(_2462_),
    .Y(_2463_)
);

INVX8 _13161_ (
    .A(areg_15_bF$buf3),
    .Y(_2465_)
);

OAI21X1 _13162_ (
    .A(_2551__bF$buf0),
    .B(_2465__bF$buf4),
    .C(_2294_),
    .Y(_2466_)
);

NAND3X1 _13163_ (
    .A(_2460_),
    .B(_2466_),
    .C(_2463_),
    .Y(_2467_)
);

AND2X2 _13164_ (
    .A(_2294_),
    .B(_2461_),
    .Y(_2468_)
);

OAI21X1 _13165_ (
    .A(_2468_),
    .B(_2462_),
    .C(_2459_),
    .Y(_2469_)
);

NAND3X1 _13166_ (
    .A(_2469_),
    .B(_2467_),
    .C(_2458_),
    .Y(_2470_)
);

NOR3X1 _13167_ (
    .A(_2459_),
    .B(_2462_),
    .C(_2468_),
    .Y(_2471_)
);

AOI21X1 _13168_ (
    .A(_2466_),
    .B(_2463_),
    .C(_2460_),
    .Y(_2472_)
);

OAI21X1 _13169_ (
    .A(_2472_),
    .B(_2471_),
    .C(_2457_),
    .Y(_2473_)
);

NAND3X1 _13170_ (
    .A(_2456_),
    .B(_2470_),
    .C(_2473_),
    .Y(_2474_)
);

XNOR2X1 _13171_ (
    .A(_2455_),
    .B(_2449_),
    .Y(_2476_)
);

NOR3X1 _13172_ (
    .A(_2471_),
    .B(_2457_),
    .C(_2472_),
    .Y(_2477_)
);

AOI21X1 _13173_ (
    .A(_2469_),
    .B(_2467_),
    .C(_2458_),
    .Y(_2478_)
);

OAI21X1 _13174_ (
    .A(_2477_),
    .B(_2478_),
    .C(_2476_),
    .Y(_2479_)
);

AOI21X1 _13175_ (
    .A(_2474_),
    .B(_2479_),
    .C(_2448_),
    .Y(_2480_)
);

AOI21X1 _13176_ (
    .A(_2217_),
    .B(_2298_),
    .C(_2302_),
    .Y(_2481_)
);

OAI21X1 _13177_ (
    .A(_2472_),
    .B(_2471_),
    .C(_2458_),
    .Y(_2482_)
);

NAND3X1 _13178_ (
    .A(_2457_),
    .B(_2469_),
    .C(_2467_),
    .Y(_2483_)
);

AOI21X1 _13179_ (
    .A(_2483_),
    .B(_2482_),
    .C(_2476_),
    .Y(_2484_)
);

AOI21X1 _13180_ (
    .A(_2470_),
    .B(_2473_),
    .C(_2456_),
    .Y(_2485_)
);

NOR3X1 _13181_ (
    .A(_2484_),
    .B(_2485_),
    .C(_2481_),
    .Y(_2487_)
);

OAI21X1 _13182_ (
    .A(_2487_),
    .B(_2480_),
    .C(_2447_),
    .Y(_2488_)
);

AOI21X1 _13183_ (
    .A(_2445_),
    .B(_2444_),
    .C(_2443_),
    .Y(_2489_)
);

AOI21X1 _13184_ (
    .A(_2440_),
    .B(_2434_),
    .C(_2425_),
    .Y(_2490_)
);

NOR2X1 _13185_ (
    .A(_2489_),
    .B(_2490_),
    .Y(_2491_)
);

OAI21X1 _13186_ (
    .A(_2484_),
    .B(_2485_),
    .C(_2481_),
    .Y(_2492_)
);

NAND3X1 _13187_ (
    .A(_2448_),
    .B(_2474_),
    .C(_2479_),
    .Y(_2493_)
);

NAND3X1 _13188_ (
    .A(_2492_),
    .B(_2493_),
    .C(_2491_),
    .Y(_2494_)
);

NAND3X1 _13189_ (
    .A(_2423_),
    .B(_2488_),
    .C(_2494_),
    .Y(_2495_)
);

AOI21X1 _13190_ (
    .A(_2314_),
    .B(_2313_),
    .C(_2311_),
    .Y(_2496_)
);

AOI21X1 _13191_ (
    .A(_2492_),
    .B(_2493_),
    .C(_2491_),
    .Y(_2498_)
);

NOR3X1 _13192_ (
    .A(_2447_),
    .B(_2480_),
    .C(_2487_),
    .Y(_2499_)
);

OAI21X1 _13193_ (
    .A(_2499_),
    .B(_2498_),
    .C(_2496_),
    .Y(_2500_)
);

NAND3X1 _13194_ (
    .A(_2422_),
    .B(_2495_),
    .C(_2500_),
    .Y(_2501_)
);

AND2X2 _13195_ (
    .A(_2415_),
    .B(_2421_),
    .Y(_2502_)
);

OAI21X1 _13196_ (
    .A(_2499_),
    .B(_2498_),
    .C(_2423_),
    .Y(_2503_)
);

NAND3X1 _13197_ (
    .A(_2494_),
    .B(_2488_),
    .C(_2496_),
    .Y(_2504_)
);

NAND3X1 _13198_ (
    .A(_2503_),
    .B(_2504_),
    .C(_2502_),
    .Y(_2505_)
);

NAND3X1 _13199_ (
    .A(_2501_),
    .B(_2505_),
    .C(_2377_),
    .Y(_2506_)
);

NOR3X1 _13200_ (
    .A(_2318_),
    .B(_2319_),
    .C(_2320_),
    .Y(_2507_)
);

AOI21X1 _13201_ (
    .A(_1881_),
    .B(_2321_),
    .C(_2507_),
    .Y(_2509_)
);

AOI21X1 _13202_ (
    .A(_2504_),
    .B(_2503_),
    .C(_2502_),
    .Y(_2510_)
);

AOI21X1 _13203_ (
    .A(_2495_),
    .B(_2500_),
    .C(_2422_),
    .Y(_2511_)
);

OAI21X1 _13204_ (
    .A(_2510_),
    .B(_2511_),
    .C(_2509_),
    .Y(_2512_)
);

NAND3X1 _13205_ (
    .A(_2374_),
    .B(_2506_),
    .C(_2512_),
    .Y(_2513_)
);

OAI21X1 _13206_ (
    .A(_2510_),
    .B(_2511_),
    .C(_2377_),
    .Y(_2514_)
);

NAND3X1 _13207_ (
    .A(_2501_),
    .B(_2505_),
    .C(_2509_),
    .Y(_2515_)
);

NAND3X1 _13208_ (
    .A(_2373_),
    .B(_2514_),
    .C(_2515_),
    .Y(_2516_)
);

NAND3X1 _13209_ (
    .A(_2516_),
    .B(_2361_),
    .C(_2513_),
    .Y(_2517_)
);

AOI21X1 _13210_ (
    .A(_1467_),
    .B(_2331_),
    .C(_2333_),
    .Y(_2518_)
);

AOI21X1 _13211_ (
    .A(_2514_),
    .B(_2515_),
    .C(_2373_),
    .Y(_2520_)
);

AOI21X1 _13212_ (
    .A(_2506_),
    .B(_2512_),
    .C(_2374_),
    .Y(_2521_)
);

OAI21X1 _13213_ (
    .A(_2520_),
    .B(_2521_),
    .C(_2518_),
    .Y(_2522_)
);

NAND3X1 _13214_ (
    .A(_2360_),
    .B(_2517_),
    .C(_2522_),
    .Y(_2523_)
);

OAI21X1 _13215_ (
    .A(_2520_),
    .B(_2521_),
    .C(_2361_),
    .Y(_2524_)
);

NAND3X1 _13216_ (
    .A(_2513_),
    .B(_2516_),
    .C(_2518_),
    .Y(_2525_)
);

NAND3X1 _13217_ (
    .A(_2359_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_)
);

NAND3X1 _13218_ (
    .A(_2358_),
    .B(_2523_),
    .C(_2526_),
    .Y(_2527_)
);

NAND3X1 _13219_ (
    .A(_2359_),
    .B(_2517_),
    .C(_2522_),
    .Y(_2528_)
);

NAND3X1 _13220_ (
    .A(_2360_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2529_)
);

NAND3X1 _13221_ (
    .A(_2336_),
    .B(_2528_),
    .C(_2529_),
    .Y(_2531_)
);

NAND2X1 _13222_ (
    .A(_2527_),
    .B(_2531_),
    .Y(_2532_)
);

OAI21X1 _13223_ (
    .A(_2351_),
    .B(_2346_),
    .C(_2341_),
    .Y(_2533_)
);

OR2X2 _13224_ (
    .A(_2533_),
    .B(_2532_),
    .Y(_2534_)
);

NAND2X1 _13225_ (
    .A(_2532_),
    .B(_2533_),
    .Y(_2535_)
);

NAND2X1 _13226_ (
    .A(_2535_),
    .B(_2534_),
    .Y(_2536_)
);

XNOR2X1 _13227_ (
    .A(_2356_),
    .B(_2536_),
    .Y(_0_[15])
);

AOI22X1 _13228_ (
    .A(_2349_),
    .B(_2352_),
    .C(_2534_),
    .D(_2535_),
    .Y(_2537_)
);

NOR2X1 _13229_ (
    .A(_2346_),
    .B(_2345_),
    .Y(_2538_)
);

INVX1 _13230_ (
    .A(_2538_),
    .Y(_2539_)
);

NOR2X1 _13231_ (
    .A(_2532_),
    .B(_2533_),
    .Y(_2541_)
);

AND2X2 _13232_ (
    .A(_2533_),
    .B(_2532_),
    .Y(_2542_)
);

OAI21X1 _13233_ (
    .A(_2542_),
    .B(_2541_),
    .C(_2355_),
    .Y(_2543_)
);

OAI21X1 _13234_ (
    .A(_2539_),
    .B(_2532_),
    .C(_2543_),
    .Y(_2544_)
);

AOI21X1 _13235_ (
    .A(_2537_),
    .B(_1412_),
    .C(_2544_),
    .Y(_2545_)
);

NAND3X1 _13236_ (
    .A(_2336_),
    .B(_2523_),
    .C(_2526_),
    .Y(_2546_)
);

NAND3X1 _13237_ (
    .A(_2358_),
    .B(_2528_),
    .C(_2529_),
    .Y(_2547_)
);

AOI21X1 _13238_ (
    .A(_2546_),
    .B(_2547_),
    .C(_2341_),
    .Y(_2548_)
);

AOI21X1 _13239_ (
    .A(_2528_),
    .B(_2529_),
    .C(_2336_),
    .Y(_2549_)
);

AOI21X1 _13240_ (
    .A(_2516_),
    .B(_2513_),
    .C(_2361_),
    .Y(_2550_)
);

OAI21X1 _13241_ (
    .A(_2550_),
    .B(_2359_),
    .C(_2517_),
    .Y(_2552_)
);

NAND2X1 _13242_ (
    .A(_2370_),
    .B(_2372_),
    .Y(_2553_)
);

INVX2 _13243_ (
    .A(_2553_),
    .Y(_2554_)
);

AOI21X1 _13244_ (
    .A(_2501_),
    .B(_2505_),
    .C(_2377_),
    .Y(_2555_)
);

OAI21X1 _13245_ (
    .A(_2555_),
    .B(_2373_),
    .C(_2506_),
    .Y(_2556_)
);

INVX1 _13246_ (
    .A(_2363_),
    .Y(_2557_)
);

NAND2X1 _13247_ (
    .A(areg_1_bF$buf4),
    .B(breg_16_bF$buf5),
    .Y(_2558_)
);

OR2X2 _13248_ (
    .A(_2557_),
    .B(_2558_),
    .Y(_2559_)
);

INVX8 _13249_ (
    .A(breg_16_bF$buf4),
    .Y(_2560_)
);

NAND2X1 _13250_ (
    .A(areg_1_bF$buf3),
    .B(breg_15_bF$buf4),
    .Y(_2561_)
);

OAI21X1 _13251_ (
    .A(_2376__bF$buf0),
    .B(_2560__bF$buf4),
    .C(_2561_),
    .Y(_2563_)
);

AND2X2 _13252_ (
    .A(_2559_),
    .B(_2563_),
    .Y(_2564_)
);

OAI21X1 _13253_ (
    .A(_1511_),
    .B(_2381_),
    .C(_2385_),
    .Y(_2565_)
);

NAND2X1 _13254_ (
    .A(_2564_),
    .B(_2565_),
    .Y(_2566_)
);

INVX1 _13255_ (
    .A(_2566_),
    .Y(_2567_)
);

NOR2X1 _13256_ (
    .A(_2564_),
    .B(_2565_),
    .Y(_2568_)
);

OAI21X1 _13257_ (
    .A(_2567_),
    .B(_2568_),
    .C(_2368_),
    .Y(_2569_)
);

NOR2X1 _13258_ (
    .A(_2568_),
    .B(_2567_),
    .Y(_2570_)
);

NAND2X1 _13259_ (
    .A(_2369_),
    .B(_2570_),
    .Y(_2571_)
);

AND2X2 _13260_ (
    .A(_2571_),
    .B(_2569_),
    .Y(_2572_)
);

NAND2X1 _13261_ (
    .A(_2414_),
    .B(_2409_),
    .Y(_2574_)
);

OAI21X1 _13262_ (
    .A(_2574_),
    .B(_2378_),
    .C(_2409_),
    .Y(_2575_)
);

XNOR2X1 _13263_ (
    .A(_2575_),
    .B(_2572_),
    .Y(_2576_)
);

INVX2 _13264_ (
    .A(_2576_),
    .Y(_2577_)
);

AOI21X1 _13265_ (
    .A(_2488_),
    .B(_2494_),
    .C(_2423_),
    .Y(_2578_)
);

OAI21X1 _13266_ (
    .A(_2502_),
    .B(_2578_),
    .C(_2495_),
    .Y(_2579_)
);

AOI21X1 _13267_ (
    .A(_2391_),
    .B(_2396_),
    .C(_2410_),
    .Y(_2580_)
);

NOR2X1 _13268_ (
    .A(_2519__bF$buf3),
    .B(_2379_),
    .Y(_2581_)
);

INVX1 _13269_ (
    .A(_2581_),
    .Y(_2582_)
);

NAND2X1 _13270_ (
    .A(areg_4_bF$buf4),
    .B(breg_12_bF$buf0),
    .Y(_2583_)
);

NOR2X1 _13271_ (
    .A(_2381_),
    .B(_2583_),
    .Y(_2585_)
);

INVX8 _13272_ (
    .A(breg_12_bF$buf4),
    .Y(_2586_)
);

OAI21X1 _13273_ (
    .A(_2562__bF$buf1),
    .B(_2586__bF$buf4),
    .C(_2381_),
    .Y(_2587_)
);

INVX1 _13274_ (
    .A(_2587_),
    .Y(_2588_)
);

NOR2X1 _13275_ (
    .A(_2585_),
    .B(_2588_),
    .Y(_2589_)
);

XNOR2X1 _13276_ (
    .A(_2589_),
    .B(_2582_),
    .Y(_2590_)
);

NAND2X1 _13277_ (
    .A(areg_6_bF$buf0),
    .B(breg_9_bF$buf4),
    .Y(_2591_)
);

NOR2X1 _13278_ (
    .A(_1598_),
    .B(_2591_),
    .Y(_2592_)
);

AOI21X1 _13279_ (
    .A(_2392_),
    .B(_2394_),
    .C(_2592_),
    .Y(_2593_)
);

INVX2 _13280_ (
    .A(_2593_),
    .Y(_2594_)
);

NOR2X1 _13281_ (
    .A(_2825__bF$buf2),
    .B(_8555_),
    .Y(_2595_)
);

NAND2X1 _13282_ (
    .A(areg_7_bF$buf2),
    .B(breg_10_bF$buf2),
    .Y(_2596_)
);

OAI21X1 _13283_ (
    .A(_4434__bF$buf2),
    .B(_6044__bF$buf0),
    .C(_2393_),
    .Y(_2597_)
);

OAI21X1 _13284_ (
    .A(_2591_),
    .B(_2596_),
    .C(_2597_),
    .Y(_2598_)
);

XNOR2X1 _13285_ (
    .A(_2598_),
    .B(_2595_),
    .Y(_2599_)
);

NAND2X1 _13286_ (
    .A(_2594_),
    .B(_2599_),
    .Y(_2600_)
);

INVX1 _13287_ (
    .A(_2595_),
    .Y(_2601_)
);

XNOR2X1 _13288_ (
    .A(_2598_),
    .B(_2601_),
    .Y(_2602_)
);

NAND2X1 _13289_ (
    .A(_2593_),
    .B(_2602_),
    .Y(_2603_)
);

NAND3X1 _13290_ (
    .A(_2590_),
    .B(_2600_),
    .C(_2603_),
    .Y(_2604_)
);

XNOR2X1 _13291_ (
    .A(_2589_),
    .B(_2581_),
    .Y(_2606_)
);

NAND2X1 _13292_ (
    .A(_2594_),
    .B(_2602_),
    .Y(_2607_)
);

NAND2X1 _13293_ (
    .A(_2593_),
    .B(_2599_),
    .Y(_2608_)
);

NAND3X1 _13294_ (
    .A(_2606_),
    .B(_2607_),
    .C(_2608_),
    .Y(_2609_)
);

NOR2X1 _13295_ (
    .A(_2433_),
    .B(_2430_),
    .Y(_2610_)
);

OAI21X1 _13296_ (
    .A(_2610_),
    .B(_2443_),
    .C(_2434_),
    .Y(_2611_)
);

NAND3X1 _13297_ (
    .A(_2604_),
    .B(_2609_),
    .C(_2611_),
    .Y(_2612_)
);

AOI21X1 _13298_ (
    .A(_2608_),
    .B(_2607_),
    .C(_2606_),
    .Y(_2613_)
);

AOI21X1 _13299_ (
    .A(_2600_),
    .B(_2603_),
    .C(_2590_),
    .Y(_2614_)
);

AND2X2 _13300_ (
    .A(_2430_),
    .B(_2433_),
    .Y(_2615_)
);

AOI21X1 _13301_ (
    .A(_2425_),
    .B(_2440_),
    .C(_2615_),
    .Y(_2618_)
);

OAI21X1 _13302_ (
    .A(_2613_),
    .B(_2614_),
    .C(_2618_),
    .Y(_2619_)
);

NAND3X1 _13303_ (
    .A(_2580_),
    .B(_2619_),
    .C(_2612_),
    .Y(_2620_)
);

OAI21X1 _13304_ (
    .A(_2390_),
    .B(_2400_),
    .C(_2402_),
    .Y(_2621_)
);

NOR3X1 _13305_ (
    .A(_2613_),
    .B(_2614_),
    .C(_2618_),
    .Y(_2622_)
);

AOI21X1 _13306_ (
    .A(_2604_),
    .B(_2609_),
    .C(_2611_),
    .Y(_2623_)
);

OAI21X1 _13307_ (
    .A(_2622_),
    .B(_2623_),
    .C(_2621_),
    .Y(_2624_)
);

NAND2X1 _13308_ (
    .A(_2620_),
    .B(_2624_),
    .Y(_2625_)
);

OAI21X1 _13309_ (
    .A(_2480_),
    .B(_2447_),
    .C(_2493_),
    .Y(_2626_)
);

NOR2X1 _13310_ (
    .A(_1936_),
    .B(_2435_),
    .Y(_2627_)
);

OR2X2 _13311_ (
    .A(_2437_),
    .B(_2627_),
    .Y(_2629_)
);

NOR2X1 _13312_ (
    .A(_5190__bF$buf0),
    .B(_5420__bF$buf1),
    .Y(_2630_)
);

NAND2X1 _13313_ (
    .A(breg_7_bF$buf0),
    .B(areg_10_bF$buf3),
    .Y(_2631_)
);

OAI21X1 _13314_ (
    .A(_5453__bF$buf5),
    .B(_7711__bF$buf0),
    .C(_2427_),
    .Y(_2632_)
);

OAI21X1 _13315_ (
    .A(_2435_),
    .B(_2631_),
    .C(_2632_),
    .Y(_2633_)
);

XNOR2X1 _13316_ (
    .A(_2633_),
    .B(_2630_),
    .Y(_2634_)
);

NAND2X1 _13317_ (
    .A(breg_4_bF$buf4),
    .B(areg_12_bF$buf3),
    .Y(_2635_)
);

OAI22X1 _13318_ (
    .A(_2174_),
    .B(_2635_),
    .C(_2450_),
    .D(_2454_),
    .Y(_2636_)
);

NAND2X1 _13319_ (
    .A(_2636_),
    .B(_2634_),
    .Y(_2637_)
);

NAND2X1 _13320_ (
    .A(breg_6_bF$buf5),
    .B(areg_10_bF$buf2),
    .Y(_2638_)
);

XOR2X1 _13321_ (
    .A(_2427_),
    .B(_2638_),
    .Y(_2640_)
);

AND2X2 _13322_ (
    .A(_2640_),
    .B(_2630_),
    .Y(_2641_)
);

NOR2X1 _13323_ (
    .A(_2630_),
    .B(_2640_),
    .Y(_2642_)
);

INVX1 _13324_ (
    .A(_2636_),
    .Y(_2643_)
);

OAI21X1 _13325_ (
    .A(_2641_),
    .B(_2642_),
    .C(_2643_),
    .Y(_2644_)
);

NAND3X1 _13326_ (
    .A(_2644_),
    .B(_2629_),
    .C(_2637_),
    .Y(_2645_)
);

NOR2X1 _13327_ (
    .A(_2627_),
    .B(_2437_),
    .Y(_2646_)
);

NAND2X1 _13328_ (
    .A(_2643_),
    .B(_2634_),
    .Y(_2647_)
);

OAI21X1 _13329_ (
    .A(_2641_),
    .B(_2642_),
    .C(_2636_),
    .Y(_2648_)
);

NAND3X1 _13330_ (
    .A(_2646_),
    .B(_2648_),
    .C(_2647_),
    .Y(_2649_)
);

NAND2X1 _13331_ (
    .A(_2645_),
    .B(_2649_),
    .Y(_2651_)
);

OAI21X1 _13332_ (
    .A(_2478_),
    .B(_2476_),
    .C(_2470_),
    .Y(_2652_)
);

NOR2X1 _13333_ (
    .A(_4258__bF$buf2),
    .B(_9104__bF$buf0),
    .Y(_2653_)
);

INVX1 _13334_ (
    .A(_2653_),
    .Y(_2654_)
);

NAND2X1 _13335_ (
    .A(breg_3_bF$buf5),
    .B(areg_13_bF$buf0),
    .Y(_2655_)
);

NOR2X1 _13336_ (
    .A(_2635_),
    .B(_2655_),
    .Y(_2656_)
);

AND2X2 _13337_ (
    .A(_2635_),
    .B(_2655_),
    .Y(_2657_)
);

NOR2X1 _13338_ (
    .A(_2656_),
    .B(_2657_),
    .Y(_2658_)
);

XNOR2X1 _13339_ (
    .A(_2658_),
    .B(_2654_),
    .Y(_2659_)
);

AOI21X1 _13340_ (
    .A(_2460_),
    .B(_2466_),
    .C(_2462_),
    .Y(_2660_)
);

INVX2 _13341_ (
    .A(_2660_),
    .Y(_2662_)
);

NAND2X1 _13342_ (
    .A(breg_2_bF$buf2),
    .B(areg_14_bF$buf1),
    .Y(_2663_)
);

INVX2 _13343_ (
    .A(_2663_),
    .Y(_2664_)
);

NAND2X1 _13344_ (
    .A(breg_1_bF$buf4),
    .B(areg_15_bF$buf2),
    .Y(_2665_)
);

NAND2X1 _13345_ (
    .A(breg_0_bF$buf3),
    .B(areg_16_bF$buf5),
    .Y(_2666_)
);

NOR2X1 _13346_ (
    .A(_2665_),
    .B(_2666_),
    .Y(_2667_)
);

INVX1 _13347_ (
    .A(_2667_),
    .Y(_2668_)
);

INVX8 _13348_ (
    .A(areg_16_bF$buf4),
    .Y(_2669_)
);

OAI21X1 _13349_ (
    .A(_2551__bF$buf3),
    .B(_2669__bF$buf3),
    .C(_2665_),
    .Y(_2670_)
);

NAND3X1 _13350_ (
    .A(_2664_),
    .B(_2670_),
    .C(_2668_),
    .Y(_2671_)
);

AND2X2 _13351_ (
    .A(_2665_),
    .B(_2666_),
    .Y(_2673_)
);

OAI21X1 _13352_ (
    .A(_2673_),
    .B(_2667_),
    .C(_2663_),
    .Y(_2674_)
);

NAND3X1 _13353_ (
    .A(_2674_),
    .B(_2671_),
    .C(_2662_),
    .Y(_2675_)
);

NOR3X1 _13354_ (
    .A(_2663_),
    .B(_2667_),
    .C(_2673_),
    .Y(_2676_)
);

AOI21X1 _13355_ (
    .A(_2670_),
    .B(_2668_),
    .C(_2664_),
    .Y(_2677_)
);

OAI21X1 _13356_ (
    .A(_2677_),
    .B(_2676_),
    .C(_2660_),
    .Y(_2678_)
);

NAND3X1 _13357_ (
    .A(_2675_),
    .B(_2659_),
    .C(_2678_),
    .Y(_2679_)
);

XNOR2X1 _13358_ (
    .A(_2658_),
    .B(_2653_),
    .Y(_2680_)
);

NOR3X1 _13359_ (
    .A(_2676_),
    .B(_2660_),
    .C(_2677_),
    .Y(_2681_)
);

AOI21X1 _13360_ (
    .A(_2674_),
    .B(_2671_),
    .C(_2662_),
    .Y(_2682_)
);

OAI21X1 _13361_ (
    .A(_2681_),
    .B(_2682_),
    .C(_2680_),
    .Y(_2684_)
);

AOI21X1 _13362_ (
    .A(_2679_),
    .B(_2684_),
    .C(_2652_),
    .Y(_2685_)
);

AOI21X1 _13363_ (
    .A(_2456_),
    .B(_2473_),
    .C(_2477_),
    .Y(_2686_)
);

OAI21X1 _13364_ (
    .A(_2677_),
    .B(_2676_),
    .C(_2662_),
    .Y(_2687_)
);

NAND3X1 _13365_ (
    .A(_2660_),
    .B(_2674_),
    .C(_2671_),
    .Y(_2688_)
);

AOI21X1 _13366_ (
    .A(_2688_),
    .B(_2687_),
    .C(_2680_),
    .Y(_2689_)
);

AOI21X1 _13367_ (
    .A(_2675_),
    .B(_2678_),
    .C(_2659_),
    .Y(_2690_)
);

NOR3X1 _13368_ (
    .A(_2689_),
    .B(_2690_),
    .C(_2686_),
    .Y(_2691_)
);

OAI21X1 _13369_ (
    .A(_2691_),
    .B(_2685_),
    .C(_2651_),
    .Y(_2692_)
);

AND2X2 _13370_ (
    .A(_2645_),
    .B(_2649_),
    .Y(_2693_)
);

OAI21X1 _13371_ (
    .A(_2689_),
    .B(_2690_),
    .C(_2686_),
    .Y(_2695_)
);

NAND3X1 _13372_ (
    .A(_2652_),
    .B(_2679_),
    .C(_2684_),
    .Y(_2696_)
);

NAND3X1 _13373_ (
    .A(_2696_),
    .B(_2695_),
    .C(_2693_),
    .Y(_2697_)
);

NAND3X1 _13374_ (
    .A(_2626_),
    .B(_2692_),
    .C(_2697_),
    .Y(_2698_)
);

AOI21X1 _13375_ (
    .A(_2492_),
    .B(_2491_),
    .C(_2487_),
    .Y(_2699_)
);

AOI21X1 _13376_ (
    .A(_2696_),
    .B(_2695_),
    .C(_2693_),
    .Y(_2700_)
);

NOR3X1 _13377_ (
    .A(_2651_),
    .B(_2685_),
    .C(_2691_),
    .Y(_2701_)
);

OAI21X1 _13378_ (
    .A(_2701_),
    .B(_2700_),
    .C(_2699_),
    .Y(_2702_)
);

NAND3X1 _13379_ (
    .A(_2698_),
    .B(_2702_),
    .C(_2625_),
    .Y(_2703_)
);

NAND3X1 _13380_ (
    .A(_2621_),
    .B(_2619_),
    .C(_2612_),
    .Y(_2704_)
);

OAI21X1 _13381_ (
    .A(_2622_),
    .B(_2623_),
    .C(_2580_),
    .Y(_2706_)
);

NAND2X1 _13382_ (
    .A(_2704_),
    .B(_2706_),
    .Y(_2707_)
);

OAI21X1 _13383_ (
    .A(_2701_),
    .B(_2700_),
    .C(_2626_),
    .Y(_2708_)
);

NAND3X1 _13384_ (
    .A(_2692_),
    .B(_2697_),
    .C(_2699_),
    .Y(_2709_)
);

NAND3X1 _13385_ (
    .A(_2709_),
    .B(_2708_),
    .C(_2707_),
    .Y(_2710_)
);

NAND3X1 _13386_ (
    .A(_2703_),
    .B(_2710_),
    .C(_2579_),
    .Y(_2711_)
);

NOR3X1 _13387_ (
    .A(_2499_),
    .B(_2498_),
    .C(_2496_),
    .Y(_2712_)
);

AOI21X1 _13388_ (
    .A(_2422_),
    .B(_2500_),
    .C(_2712_),
    .Y(_2713_)
);

AOI21X1 _13389_ (
    .A(_2709_),
    .B(_2708_),
    .C(_2707_),
    .Y(_2714_)
);

AOI21X1 _13390_ (
    .A(_2698_),
    .B(_2702_),
    .C(_2625_),
    .Y(_2715_)
);

OAI21X1 _13391_ (
    .A(_2714_),
    .B(_2715_),
    .C(_2713_),
    .Y(_2717_)
);

NAND3X1 _13392_ (
    .A(_2711_),
    .B(_2577_),
    .C(_2717_),
    .Y(_2718_)
);

OAI21X1 _13393_ (
    .A(_2714_),
    .B(_2715_),
    .C(_2579_),
    .Y(_2719_)
);

NAND3X1 _13394_ (
    .A(_2703_),
    .B(_2710_),
    .C(_2713_),
    .Y(_2720_)
);

NAND3X1 _13395_ (
    .A(_2576_),
    .B(_2719_),
    .C(_2720_),
    .Y(_2721_)
);

NAND3X1 _13396_ (
    .A(_2721_),
    .B(_2556_),
    .C(_2718_),
    .Y(_2722_)
);

NOR3X1 _13397_ (
    .A(_2510_),
    .B(_2511_),
    .C(_2509_),
    .Y(_2723_)
);

AOI21X1 _13398_ (
    .A(_2374_),
    .B(_2512_),
    .C(_2723_),
    .Y(_2724_)
);

AOI21X1 _13399_ (
    .A(_2719_),
    .B(_2720_),
    .C(_2576_),
    .Y(_2725_)
);

AOI21X1 _13400_ (
    .A(_2711_),
    .B(_2717_),
    .C(_2577_),
    .Y(_2726_)
);

OAI21X1 _13401_ (
    .A(_2725_),
    .B(_2726_),
    .C(_2724_),
    .Y(_2728_)
);

NAND3X1 _13402_ (
    .A(_2554_),
    .B(_2722_),
    .C(_2728_),
    .Y(_2729_)
);

OAI21X1 _13403_ (
    .A(_2725_),
    .B(_2726_),
    .C(_2556_),
    .Y(_2730_)
);

NAND3X1 _13404_ (
    .A(_2718_),
    .B(_2721_),
    .C(_2724_),
    .Y(_2731_)
);

NAND3X1 _13405_ (
    .A(_2553_),
    .B(_2730_),
    .C(_2731_),
    .Y(_2732_)
);

NAND3X1 _13406_ (
    .A(_2729_),
    .B(_2552_),
    .C(_2732_),
    .Y(_2733_)
);

NOR3X1 _13407_ (
    .A(_2520_),
    .B(_2521_),
    .C(_2518_),
    .Y(_2734_)
);

AOI21X1 _13408_ (
    .A(_2360_),
    .B(_2522_),
    .C(_2734_),
    .Y(_2735_)
);

AOI21X1 _13409_ (
    .A(_2730_),
    .B(_2731_),
    .C(_2553_),
    .Y(_2736_)
);

AOI21X1 _13410_ (
    .A(_2722_),
    .B(_2728_),
    .C(_2554_),
    .Y(_2737_)
);

OAI21X1 _13411_ (
    .A(_2736_),
    .B(_2737_),
    .C(_2735_),
    .Y(_2739_)
);

NAND3X1 _13412_ (
    .A(_2733_),
    .B(_2549_),
    .C(_2739_),
    .Y(_2740_)
);

OAI21X1 _13413_ (
    .A(_2736_),
    .B(_2737_),
    .C(_2552_),
    .Y(_2741_)
);

NAND3X1 _13414_ (
    .A(_2729_),
    .B(_2732_),
    .C(_2735_),
    .Y(_2742_)
);

NAND3X1 _13415_ (
    .A(_2527_),
    .B(_2741_),
    .C(_2742_),
    .Y(_2743_)
);

NAND3X1 _13416_ (
    .A(_2548_),
    .B(_2740_),
    .C(_2743_),
    .Y(_2744_)
);

NAND3X1 _13417_ (
    .A(_2350_),
    .B(_2531_),
    .C(_2527_),
    .Y(_2745_)
);

NAND3X1 _13418_ (
    .A(_2527_),
    .B(_2733_),
    .C(_2739_),
    .Y(_2746_)
);

NAND3X1 _13419_ (
    .A(_2549_),
    .B(_2741_),
    .C(_2742_),
    .Y(_2747_)
);

NAND3X1 _13420_ (
    .A(_2745_),
    .B(_2746_),
    .C(_2747_),
    .Y(_2748_)
);

NAND2X1 _13421_ (
    .A(_2748_),
    .B(_2744_),
    .Y(_2750_)
);

XOR2X1 _13422_ (
    .A(_2545_),
    .B(_2750_),
    .Y(_0_[16])
);

OAI21X1 _13423_ (
    .A(_2545_),
    .B(_2750_),
    .C(_2744_),
    .Y(_2751_)
);

AOI21X1 _13424_ (
    .A(_2741_),
    .B(_2742_),
    .C(_2527_),
    .Y(_2752_)
);

NOR3X1 _13425_ (
    .A(_2736_),
    .B(_2737_),
    .C(_2735_),
    .Y(_2753_)
);

AOI21X1 _13426_ (
    .A(_2721_),
    .B(_2718_),
    .C(_2556_),
    .Y(_2754_)
);

OAI21X1 _13427_ (
    .A(_2754_),
    .B(_2553_),
    .C(_2722_),
    .Y(_2755_)
);

NAND2X1 _13428_ (
    .A(_2572_),
    .B(_2575_),
    .Y(_2756_)
);

INVX2 _13429_ (
    .A(_2756_),
    .Y(_2757_)
);

AOI21X1 _13430_ (
    .A(_2703_),
    .B(_2710_),
    .C(_2579_),
    .Y(_2758_)
);

OAI21X1 _13431_ (
    .A(_2758_),
    .B(_2576_),
    .C(_2711_),
    .Y(_2760_)
);

INVX1 _13432_ (
    .A(_2571_),
    .Y(_2761_)
);

OAI21X1 _13433_ (
    .A(_2623_),
    .B(_2580_),
    .C(_2612_),
    .Y(_2762_)
);

INVX4 _13434_ (
    .A(breg_17_bF$buf4),
    .Y(_2763_)
);

NOR2X1 _13435_ (
    .A(_2376__bF$buf3),
    .B(_2763_),
    .Y(_2764_)
);

NAND2X1 _13436_ (
    .A(areg_2_bF$buf2),
    .B(breg_15_bF$buf3),
    .Y(_2765_)
);

XOR2X1 _13437_ (
    .A(_2558_),
    .B(_2765_),
    .Y(_2766_)
);

NAND2X1 _13438_ (
    .A(_2764_),
    .B(_2766_),
    .Y(_2767_)
);

NAND2X1 _13439_ (
    .A(areg_2_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_2768_)
);

OAI21X1 _13440_ (
    .A(_2519__bF$buf2),
    .B(_2362__bF$buf4),
    .C(_2558_),
    .Y(_2769_)
);

OAI21X1 _13441_ (
    .A(_2561_),
    .B(_2768_),
    .C(_2769_),
    .Y(_2771_)
);

OAI21X1 _13442_ (
    .A(_2376__bF$buf2),
    .B(_2763_),
    .C(_2771_),
    .Y(_2772_)
);

AOI21X1 _13443_ (
    .A(_2581_),
    .B(_2587_),
    .C(_2585_),
    .Y(_2773_)
);

INVX1 _13444_ (
    .A(_2773_),
    .Y(_2774_)
);

NAND3X1 _13445_ (
    .A(_2772_),
    .B(_2774_),
    .C(_2767_),
    .Y(_2775_)
);

AOI21X1 _13446_ (
    .A(_2772_),
    .B(_2767_),
    .C(_2774_),
    .Y(_2776_)
);

INVX1 _13447_ (
    .A(_2776_),
    .Y(_2777_)
);

NAND2X1 _13448_ (
    .A(_2775_),
    .B(_2777_),
    .Y(_2778_)
);

OAI21X1 _13449_ (
    .A(_2557_),
    .B(_2558_),
    .C(_2566_),
    .Y(_2779_)
);

XNOR2X1 _13450_ (
    .A(_2779_),
    .B(_2778_),
    .Y(_2780_)
);

NAND2X1 _13451_ (
    .A(_2780_),
    .B(_2762_),
    .Y(_2782_)
);

AOI21X1 _13452_ (
    .A(_2621_),
    .B(_2619_),
    .C(_2622_),
    .Y(_2783_)
);

XOR2X1 _13453_ (
    .A(_2779_),
    .B(_2778_),
    .Y(_2784_)
);

NAND2X1 _13454_ (
    .A(_2784_),
    .B(_2783_),
    .Y(_2785_)
);

NAND3X1 _13455_ (
    .A(_2761_),
    .B(_2782_),
    .C(_2785_),
    .Y(_2786_)
);

NAND2X1 _13456_ (
    .A(_2780_),
    .B(_2783_),
    .Y(_2787_)
);

NAND2X1 _13457_ (
    .A(_2784_),
    .B(_2762_),
    .Y(_2788_)
);

NAND3X1 _13458_ (
    .A(_2571_),
    .B(_2788_),
    .C(_2787_),
    .Y(_2789_)
);

AND2X2 _13459_ (
    .A(_2786_),
    .B(_2789_),
    .Y(_2790_)
);

AOI21X1 _13460_ (
    .A(_2692_),
    .B(_2697_),
    .C(_2626_),
    .Y(_2791_)
);

OAI21X1 _13461_ (
    .A(_2707_),
    .B(_2791_),
    .C(_2698_),
    .Y(_2793_)
);

AOI21X1 _13462_ (
    .A(_2594_),
    .B(_2599_),
    .C(_2613_),
    .Y(_2794_)
);

NOR2X1 _13463_ (
    .A(_2792_),
    .B(_2379_),
    .Y(_2795_)
);

NAND2X1 _13464_ (
    .A(areg_5_bF$buf4),
    .B(breg_13_bF$buf0),
    .Y(_2796_)
);

NAND2X1 _13465_ (
    .A(areg_4_bF$buf3),
    .B(breg_13_bF$buf4),
    .Y(_2797_)
);

OAI21X1 _13466_ (
    .A(_2825__bF$buf1),
    .B(_2586__bF$buf3),
    .C(_2797_),
    .Y(_2798_)
);

OAI21X1 _13467_ (
    .A(_2583_),
    .B(_2796_),
    .C(_2798_),
    .Y(_2799_)
);

XNOR2X1 _13468_ (
    .A(_2799_),
    .B(_2795_),
    .Y(_2800_)
);

NAND2X1 _13469_ (
    .A(areg_7_bF$buf1),
    .B(breg_9_bF$buf3),
    .Y(_2801_)
);

NOR2X1 _13470_ (
    .A(_2393_),
    .B(_2801_),
    .Y(_2802_)
);

AOI21X1 _13471_ (
    .A(_2595_),
    .B(_2597_),
    .C(_2802_),
    .Y(_2804_)
);

INVX2 _13472_ (
    .A(_2804_),
    .Y(_2805_)
);

NOR2X1 _13473_ (
    .A(_3646__bF$buf1),
    .B(_8555_),
    .Y(_2806_)
);

NAND2X1 _13474_ (
    .A(areg_8_bF$buf1),
    .B(breg_10_bF$buf1),
    .Y(_2807_)
);

OAI21X1 _13475_ (
    .A(_5190__bF$buf3),
    .B(_6044__bF$buf5),
    .C(_2596_),
    .Y(_2808_)
);

OAI21X1 _13476_ (
    .A(_2801_),
    .B(_2807_),
    .C(_2808_),
    .Y(_2809_)
);

XNOR2X1 _13477_ (
    .A(_2809_),
    .B(_2806_),
    .Y(_2810_)
);

NAND2X1 _13478_ (
    .A(_2805_),
    .B(_2810_),
    .Y(_2811_)
);

INVX1 _13479_ (
    .A(_2806_),
    .Y(_2812_)
);

NOR2X1 _13480_ (
    .A(_2812_),
    .B(_2809_),
    .Y(_2813_)
);

NAND2X1 _13481_ (
    .A(areg_8_bF$buf0),
    .B(breg_9_bF$buf2),
    .Y(_2815_)
);

NOR2X1 _13482_ (
    .A(_2596_),
    .B(_2815_),
    .Y(_2816_)
);

INVX1 _13483_ (
    .A(_2816_),
    .Y(_2817_)
);

AOI21X1 _13484_ (
    .A(_2808_),
    .B(_2817_),
    .C(_2806_),
    .Y(_2818_)
);

OAI21X1 _13485_ (
    .A(_2813_),
    .B(_2818_),
    .C(_2804_),
    .Y(_2819_)
);

NAND3X1 _13486_ (
    .A(_2800_),
    .B(_2819_),
    .C(_2811_),
    .Y(_2820_)
);

INVX1 _13487_ (
    .A(_2800_),
    .Y(_2821_)
);

OAI21X1 _13488_ (
    .A(_2813_),
    .B(_2818_),
    .C(_2805_),
    .Y(_2822_)
);

NAND2X1 _13489_ (
    .A(_2804_),
    .B(_2810_),
    .Y(_2823_)
);

NAND3X1 _13490_ (
    .A(_2821_),
    .B(_2822_),
    .C(_2823_),
    .Y(_2824_)
);

NOR2X1 _13491_ (
    .A(_2636_),
    .B(_2634_),
    .Y(_2826_)
);

OAI21X1 _13492_ (
    .A(_2826_),
    .B(_2646_),
    .C(_2637_),
    .Y(_2827_)
);

NAND3X1 _13493_ (
    .A(_2820_),
    .B(_2824_),
    .C(_2827_),
    .Y(_2828_)
);

AOI21X1 _13494_ (
    .A(_2822_),
    .B(_2823_),
    .C(_2821_),
    .Y(_2829_)
);

AOI21X1 _13495_ (
    .A(_2819_),
    .B(_2811_),
    .C(_2800_),
    .Y(_2830_)
);

AND2X2 _13496_ (
    .A(_2634_),
    .B(_2636_),
    .Y(_2831_)
);

AOI21X1 _13497_ (
    .A(_2629_),
    .B(_2644_),
    .C(_2831_),
    .Y(_2832_)
);

OAI21X1 _13498_ (
    .A(_2829_),
    .B(_2830_),
    .C(_2832_),
    .Y(_2833_)
);

NAND3X1 _13499_ (
    .A(_2794_),
    .B(_2833_),
    .C(_2828_),
    .Y(_2834_)
);

OAI21X1 _13500_ (
    .A(_2593_),
    .B(_2602_),
    .C(_2604_),
    .Y(_2835_)
);

NOR3X1 _13501_ (
    .A(_2829_),
    .B(_2830_),
    .C(_2832_),
    .Y(_2837_)
);

AOI21X1 _13502_ (
    .A(_2820_),
    .B(_2824_),
    .C(_2827_),
    .Y(_2838_)
);

OAI21X1 _13503_ (
    .A(_2837_),
    .B(_2838_),
    .C(_2835_),
    .Y(_2839_)
);

NAND2X1 _13504_ (
    .A(_2834_),
    .B(_2839_),
    .Y(_2840_)
);

OAI21X1 _13505_ (
    .A(_2685_),
    .B(_2651_),
    .C(_2696_),
    .Y(_2841_)
);

NAND2X1 _13506_ (
    .A(_2630_),
    .B(_2640_),
    .Y(_2842_)
);

OAI21X1 _13507_ (
    .A(_2435_),
    .B(_2631_),
    .C(_2842_),
    .Y(_2843_)
);

NOR2X1 _13508_ (
    .A(_5420__bF$buf0),
    .B(_6582__bF$buf0),
    .Y(_2844_)
);

NAND2X1 _13509_ (
    .A(breg_6_bF$buf4),
    .B(areg_11_bF$buf3),
    .Y(_2845_)
);

XOR2X1 _13510_ (
    .A(_2631_),
    .B(_2845_),
    .Y(_2846_)
);

NAND2X1 _13511_ (
    .A(_2844_),
    .B(_2846_),
    .Y(_2848_)
);

NAND2X1 _13512_ (
    .A(breg_7_bF$buf5),
    .B(areg_11_bF$buf2),
    .Y(_2849_)
);

OAI21X1 _13513_ (
    .A(_5453__bF$buf4),
    .B(_9104__bF$buf3),
    .C(_2631_),
    .Y(_2850_)
);

OAI21X1 _13514_ (
    .A(_2638_),
    .B(_2849_),
    .C(_2850_),
    .Y(_2851_)
);

OAI21X1 _13515_ (
    .A(_5420__bF$buf3),
    .B(_6582__bF$buf3),
    .C(_2851_),
    .Y(_2852_)
);

OAI21X1 _13516_ (
    .A(_2365_),
    .B(_549__bF$buf3),
    .C(_2635_),
    .Y(_2853_)
);

AOI21X1 _13517_ (
    .A(_2653_),
    .B(_2853_),
    .C(_2656_),
    .Y(_2854_)
);

INVX2 _13518_ (
    .A(_2854_),
    .Y(_2855_)
);

NAND3X1 _13519_ (
    .A(_2852_),
    .B(_2855_),
    .C(_2848_),
    .Y(_2856_)
);

INVX1 _13520_ (
    .A(_2844_),
    .Y(_2857_)
);

NOR2X1 _13521_ (
    .A(_2857_),
    .B(_2851_),
    .Y(_2859_)
);

NOR2X1 _13522_ (
    .A(_2844_),
    .B(_2846_),
    .Y(_2860_)
);

OAI21X1 _13523_ (
    .A(_2860_),
    .B(_2859_),
    .C(_2854_),
    .Y(_2861_)
);

NAND3X1 _13524_ (
    .A(_2843_),
    .B(_2856_),
    .C(_2861_),
    .Y(_2862_)
);

NOR2X1 _13525_ (
    .A(_2427_),
    .B(_2638_),
    .Y(_2863_)
);

NOR2X1 _13526_ (
    .A(_2863_),
    .B(_2641_),
    .Y(_2864_)
);

NOR3X1 _13527_ (
    .A(_2859_),
    .B(_2854_),
    .C(_2860_),
    .Y(_2865_)
);

AOI21X1 _13528_ (
    .A(_2852_),
    .B(_2848_),
    .C(_2855_),
    .Y(_2866_)
);

OAI21X1 _13529_ (
    .A(_2865_),
    .B(_2866_),
    .C(_2864_),
    .Y(_2867_)
);

NAND2X1 _13530_ (
    .A(_2862_),
    .B(_2867_),
    .Y(_2868_)
);

OAI21X1 _13531_ (
    .A(_2682_),
    .B(_2680_),
    .C(_2675_),
    .Y(_2870_)
);

NAND2X1 _13532_ (
    .A(breg_5_bF$buf2),
    .B(areg_12_bF$buf2),
    .Y(_2871_)
);

NAND2X1 _13533_ (
    .A(breg_4_bF$buf3),
    .B(areg_13_bF$buf4),
    .Y(_2872_)
);

NAND2X1 _13534_ (
    .A(breg_3_bF$buf4),
    .B(areg_14_bF$buf0),
    .Y(_2873_)
);

XOR2X1 _13535_ (
    .A(_2872_),
    .B(_2873_),
    .Y(_2874_)
);

XNOR2X1 _13536_ (
    .A(_2874_),
    .B(_2871_),
    .Y(_2875_)
);

AOI21X1 _13537_ (
    .A(_2664_),
    .B(_2670_),
    .C(_2667_),
    .Y(_2876_)
);

INVX2 _13538_ (
    .A(_2876_),
    .Y(_2877_)
);

NAND2X1 _13539_ (
    .A(breg_2_bF$buf1),
    .B(areg_15_bF$buf1),
    .Y(_2878_)
);

INVX2 _13540_ (
    .A(_2878_),
    .Y(_2879_)
);

NAND2X1 _13541_ (
    .A(breg_1_bF$buf3),
    .B(areg_16_bF$buf3),
    .Y(_2881_)
);

NAND2X1 _13542_ (
    .A(breg_0_bF$buf2),
    .B(areg_17_bF$buf5),
    .Y(_2882_)
);

OR2X2 _13543_ (
    .A(_2881_),
    .B(_2882_),
    .Y(_2883_)
);

INVX8 _13544_ (
    .A(areg_17_bF$buf4),
    .Y(_2884_)
);

OAI21X1 _13545_ (
    .A(_2551__bF$buf2),
    .B(_2884__bF$buf3),
    .C(_2881_),
    .Y(_2885_)
);

NAND3X1 _13546_ (
    .A(_2879_),
    .B(_2885_),
    .C(_2883_),
    .Y(_2886_)
);

NOR2X1 _13547_ (
    .A(_2881_),
    .B(_2882_),
    .Y(_2887_)
);

AND2X2 _13548_ (
    .A(_2881_),
    .B(_2882_),
    .Y(_2888_)
);

OAI21X1 _13549_ (
    .A(_2888_),
    .B(_2887_),
    .C(_2878_),
    .Y(_2889_)
);

NAND3X1 _13550_ (
    .A(_2886_),
    .B(_2889_),
    .C(_2877_),
    .Y(_2890_)
);

NOR3X1 _13551_ (
    .A(_2878_),
    .B(_2887_),
    .C(_2888_),
    .Y(_2891_)
);

AOI21X1 _13552_ (
    .A(_2885_),
    .B(_2883_),
    .C(_2879_),
    .Y(_2892_)
);

OAI21X1 _13553_ (
    .A(_2891_),
    .B(_2892_),
    .C(_2876_),
    .Y(_2893_)
);

NAND3X1 _13554_ (
    .A(_2875_),
    .B(_2893_),
    .C(_2890_),
    .Y(_2894_)
);

INVX2 _13555_ (
    .A(_2871_),
    .Y(_2895_)
);

XNOR2X1 _13556_ (
    .A(_2874_),
    .B(_2895_),
    .Y(_2896_)
);

NOR3X1 _13557_ (
    .A(_2892_),
    .B(_2876_),
    .C(_2891_),
    .Y(_2897_)
);

AOI21X1 _13558_ (
    .A(_2889_),
    .B(_2886_),
    .C(_2877_),
    .Y(_2898_)
);

OAI21X1 _13559_ (
    .A(_2898_),
    .B(_2897_),
    .C(_2896_),
    .Y(_2899_)
);

AOI21X1 _13560_ (
    .A(_2894_),
    .B(_2899_),
    .C(_2870_),
    .Y(_2900_)
);

AOI21X1 _13561_ (
    .A(_2659_),
    .B(_2678_),
    .C(_2681_),
    .Y(_2903_)
);

OAI21X1 _13562_ (
    .A(_2891_),
    .B(_2892_),
    .C(_2877_),
    .Y(_2904_)
);

NAND3X1 _13563_ (
    .A(_2876_),
    .B(_2889_),
    .C(_2886_),
    .Y(_2905_)
);

AOI21X1 _13564_ (
    .A(_2905_),
    .B(_2904_),
    .C(_2896_),
    .Y(_2906_)
);

AOI21X1 _13565_ (
    .A(_2893_),
    .B(_2890_),
    .C(_2875_),
    .Y(_2907_)
);

NOR3X1 _13566_ (
    .A(_2907_),
    .B(_2906_),
    .C(_2903_),
    .Y(_2908_)
);

OAI21X1 _13567_ (
    .A(_2908_),
    .B(_2900_),
    .C(_2868_),
    .Y(_2909_)
);

NAND3X1 _13568_ (
    .A(_2854_),
    .B(_2852_),
    .C(_2848_),
    .Y(_2910_)
);

OAI21X1 _13569_ (
    .A(_2860_),
    .B(_2859_),
    .C(_2855_),
    .Y(_2911_)
);

AOI21X1 _13570_ (
    .A(_2910_),
    .B(_2911_),
    .C(_2864_),
    .Y(_2912_)
);

AOI21X1 _13571_ (
    .A(_2856_),
    .B(_2861_),
    .C(_2843_),
    .Y(_2914_)
);

NOR2X1 _13572_ (
    .A(_2912_),
    .B(_2914_),
    .Y(_2915_)
);

OAI21X1 _13573_ (
    .A(_2907_),
    .B(_2906_),
    .C(_2903_),
    .Y(_2916_)
);

NAND3X1 _13574_ (
    .A(_2894_),
    .B(_2899_),
    .C(_2870_),
    .Y(_2917_)
);

NAND3X1 _13575_ (
    .A(_2916_),
    .B(_2917_),
    .C(_2915_),
    .Y(_2918_)
);

NAND3X1 _13576_ (
    .A(_2918_),
    .B(_2909_),
    .C(_2841_),
    .Y(_2919_)
);

AOI21X1 _13577_ (
    .A(_2695_),
    .B(_2693_),
    .C(_2691_),
    .Y(_2920_)
);

AOI21X1 _13578_ (
    .A(_2917_),
    .B(_2916_),
    .C(_2915_),
    .Y(_2921_)
);

NOR3X1 _13579_ (
    .A(_2868_),
    .B(_2900_),
    .C(_2908_),
    .Y(_2922_)
);

OAI21X1 _13580_ (
    .A(_2922_),
    .B(_2921_),
    .C(_2920_),
    .Y(_2923_)
);

NAND3X1 _13581_ (
    .A(_2919_),
    .B(_2923_),
    .C(_2840_),
    .Y(_2925_)
);

NAND3X1 _13582_ (
    .A(_2820_),
    .B(_2824_),
    .C(_2832_),
    .Y(_2926_)
);

OAI21X1 _13583_ (
    .A(_2829_),
    .B(_2830_),
    .C(_2827_),
    .Y(_2927_)
);

AOI21X1 _13584_ (
    .A(_2927_),
    .B(_2926_),
    .C(_2835_),
    .Y(_2928_)
);

AOI21X1 _13585_ (
    .A(_2833_),
    .B(_2828_),
    .C(_2794_),
    .Y(_2929_)
);

NOR2X1 _13586_ (
    .A(_2929_),
    .B(_2928_),
    .Y(_2930_)
);

OAI21X1 _13587_ (
    .A(_2922_),
    .B(_2921_),
    .C(_2841_),
    .Y(_2931_)
);

NAND3X1 _13588_ (
    .A(_2909_),
    .B(_2918_),
    .C(_2920_),
    .Y(_2932_)
);

NAND3X1 _13589_ (
    .A(_2931_),
    .B(_2932_),
    .C(_2930_),
    .Y(_2933_)
);

NAND3X1 _13590_ (
    .A(_2933_),
    .B(_2925_),
    .C(_2793_),
    .Y(_2934_)
);

NOR3X1 _13591_ (
    .A(_2699_),
    .B(_2700_),
    .C(_2701_),
    .Y(_2936_)
);

AOI21X1 _13592_ (
    .A(_2625_),
    .B(_2702_),
    .C(_2936_),
    .Y(_2937_)
);

AOI21X1 _13593_ (
    .A(_2931_),
    .B(_2932_),
    .C(_2930_),
    .Y(_2938_)
);

AOI21X1 _13594_ (
    .A(_2919_),
    .B(_2923_),
    .C(_2840_),
    .Y(_2939_)
);

OAI21X1 _13595_ (
    .A(_2939_),
    .B(_2938_),
    .C(_2937_),
    .Y(_2940_)
);

NAND3X1 _13596_ (
    .A(_2790_),
    .B(_2934_),
    .C(_2940_),
    .Y(_2941_)
);

NAND2X1 _13597_ (
    .A(_2786_),
    .B(_2789_),
    .Y(_2942_)
);

OAI21X1 _13598_ (
    .A(_2939_),
    .B(_2938_),
    .C(_2793_),
    .Y(_2943_)
);

NAND3X1 _13599_ (
    .A(_2925_),
    .B(_2933_),
    .C(_2937_),
    .Y(_2944_)
);

NAND3X1 _13600_ (
    .A(_2942_),
    .B(_2943_),
    .C(_2944_),
    .Y(_2945_)
);

NAND3X1 _13601_ (
    .A(_2941_),
    .B(_2945_),
    .C(_2760_),
    .Y(_2947_)
);

NOR3X1 _13602_ (
    .A(_2714_),
    .B(_2715_),
    .C(_2713_),
    .Y(_2948_)
);

AOI21X1 _13603_ (
    .A(_2577_),
    .B(_2717_),
    .C(_2948_),
    .Y(_2949_)
);

AOI21X1 _13604_ (
    .A(_2943_),
    .B(_2944_),
    .C(_2942_),
    .Y(_2950_)
);

AOI21X1 _13605_ (
    .A(_2934_),
    .B(_2940_),
    .C(_2790_),
    .Y(_2951_)
);

OAI21X1 _13606_ (
    .A(_2950_),
    .B(_2951_),
    .C(_2949_),
    .Y(_2952_)
);

NAND3X1 _13607_ (
    .A(_2757_),
    .B(_2947_),
    .C(_2952_),
    .Y(_2953_)
);

OAI21X1 _13608_ (
    .A(_2950_),
    .B(_2951_),
    .C(_2760_),
    .Y(_2954_)
);

NAND3X1 _13609_ (
    .A(_2941_),
    .B(_2945_),
    .C(_2949_),
    .Y(_2955_)
);

NAND3X1 _13610_ (
    .A(_2756_),
    .B(_2954_),
    .C(_2955_),
    .Y(_2956_)
);

NAND3X1 _13611_ (
    .A(_2953_),
    .B(_2956_),
    .C(_2755_),
    .Y(_2958_)
);

NOR3X1 _13612_ (
    .A(_2725_),
    .B(_2726_),
    .C(_2724_),
    .Y(_2959_)
);

AOI21X1 _13613_ (
    .A(_2554_),
    .B(_2728_),
    .C(_2959_),
    .Y(_2960_)
);

AOI21X1 _13614_ (
    .A(_2954_),
    .B(_2955_),
    .C(_2756_),
    .Y(_2961_)
);

AOI21X1 _13615_ (
    .A(_2947_),
    .B(_2952_),
    .C(_2757_),
    .Y(_2962_)
);

OAI21X1 _13616_ (
    .A(_2961_),
    .B(_2962_),
    .C(_2960_),
    .Y(_2963_)
);

NAND3X1 _13617_ (
    .A(_2958_),
    .B(_2963_),
    .C(_2753_),
    .Y(_2964_)
);

OAI21X1 _13618_ (
    .A(_2961_),
    .B(_2962_),
    .C(_2755_),
    .Y(_2965_)
);

NAND3X1 _13619_ (
    .A(_2953_),
    .B(_2956_),
    .C(_2960_),
    .Y(_2966_)
);

NAND3X1 _13620_ (
    .A(_2733_),
    .B(_2965_),
    .C(_2966_),
    .Y(_2967_)
);

NAND3X1 _13621_ (
    .A(_2752_),
    .B(_2967_),
    .C(_2964_),
    .Y(_2969_)
);

AOI21X1 _13622_ (
    .A(_2965_),
    .B(_2966_),
    .C(_2733_),
    .Y(_2970_)
);

NOR2X1 _13623_ (
    .A(_2737_),
    .B(_2736_),
    .Y(_2971_)
);

AOI22X1 _13624_ (
    .A(_2552_),
    .B(_2971_),
    .C(_2963_),
    .D(_2958_),
    .Y(_2972_)
);

OAI21X1 _13625_ (
    .A(_2970_),
    .B(_2972_),
    .C(_2740_),
    .Y(_2973_)
);

NAND2X1 _13626_ (
    .A(_2973_),
    .B(_2969_),
    .Y(_2974_)
);

XNOR2X1 _13627_ (
    .A(_2751_),
    .B(_2974_),
    .Y(_0_[17])
);

NOR2X1 _13628_ (
    .A(_2972_),
    .B(_2970_),
    .Y(_2975_)
);

NAND2X1 _13629_ (
    .A(_2744_),
    .B(_2969_),
    .Y(_2976_)
);

OAI21X1 _13630_ (
    .A(_2752_),
    .B(_2975_),
    .C(_2976_),
    .Y(_2977_)
);

OR2X2 _13631_ (
    .A(_2974_),
    .B(_2750_),
    .Y(_2979_)
);

OAI21X1 _13632_ (
    .A(_2545_),
    .B(_2979_),
    .C(_2977_),
    .Y(_2980_)
);

NOR3X1 _13633_ (
    .A(_2961_),
    .B(_2962_),
    .C(_2960_),
    .Y(_2981_)
);

AOI21X1 _13634_ (
    .A(_2941_),
    .B(_2945_),
    .C(_2760_),
    .Y(_2982_)
);

OAI21X1 _13635_ (
    .A(_2982_),
    .B(_2756_),
    .C(_2947_),
    .Y(_2983_)
);

OAI21X1 _13636_ (
    .A(_2783_),
    .B(_2784_),
    .C(_2786_),
    .Y(_2984_)
);

INVX2 _13637_ (
    .A(_2984_),
    .Y(_2985_)
);

AOI21X1 _13638_ (
    .A(_2933_),
    .B(_2925_),
    .C(_2793_),
    .Y(_2986_)
);

OAI21X1 _13639_ (
    .A(_2986_),
    .B(_2942_),
    .C(_2934_),
    .Y(_2987_)
);

NOR2X1 _13640_ (
    .A(_2566_),
    .B(_2778_),
    .Y(_2988_)
);

NAND2X1 _13641_ (
    .A(areg[0]),
    .B(breg_18_bF$buf5),
    .Y(_2990_)
);

OAI21X1 _13642_ (
    .A(_2558_),
    .B(_2765_),
    .C(_2767_),
    .Y(_2991_)
);

NOR2X1 _13643_ (
    .A(_2661_),
    .B(_2763_),
    .Y(_2992_)
);

NAND2X1 _13644_ (
    .A(areg_3_bF$buf1),
    .B(breg_15_bF$buf2),
    .Y(_2993_)
);

XOR2X1 _13645_ (
    .A(_2768_),
    .B(_2993_),
    .Y(_2994_)
);

NAND2X1 _13646_ (
    .A(_2992_),
    .B(_2994_),
    .Y(_2995_)
);

NAND2X1 _13647_ (
    .A(areg_3_bF$buf0),
    .B(breg_16_bF$buf2),
    .Y(_2996_)
);

OAI21X1 _13648_ (
    .A(_2792_),
    .B(_2362__bF$buf3),
    .C(_2768_),
    .Y(_2997_)
);

OAI21X1 _13649_ (
    .A(_2765_),
    .B(_2996_),
    .C(_2997_),
    .Y(_2998_)
);

OAI21X1 _13650_ (
    .A(_2661_),
    .B(_2763_),
    .C(_2998_),
    .Y(_2999_)
);

NAND2X1 _13651_ (
    .A(areg_5_bF$buf3),
    .B(breg_12_bF$buf3),
    .Y(_3001_)
);

NOR2X1 _13652_ (
    .A(_2797_),
    .B(_3001_),
    .Y(_3002_)
);

AOI21X1 _13653_ (
    .A(_2795_),
    .B(_2798_),
    .C(_3002_),
    .Y(_3003_)
);

INVX2 _13654_ (
    .A(_3003_),
    .Y(_3004_)
);

NAND3X1 _13655_ (
    .A(_2999_),
    .B(_3004_),
    .C(_2995_),
    .Y(_3005_)
);

INVX1 _13656_ (
    .A(_2992_),
    .Y(_3006_)
);

NOR2X1 _13657_ (
    .A(_3006_),
    .B(_2998_),
    .Y(_3007_)
);

NOR2X1 _13658_ (
    .A(_2992_),
    .B(_2994_),
    .Y(_3008_)
);

OAI21X1 _13659_ (
    .A(_3008_),
    .B(_3007_),
    .C(_3003_),
    .Y(_3009_)
);

NAND3X1 _13660_ (
    .A(_2991_),
    .B(_3005_),
    .C(_3009_),
    .Y(_3010_)
);

NOR2X1 _13661_ (
    .A(_2558_),
    .B(_2765_),
    .Y(_3012_)
);

INVX1 _13662_ (
    .A(_2764_),
    .Y(_3013_)
);

NOR2X1 _13663_ (
    .A(_3013_),
    .B(_2771_),
    .Y(_3014_)
);

NOR2X1 _13664_ (
    .A(_3012_),
    .B(_3014_),
    .Y(_3015_)
);

NAND3X1 _13665_ (
    .A(_3003_),
    .B(_2999_),
    .C(_2995_),
    .Y(_3016_)
);

OAI21X1 _13666_ (
    .A(_3008_),
    .B(_3007_),
    .C(_3004_),
    .Y(_3017_)
);

NAND3X1 _13667_ (
    .A(_3015_),
    .B(_3016_),
    .C(_3017_),
    .Y(_3018_)
);

AOI21X1 _13668_ (
    .A(_2559_),
    .B(_2775_),
    .C(_2776_),
    .Y(_3019_)
);

AOI21X1 _13669_ (
    .A(_3018_),
    .B(_3010_),
    .C(_3019_),
    .Y(_3020_)
);

AOI21X1 _13670_ (
    .A(_3016_),
    .B(_3017_),
    .C(_3015_),
    .Y(_3021_)
);

AOI21X1 _13671_ (
    .A(_3005_),
    .B(_3009_),
    .C(_2991_),
    .Y(_3023_)
);

INVX1 _13672_ (
    .A(_2559_),
    .Y(_3024_)
);

NOR2X1 _13673_ (
    .A(_2764_),
    .B(_2766_),
    .Y(_3025_)
);

NOR3X1 _13674_ (
    .A(_3014_),
    .B(_2773_),
    .C(_3025_),
    .Y(_3026_)
);

OAI21X1 _13675_ (
    .A(_3026_),
    .B(_3024_),
    .C(_2777_),
    .Y(_3027_)
);

NOR3X1 _13676_ (
    .A(_3021_),
    .B(_3023_),
    .C(_3027_),
    .Y(_3028_)
);

OAI21X1 _13677_ (
    .A(_3028_),
    .B(_3020_),
    .C(_2990_),
    .Y(_3029_)
);

INVX1 _13678_ (
    .A(_2990_),
    .Y(_3030_)
);

OAI21X1 _13679_ (
    .A(_3021_),
    .B(_3023_),
    .C(_3027_),
    .Y(_3031_)
);

NAND3X1 _13680_ (
    .A(_3019_),
    .B(_3010_),
    .C(_3018_),
    .Y(_3032_)
);

NAND3X1 _13681_ (
    .A(_3030_),
    .B(_3032_),
    .C(_3031_),
    .Y(_3034_)
);

OAI21X1 _13682_ (
    .A(_2838_),
    .B(_2794_),
    .C(_2828_),
    .Y(_3035_)
);

NAND3X1 _13683_ (
    .A(_3034_),
    .B(_3035_),
    .C(_3029_),
    .Y(_3036_)
);

AOI21X1 _13684_ (
    .A(_3032_),
    .B(_3031_),
    .C(_3030_),
    .Y(_3037_)
);

NOR3X1 _13685_ (
    .A(_2990_),
    .B(_3020_),
    .C(_3028_),
    .Y(_3038_)
);

AOI21X1 _13686_ (
    .A(_2835_),
    .B(_2833_),
    .C(_2837_),
    .Y(_3039_)
);

OAI21X1 _13687_ (
    .A(_3038_),
    .B(_3037_),
    .C(_3039_),
    .Y(_3040_)
);

NAND3X1 _13688_ (
    .A(_2988_),
    .B(_3036_),
    .C(_3040_),
    .Y(_3041_)
);

INVX1 _13689_ (
    .A(_2988_),
    .Y(_3042_)
);

NAND3X1 _13690_ (
    .A(_3034_),
    .B(_3029_),
    .C(_3039_),
    .Y(_3043_)
);

OAI21X1 _13691_ (
    .A(_3038_),
    .B(_3037_),
    .C(_3035_),
    .Y(_3045_)
);

NAND3X1 _13692_ (
    .A(_3042_),
    .B(_3043_),
    .C(_3045_),
    .Y(_3046_)
);

NAND2X1 _13693_ (
    .A(_3041_),
    .B(_3046_),
    .Y(_3047_)
);

AOI21X1 _13694_ (
    .A(_2918_),
    .B(_2909_),
    .C(_2841_),
    .Y(_3048_)
);

OAI21X1 _13695_ (
    .A(_2930_),
    .B(_3048_),
    .C(_2919_),
    .Y(_3049_)
);

AOI21X1 _13696_ (
    .A(_2805_),
    .B(_2810_),
    .C(_2829_),
    .Y(_3050_)
);

NOR2X1 _13697_ (
    .A(_2562__bF$buf0),
    .B(_2379_),
    .Y(_3051_)
);

INVX1 _13698_ (
    .A(_3051_),
    .Y(_3052_)
);

NAND2X1 _13699_ (
    .A(areg_6_bF$buf4),
    .B(breg_12_bF$buf2),
    .Y(_3053_)
);

NOR2X1 _13700_ (
    .A(_2796_),
    .B(_3053_),
    .Y(_3054_)
);

AND2X2 _13701_ (
    .A(_2796_),
    .B(_3053_),
    .Y(_3056_)
);

NOR2X1 _13702_ (
    .A(_3054_),
    .B(_3056_),
    .Y(_3057_)
);

XNOR2X1 _13703_ (
    .A(_3057_),
    .B(_3052_),
    .Y(_3058_)
);

AOI21X1 _13704_ (
    .A(_2806_),
    .B(_2808_),
    .C(_2816_),
    .Y(_3059_)
);

INVX1 _13705_ (
    .A(_3059_),
    .Y(_3060_)
);

NOR2X1 _13706_ (
    .A(_4434__bF$buf1),
    .B(_8555_),
    .Y(_3061_)
);

NAND2X1 _13707_ (
    .A(areg_9_bF$buf1),
    .B(breg_9_bF$buf1),
    .Y(_3062_)
);

NOR2X1 _13708_ (
    .A(_2807_),
    .B(_3062_),
    .Y(_3063_)
);

AND2X2 _13709_ (
    .A(_2807_),
    .B(_3062_),
    .Y(_3064_)
);

NOR2X1 _13710_ (
    .A(_3063_),
    .B(_3064_),
    .Y(_3065_)
);

NAND2X1 _13711_ (
    .A(_3061_),
    .B(_3065_),
    .Y(_3067_)
);

INVX1 _13712_ (
    .A(_3061_),
    .Y(_3068_)
);

OAI21X1 _13713_ (
    .A(_3064_),
    .B(_3063_),
    .C(_3068_),
    .Y(_3069_)
);

NAND3X1 _13714_ (
    .A(_3069_),
    .B(_3060_),
    .C(_3067_),
    .Y(_3070_)
);

NAND2X1 _13715_ (
    .A(areg_9_bF$buf0),
    .B(breg_10_bF$buf0),
    .Y(_3071_)
);

OAI21X1 _13716_ (
    .A(_6582__bF$buf2),
    .B(_6044__bF$buf4),
    .C(_2807_),
    .Y(_3072_)
);

OAI21X1 _13717_ (
    .A(_2815_),
    .B(_3071_),
    .C(_3072_),
    .Y(_3073_)
);

NOR2X1 _13718_ (
    .A(_3068_),
    .B(_3073_),
    .Y(_3074_)
);

INVX1 _13719_ (
    .A(_3069_),
    .Y(_3075_)
);

OAI21X1 _13720_ (
    .A(_3075_),
    .B(_3074_),
    .C(_3059_),
    .Y(_3076_)
);

NAND3X1 _13721_ (
    .A(_3058_),
    .B(_3070_),
    .C(_3076_),
    .Y(_3078_)
);

INVX1 _13722_ (
    .A(_3058_),
    .Y(_3079_)
);

OAI21X1 _13723_ (
    .A(_3075_),
    .B(_3074_),
    .C(_3060_),
    .Y(_3080_)
);

NAND3X1 _13724_ (
    .A(_3059_),
    .B(_3069_),
    .C(_3067_),
    .Y(_3081_)
);

NAND3X1 _13725_ (
    .A(_3080_),
    .B(_3081_),
    .C(_3079_),
    .Y(_3082_)
);

OAI21X1 _13726_ (
    .A(_2864_),
    .B(_2866_),
    .C(_2856_),
    .Y(_3083_)
);

NAND3X1 _13727_ (
    .A(_3083_),
    .B(_3078_),
    .C(_3082_),
    .Y(_3084_)
);

AOI21X1 _13728_ (
    .A(_3081_),
    .B(_3080_),
    .C(_3079_),
    .Y(_3085_)
);

AOI21X1 _13729_ (
    .A(_3070_),
    .B(_3076_),
    .C(_3058_),
    .Y(_3086_)
);

AOI21X1 _13730_ (
    .A(_2843_),
    .B(_2861_),
    .C(_2865_),
    .Y(_3087_)
);

OAI21X1 _13731_ (
    .A(_3085_),
    .B(_3086_),
    .C(_3087_),
    .Y(_3089_)
);

NAND3X1 _13732_ (
    .A(_3050_),
    .B(_3084_),
    .C(_3089_),
    .Y(_3090_)
);

NAND2X1 _13733_ (
    .A(_2811_),
    .B(_2820_),
    .Y(_3091_)
);

NAND3X1 _13734_ (
    .A(_3087_),
    .B(_3078_),
    .C(_3082_),
    .Y(_3092_)
);

OAI21X1 _13735_ (
    .A(_3085_),
    .B(_3086_),
    .C(_3083_),
    .Y(_3093_)
);

NAND3X1 _13736_ (
    .A(_3091_),
    .B(_3092_),
    .C(_3093_),
    .Y(_3094_)
);

AND2X2 _13737_ (
    .A(_3090_),
    .B(_3094_),
    .Y(_3095_)
);

OAI21X1 _13738_ (
    .A(_2868_),
    .B(_2900_),
    .C(_2917_),
    .Y(_3096_)
);

NOR2X1 _13739_ (
    .A(_2631_),
    .B(_2845_),
    .Y(_3097_)
);

NOR2X1 _13740_ (
    .A(_3097_),
    .B(_2859_),
    .Y(_3098_)
);

NAND2X1 _13741_ (
    .A(breg[8]),
    .B(areg_10_bF$buf1),
    .Y(_3100_)
);

INVX1 _13742_ (
    .A(_3100_),
    .Y(_3101_)
);

AND2X2 _13743_ (
    .A(breg_7_bF$buf4),
    .B(areg_11_bF$buf1),
    .Y(_3102_)
);

AND2X2 _13744_ (
    .A(breg_6_bF$buf3),
    .B(areg_12_bF$buf1),
    .Y(_3103_)
);

NAND2X1 _13745_ (
    .A(_3102_),
    .B(_3103_),
    .Y(_3104_)
);

OAI21X1 _13746_ (
    .A(_5453__bF$buf3),
    .B(_10869__bF$buf2),
    .C(_2849_),
    .Y(_3105_)
);

NAND3X1 _13747_ (
    .A(_3101_),
    .B(_3105_),
    .C(_3104_),
    .Y(_3106_)
);

OAI21X1 _13748_ (
    .A(_4116__bF$buf2),
    .B(_9104__bF$buf2),
    .C(_3103_),
    .Y(_3107_)
);

OAI21X1 _13749_ (
    .A(_5453__bF$buf2),
    .B(_10869__bF$buf1),
    .C(_3102_),
    .Y(_3108_)
);

NAND3X1 _13750_ (
    .A(_3100_),
    .B(_3107_),
    .C(_3108_),
    .Y(_3109_)
);

NAND2X1 _13751_ (
    .A(breg_4_bF$buf2),
    .B(areg_14_bF$buf4),
    .Y(_3111_)
);

AND2X2 _13752_ (
    .A(_2872_),
    .B(_2873_),
    .Y(_3112_)
);

OAI22X1 _13753_ (
    .A(_2655_),
    .B(_3111_),
    .C(_3112_),
    .D(_2871_),
    .Y(_3113_)
);

NAND3X1 _13754_ (
    .A(_3106_),
    .B(_3109_),
    .C(_3113_),
    .Y(_3114_)
);

AOI21X1 _13755_ (
    .A(_3107_),
    .B(_3108_),
    .C(_3100_),
    .Y(_3115_)
);

AOI21X1 _13756_ (
    .A(_3105_),
    .B(_3104_),
    .C(_3101_),
    .Y(_3116_)
);

NOR2X1 _13757_ (
    .A(_2872_),
    .B(_2873_),
    .Y(_3117_)
);

OAI21X1 _13758_ (
    .A(_2365_),
    .B(_2287__bF$buf2),
    .C(_2872_),
    .Y(_3118_)
);

AOI21X1 _13759_ (
    .A(_2895_),
    .B(_3118_),
    .C(_3117_),
    .Y(_3119_)
);

OAI21X1 _13760_ (
    .A(_3115_),
    .B(_3116_),
    .C(_3119_),
    .Y(_3120_)
);

NAND3X1 _13761_ (
    .A(_3114_),
    .B(_3120_),
    .C(_3098_),
    .Y(_3121_)
);

OAI21X1 _13762_ (
    .A(_2638_),
    .B(_2849_),
    .C(_2848_),
    .Y(_3122_)
);

NOR3X1 _13763_ (
    .A(_3116_),
    .B(_3119_),
    .C(_3115_),
    .Y(_3123_)
);

AOI21X1 _13764_ (
    .A(_3106_),
    .B(_3109_),
    .C(_3113_),
    .Y(_3124_)
);

OAI21X1 _13765_ (
    .A(_3123_),
    .B(_3124_),
    .C(_3122_),
    .Y(_3125_)
);

NAND2X1 _13766_ (
    .A(_3125_),
    .B(_3121_),
    .Y(_3126_)
);

INVX2 _13767_ (
    .A(_3126_),
    .Y(_3127_)
);

OAI21X1 _13768_ (
    .A(_2898_),
    .B(_2896_),
    .C(_2890_),
    .Y(_3128_)
);

NOR2X1 _13769_ (
    .A(_4258__bF$buf1),
    .B(_549__bF$buf2),
    .Y(_3129_)
);

NAND2X1 _13770_ (
    .A(breg_3_bF$buf3),
    .B(areg_15_bF$buf0),
    .Y(_3130_)
);

OR2X2 _13771_ (
    .A(_3111_),
    .B(_3130_),
    .Y(_3132_)
);

OAI21X1 _13772_ (
    .A(_2365_),
    .B(_2465__bF$buf3),
    .C(_3111_),
    .Y(_3133_)
);

NAND3X1 _13773_ (
    .A(_3129_),
    .B(_3133_),
    .C(_3132_),
    .Y(_3134_)
);

INVX1 _13774_ (
    .A(_3129_),
    .Y(_3135_)
);

NOR2X1 _13775_ (
    .A(_3111_),
    .B(_3130_),
    .Y(_3136_)
);

AND2X2 _13776_ (
    .A(_3111_),
    .B(_3130_),
    .Y(_3137_)
);

OAI21X1 _13777_ (
    .A(_3137_),
    .B(_3136_),
    .C(_3135_),
    .Y(_3138_)
);

NAND2X1 _13778_ (
    .A(_3134_),
    .B(_3138_),
    .Y(_3139_)
);

OAI21X1 _13779_ (
    .A(_2888_),
    .B(_2878_),
    .C(_2883_),
    .Y(_3140_)
);

NAND2X1 _13780_ (
    .A(breg_2_bF$buf0),
    .B(areg_16_bF$buf2),
    .Y(_3141_)
);

AND2X2 _13781_ (
    .A(breg_0_bF$buf1),
    .B(areg_18_bF$buf5),
    .Y(_3144_)
);

OAI21X1 _13782_ (
    .A(_3220_),
    .B(_2884__bF$buf2),
    .C(_3144_),
    .Y(_3145_)
);

INVX8 _13783_ (
    .A(areg_18_bF$buf4),
    .Y(_3146_)
);

AND2X2 _13784_ (
    .A(breg_1_bF$buf2),
    .B(areg_17_bF$buf3),
    .Y(_3147_)
);

OAI21X1 _13785_ (
    .A(_2551__bF$buf1),
    .B(_3146__bF$buf3),
    .C(_3147_),
    .Y(_3148_)
);

AOI21X1 _13786_ (
    .A(_3145_),
    .B(_3148_),
    .C(_3141_),
    .Y(_3149_)
);

INVX2 _13787_ (
    .A(_3141_),
    .Y(_3150_)
);

NAND2X1 _13788_ (
    .A(_3147_),
    .B(_3144_),
    .Y(_3151_)
);

NAND2X1 _13789_ (
    .A(breg_1_bF$buf1),
    .B(areg_17_bF$buf2),
    .Y(_3152_)
);

OAI21X1 _13790_ (
    .A(_2551__bF$buf0),
    .B(_3146__bF$buf2),
    .C(_3152_),
    .Y(_3153_)
);

AOI21X1 _13791_ (
    .A(_3153_),
    .B(_3151_),
    .C(_3150_),
    .Y(_3155_)
);

OAI21X1 _13792_ (
    .A(_3149_),
    .B(_3155_),
    .C(_3140_),
    .Y(_3156_)
);

AOI21X1 _13793_ (
    .A(_2879_),
    .B(_2885_),
    .C(_2887_),
    .Y(_3157_)
);

NAND3X1 _13794_ (
    .A(_3150_),
    .B(_3153_),
    .C(_3151_),
    .Y(_3158_)
);

NAND2X1 _13795_ (
    .A(breg_0_bF$buf0),
    .B(areg_18_bF$buf3),
    .Y(_3159_)
);

NOR2X1 _13796_ (
    .A(_3152_),
    .B(_3159_),
    .Y(_3160_)
);

NOR2X1 _13797_ (
    .A(_3147_),
    .B(_3144_),
    .Y(_3161_)
);

OAI21X1 _13798_ (
    .A(_3161_),
    .B(_3160_),
    .C(_3141_),
    .Y(_3162_)
);

NAND3X1 _13799_ (
    .A(_3157_),
    .B(_3158_),
    .C(_3162_),
    .Y(_3163_)
);

AOI21X1 _13800_ (
    .A(_3156_),
    .B(_3163_),
    .C(_3139_),
    .Y(_3164_)
);

AND2X2 _13801_ (
    .A(_3138_),
    .B(_3134_),
    .Y(_3166_)
);

NAND3X1 _13802_ (
    .A(_3158_),
    .B(_3140_),
    .C(_3162_),
    .Y(_3167_)
);

OAI21X1 _13803_ (
    .A(_3149_),
    .B(_3155_),
    .C(_3157_),
    .Y(_3168_)
);

AOI21X1 _13804_ (
    .A(_3168_),
    .B(_3167_),
    .C(_3166_),
    .Y(_3169_)
);

OAI21X1 _13805_ (
    .A(_3164_),
    .B(_3169_),
    .C(_3128_),
    .Y(_3170_)
);

AOI21X1 _13806_ (
    .A(_2893_),
    .B(_2875_),
    .C(_2897_),
    .Y(_3171_)
);

NAND3X1 _13807_ (
    .A(_3168_),
    .B(_3167_),
    .C(_3166_),
    .Y(_3172_)
);

NOR3X1 _13808_ (
    .A(_3155_),
    .B(_3157_),
    .C(_3149_),
    .Y(_3173_)
);

AOI21X1 _13809_ (
    .A(_3158_),
    .B(_3162_),
    .C(_3140_),
    .Y(_3174_)
);

OAI21X1 _13810_ (
    .A(_3173_),
    .B(_3174_),
    .C(_3139_),
    .Y(_3175_)
);

NAND3X1 _13811_ (
    .A(_3172_),
    .B(_3175_),
    .C(_3171_),
    .Y(_3177_)
);

AOI21X1 _13812_ (
    .A(_3177_),
    .B(_3170_),
    .C(_3127_),
    .Y(_3178_)
);

NAND3X1 _13813_ (
    .A(_3172_),
    .B(_3175_),
    .C(_3128_),
    .Y(_3179_)
);

OAI21X1 _13814_ (
    .A(_3164_),
    .B(_3169_),
    .C(_3171_),
    .Y(_3180_)
);

AOI21X1 _13815_ (
    .A(_3180_),
    .B(_3179_),
    .C(_3126_),
    .Y(_3181_)
);

OAI21X1 _13816_ (
    .A(_3178_),
    .B(_3181_),
    .C(_3096_),
    .Y(_3182_)
);

AOI21X1 _13817_ (
    .A(_2916_),
    .B(_2915_),
    .C(_2908_),
    .Y(_3183_)
);

NAND3X1 _13818_ (
    .A(_3126_),
    .B(_3180_),
    .C(_3179_),
    .Y(_3184_)
);

NOR3X1 _13819_ (
    .A(_3164_),
    .B(_3169_),
    .C(_3171_),
    .Y(_3185_)
);

AOI21X1 _13820_ (
    .A(_3172_),
    .B(_3175_),
    .C(_3128_),
    .Y(_3186_)
);

OAI21X1 _13821_ (
    .A(_3185_),
    .B(_3186_),
    .C(_3127_),
    .Y(_3188_)
);

NAND3X1 _13822_ (
    .A(_3184_),
    .B(_3188_),
    .C(_3183_),
    .Y(_3189_)
);

AOI21X1 _13823_ (
    .A(_3182_),
    .B(_3189_),
    .C(_3095_),
    .Y(_3190_)
);

NAND2X1 _13824_ (
    .A(_3094_),
    .B(_3090_),
    .Y(_3191_)
);

NAND3X1 _13825_ (
    .A(_3184_),
    .B(_3188_),
    .C(_3096_),
    .Y(_3192_)
);

OAI21X1 _13826_ (
    .A(_3178_),
    .B(_3181_),
    .C(_3183_),
    .Y(_3193_)
);

AOI21X1 _13827_ (
    .A(_3192_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3194_)
);

OAI21X1 _13828_ (
    .A(_3190_),
    .B(_3194_),
    .C(_3049_),
    .Y(_3195_)
);

NOR3X1 _13829_ (
    .A(_2922_),
    .B(_2921_),
    .C(_2920_),
    .Y(_3196_)
);

AOI21X1 _13830_ (
    .A(_2923_),
    .B(_2840_),
    .C(_3196_),
    .Y(_3197_)
);

NAND3X1 _13831_ (
    .A(_3192_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3199_)
);

NOR3X1 _13832_ (
    .A(_3183_),
    .B(_3181_),
    .C(_3178_),
    .Y(_3200_)
);

AOI21X1 _13833_ (
    .A(_3184_),
    .B(_3188_),
    .C(_3096_),
    .Y(_3201_)
);

OAI21X1 _13834_ (
    .A(_3200_),
    .B(_3201_),
    .C(_3095_),
    .Y(_3202_)
);

NAND3X1 _13835_ (
    .A(_3199_),
    .B(_3202_),
    .C(_3197_),
    .Y(_3203_)
);

AOI21X1 _13836_ (
    .A(_3195_),
    .B(_3203_),
    .C(_3047_),
    .Y(_3204_)
);

NAND3X1 _13837_ (
    .A(_3042_),
    .B(_3036_),
    .C(_3040_),
    .Y(_3205_)
);

NAND3X1 _13838_ (
    .A(_2988_),
    .B(_3043_),
    .C(_3045_),
    .Y(_3206_)
);

NAND2X1 _13839_ (
    .A(_3205_),
    .B(_3206_),
    .Y(_3207_)
);

NAND3X1 _13840_ (
    .A(_3199_),
    .B(_3202_),
    .C(_3049_),
    .Y(_3208_)
);

OAI21X1 _13841_ (
    .A(_3190_),
    .B(_3194_),
    .C(_3197_),
    .Y(_3210_)
);

AOI21X1 _13842_ (
    .A(_3210_),
    .B(_3208_),
    .C(_3207_),
    .Y(_3211_)
);

OAI21X1 _13843_ (
    .A(_3204_),
    .B(_3211_),
    .C(_2987_),
    .Y(_3212_)
);

NOR3X1 _13844_ (
    .A(_2938_),
    .B(_2939_),
    .C(_2937_),
    .Y(_3213_)
);

AOI21X1 _13845_ (
    .A(_2790_),
    .B(_2940_),
    .C(_3213_),
    .Y(_3214_)
);

NAND3X1 _13846_ (
    .A(_3208_),
    .B(_3210_),
    .C(_3207_),
    .Y(_3215_)
);

NAND3X1 _13847_ (
    .A(_3195_),
    .B(_3203_),
    .C(_3047_),
    .Y(_3216_)
);

NAND3X1 _13848_ (
    .A(_3215_),
    .B(_3216_),
    .C(_3214_),
    .Y(_3217_)
);

AOI21X1 _13849_ (
    .A(_3212_),
    .B(_3217_),
    .C(_2985_),
    .Y(_3218_)
);

NAND3X1 _13850_ (
    .A(_3215_),
    .B(_3216_),
    .C(_2987_),
    .Y(_3219_)
);

OAI21X1 _13851_ (
    .A(_3204_),
    .B(_3211_),
    .C(_3214_),
    .Y(_3221_)
);

AOI21X1 _13852_ (
    .A(_3219_),
    .B(_3221_),
    .C(_2984_),
    .Y(_3222_)
);

OAI21X1 _13853_ (
    .A(_3218_),
    .B(_3222_),
    .C(_2983_),
    .Y(_3223_)
);

NOR3X1 _13854_ (
    .A(_2950_),
    .B(_2951_),
    .C(_2949_),
    .Y(_3224_)
);

AOI21X1 _13855_ (
    .A(_2757_),
    .B(_2952_),
    .C(_3224_),
    .Y(_3225_)
);

NAND3X1 _13856_ (
    .A(_2984_),
    .B(_3219_),
    .C(_3221_),
    .Y(_3226_)
);

NAND3X1 _13857_ (
    .A(_2985_),
    .B(_3212_),
    .C(_3217_),
    .Y(_3227_)
);

NAND3X1 _13858_ (
    .A(_3226_),
    .B(_3227_),
    .C(_3225_),
    .Y(_3228_)
);

AOI21X1 _13859_ (
    .A(_3223_),
    .B(_3228_),
    .C(_2981_),
    .Y(_3229_)
);

NAND3X1 _13860_ (
    .A(_3226_),
    .B(_2983_),
    .C(_3227_),
    .Y(_3230_)
);

OAI21X1 _13861_ (
    .A(_3218_),
    .B(_3222_),
    .C(_3225_),
    .Y(_3232_)
);

AOI21X1 _13862_ (
    .A(_3230_),
    .B(_3232_),
    .C(_2958_),
    .Y(_3233_)
);

OAI21X1 _13863_ (
    .A(_3229_),
    .B(_3233_),
    .C(_2964_),
    .Y(_3234_)
);

AOI21X1 _13864_ (
    .A(_3223_),
    .B(_3228_),
    .C(_2958_),
    .Y(_3235_)
);

AOI21X1 _13865_ (
    .A(_3230_),
    .B(_3232_),
    .C(_2981_),
    .Y(_3236_)
);

OAI21X1 _13866_ (
    .A(_3236_),
    .B(_3235_),
    .C(_2970_),
    .Y(_3237_)
);

NAND2X1 _13867_ (
    .A(_3234_),
    .B(_3237_),
    .Y(_3238_)
);

XOR2X1 _13868_ (
    .A(_2980_),
    .B(_3238_),
    .Y(_0_[18])
);

OAI21X1 _13869_ (
    .A(_3229_),
    .B(_3233_),
    .C(_2970_),
    .Y(_3239_)
);

INVX1 _13870_ (
    .A(_3239_),
    .Y(_3240_)
);

AOI21X1 _13871_ (
    .A(_3238_),
    .B(_2980_),
    .C(_3240_),
    .Y(_3242_)
);

NOR3X1 _13872_ (
    .A(_3218_),
    .B(_3222_),
    .C(_3225_),
    .Y(_3243_)
);

AOI21X1 _13873_ (
    .A(_3215_),
    .B(_3216_),
    .C(_2987_),
    .Y(_3244_)
);

OAI21X1 _13874_ (
    .A(_3244_),
    .B(_2985_),
    .C(_3219_),
    .Y(_3245_)
);

NAND2X1 _13875_ (
    .A(_3036_),
    .B(_3041_),
    .Y(_3246_)
);

AOI21X1 _13876_ (
    .A(_3199_),
    .B(_3202_),
    .C(_3049_),
    .Y(_3247_)
);

OAI21X1 _13877_ (
    .A(_3047_),
    .B(_3247_),
    .C(_3208_),
    .Y(_3248_)
);

OAI21X1 _13878_ (
    .A(_3020_),
    .B(_2990_),
    .C(_3032_),
    .Y(_3249_)
);

INVX1 _13879_ (
    .A(_3249_),
    .Y(_3250_)
);

NAND2X1 _13880_ (
    .A(areg_1_bF$buf2),
    .B(breg_19_bF$buf5),
    .Y(_3251_)
);

INVX8 _13881_ (
    .A(breg_19_bF$buf4),
    .Y(_3253_)
);

NAND2X1 _13882_ (
    .A(areg_1_bF$buf1),
    .B(breg_18_bF$buf4),
    .Y(_3254_)
);

OAI21X1 _13883_ (
    .A(_2376__bF$buf1),
    .B(_3253__bF$buf3),
    .C(_3254_),
    .Y(_3255_)
);

OAI21X1 _13884_ (
    .A(_2990_),
    .B(_3251_),
    .C(_3255_),
    .Y(_3256_)
);

INVX2 _13885_ (
    .A(_3256_),
    .Y(_3257_)
);

AOI21X1 _13886_ (
    .A(_2999_),
    .B(_2995_),
    .C(_3004_),
    .Y(_3258_)
);

OAI21X1 _13887_ (
    .A(_3258_),
    .B(_3015_),
    .C(_3005_),
    .Y(_3259_)
);

OAI21X1 _13888_ (
    .A(_2765_),
    .B(_2996_),
    .C(_2995_),
    .Y(_3260_)
);

NOR2X1 _13889_ (
    .A(_2519__bF$buf1),
    .B(_2763_),
    .Y(_3261_)
);

NAND2X1 _13890_ (
    .A(areg_4_bF$buf2),
    .B(breg_15_bF$buf1),
    .Y(_3262_)
);

XOR2X1 _13891_ (
    .A(_2996_),
    .B(_3262_),
    .Y(_3264_)
);

NAND2X1 _13892_ (
    .A(_3261_),
    .B(_3264_),
    .Y(_3265_)
);

NAND2X1 _13893_ (
    .A(areg_4_bF$buf1),
    .B(breg_16_bF$buf1),
    .Y(_3266_)
);

OAI21X1 _13894_ (
    .A(_2562__bF$buf4),
    .B(_2362__bF$buf2),
    .C(_2996_),
    .Y(_3267_)
);

OAI21X1 _13895_ (
    .A(_2993_),
    .B(_3266_),
    .C(_3267_),
    .Y(_3268_)
);

OAI21X1 _13896_ (
    .A(_2519__bF$buf0),
    .B(_2763_),
    .C(_3268_),
    .Y(_3269_)
);

OAI21X1 _13897_ (
    .A(_3646__bF$buf0),
    .B(_2586__bF$buf2),
    .C(_2796_),
    .Y(_3270_)
);

AOI21X1 _13898_ (
    .A(_3051_),
    .B(_3270_),
    .C(_3054_),
    .Y(_3271_)
);

INVX1 _13899_ (
    .A(_3271_),
    .Y(_3272_)
);

NAND3X1 _13900_ (
    .A(_3269_),
    .B(_3272_),
    .C(_3265_),
    .Y(_3273_)
);

INVX1 _13901_ (
    .A(_3261_),
    .Y(_3275_)
);

NOR2X1 _13902_ (
    .A(_3275_),
    .B(_3268_),
    .Y(_3276_)
);

NOR2X1 _13903_ (
    .A(_3261_),
    .B(_3264_),
    .Y(_3277_)
);

OAI21X1 _13904_ (
    .A(_3277_),
    .B(_3276_),
    .C(_3271_),
    .Y(_3278_)
);

NAND3X1 _13905_ (
    .A(_3260_),
    .B(_3273_),
    .C(_3278_),
    .Y(_3279_)
);

NOR2X1 _13906_ (
    .A(_2768_),
    .B(_2993_),
    .Y(_3280_)
);

NOR2X1 _13907_ (
    .A(_3280_),
    .B(_3007_),
    .Y(_3281_)
);

NOR3X1 _13908_ (
    .A(_3276_),
    .B(_3271_),
    .C(_3277_),
    .Y(_3282_)
);

AOI21X1 _13909_ (
    .A(_3269_),
    .B(_3265_),
    .C(_3272_),
    .Y(_3283_)
);

OAI21X1 _13910_ (
    .A(_3282_),
    .B(_3283_),
    .C(_3281_),
    .Y(_3284_)
);

NAND3X1 _13911_ (
    .A(_3259_),
    .B(_3279_),
    .C(_3284_),
    .Y(_3286_)
);

INVX1 _13912_ (
    .A(_3259_),
    .Y(_3287_)
);

NOR3X1 _13913_ (
    .A(_3281_),
    .B(_3283_),
    .C(_3282_),
    .Y(_3288_)
);

AOI21X1 _13914_ (
    .A(_3273_),
    .B(_3278_),
    .C(_3260_),
    .Y(_3289_)
);

OAI21X1 _13915_ (
    .A(_3288_),
    .B(_3289_),
    .C(_3287_),
    .Y(_3290_)
);

NAND3X1 _13916_ (
    .A(_3257_),
    .B(_3286_),
    .C(_3290_),
    .Y(_3291_)
);

OAI21X1 _13917_ (
    .A(_3288_),
    .B(_3289_),
    .C(_3259_),
    .Y(_3292_)
);

NAND3X1 _13918_ (
    .A(_3279_),
    .B(_3284_),
    .C(_3287_),
    .Y(_3293_)
);

NAND3X1 _13919_ (
    .A(_3256_),
    .B(_3292_),
    .C(_3293_),
    .Y(_3294_)
);

AOI21X1 _13920_ (
    .A(_3078_),
    .B(_3082_),
    .C(_3083_),
    .Y(_3295_)
);

OAI21X1 _13921_ (
    .A(_3295_),
    .B(_3050_),
    .C(_3084_),
    .Y(_3297_)
);

NAND3X1 _13922_ (
    .A(_3291_),
    .B(_3297_),
    .C(_3294_),
    .Y(_3298_)
);

AOI21X1 _13923_ (
    .A(_3292_),
    .B(_3293_),
    .C(_3256_),
    .Y(_3299_)
);

AOI21X1 _13924_ (
    .A(_3286_),
    .B(_3290_),
    .C(_3257_),
    .Y(_3300_)
);

NOR3X1 _13925_ (
    .A(_3086_),
    .B(_3087_),
    .C(_3085_),
    .Y(_3301_)
);

AOI21X1 _13926_ (
    .A(_3091_),
    .B(_3089_),
    .C(_3301_),
    .Y(_3302_)
);

OAI21X1 _13927_ (
    .A(_3299_),
    .B(_3300_),
    .C(_3302_),
    .Y(_3303_)
);

NAND3X1 _13928_ (
    .A(_3298_),
    .B(_3250_),
    .C(_3303_),
    .Y(_3304_)
);

NAND3X1 _13929_ (
    .A(_3291_),
    .B(_3302_),
    .C(_3294_),
    .Y(_3305_)
);

OAI21X1 _13930_ (
    .A(_3299_),
    .B(_3300_),
    .C(_3297_),
    .Y(_3306_)
);

NAND3X1 _13931_ (
    .A(_3249_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3308_)
);

NAND2X1 _13932_ (
    .A(_3308_),
    .B(_3304_),
    .Y(_3309_)
);

OAI21X1 _13933_ (
    .A(_3095_),
    .B(_3201_),
    .C(_3192_),
    .Y(_3310_)
);

NAND2X1 _13934_ (
    .A(_3070_),
    .B(_3078_),
    .Y(_3311_)
);

NOR2X1 _13935_ (
    .A(_2825__bF$buf0),
    .B(_2379_),
    .Y(_3312_)
);

INVX1 _13936_ (
    .A(_3312_),
    .Y(_3313_)
);

NAND2X1 _13937_ (
    .A(areg_6_bF$buf3),
    .B(breg_13_bF$buf3),
    .Y(_3314_)
);

NAND2X1 _13938_ (
    .A(areg_7_bF$buf0),
    .B(breg_12_bF$buf1),
    .Y(_3315_)
);

NOR2X1 _13939_ (
    .A(_3314_),
    .B(_3315_),
    .Y(_3316_)
);

AND2X2 _13940_ (
    .A(_3314_),
    .B(_3315_),
    .Y(_3317_)
);

NOR2X1 _13941_ (
    .A(_3316_),
    .B(_3317_),
    .Y(_3319_)
);

XNOR2X1 _13942_ (
    .A(_3319_),
    .B(_3313_),
    .Y(_3320_)
);

AOI21X1 _13943_ (
    .A(_3061_),
    .B(_3072_),
    .C(_3063_),
    .Y(_3321_)
);

INVX1 _13944_ (
    .A(_3321_),
    .Y(_3322_)
);

NAND2X1 _13945_ (
    .A(areg_8_bF$buf4),
    .B(breg_11_bF$buf3),
    .Y(_3323_)
);

INVX2 _13946_ (
    .A(_3323_),
    .Y(_3324_)
);

AND2X2 _13947_ (
    .A(areg_9_bF$buf4),
    .B(breg_10_bF$buf5),
    .Y(_3325_)
);

AND2X2 _13948_ (
    .A(breg_9_bF$buf0),
    .B(areg_10_bF$buf0),
    .Y(_3326_)
);

NAND2X1 _13949_ (
    .A(_3325_),
    .B(_3326_),
    .Y(_3327_)
);

OAI21X1 _13950_ (
    .A(_6044__bF$buf3),
    .B(_7711__bF$buf3),
    .C(_3071_),
    .Y(_3328_)
);

NAND3X1 _13951_ (
    .A(_3324_),
    .B(_3328_),
    .C(_3327_),
    .Y(_3330_)
);

NAND2X1 _13952_ (
    .A(areg_10_bF$buf4),
    .B(breg_10_bF$buf4),
    .Y(_3331_)
);

NOR2X1 _13953_ (
    .A(_3062_),
    .B(_3331_),
    .Y(_3332_)
);

NOR2X1 _13954_ (
    .A(_3325_),
    .B(_3326_),
    .Y(_3333_)
);

OAI21X1 _13955_ (
    .A(_3333_),
    .B(_3332_),
    .C(_3323_),
    .Y(_3334_)
);

NAND3X1 _13956_ (
    .A(_3330_),
    .B(_3334_),
    .C(_3322_),
    .Y(_3335_)
);

NOR3X1 _13957_ (
    .A(_3323_),
    .B(_3332_),
    .C(_3333_),
    .Y(_3336_)
);

AOI21X1 _13958_ (
    .A(_3328_),
    .B(_3327_),
    .C(_3324_),
    .Y(_3337_)
);

OAI21X1 _13959_ (
    .A(_3336_),
    .B(_3337_),
    .C(_3321_),
    .Y(_3338_)
);

NAND3X1 _13960_ (
    .A(_3338_),
    .B(_3335_),
    .C(_3320_),
    .Y(_3339_)
);

XNOR2X1 _13961_ (
    .A(_3319_),
    .B(_3312_),
    .Y(_3340_)
);

OAI21X1 _13962_ (
    .A(_3336_),
    .B(_3337_),
    .C(_3322_),
    .Y(_3341_)
);

NAND3X1 _13963_ (
    .A(_3321_),
    .B(_3330_),
    .C(_3334_),
    .Y(_3342_)
);

NAND3X1 _13964_ (
    .A(_3341_),
    .B(_3342_),
    .C(_3340_),
    .Y(_3343_)
);

OAI21X1 _13965_ (
    .A(_3098_),
    .B(_3124_),
    .C(_3114_),
    .Y(_3344_)
);

AOI21X1 _13966_ (
    .A(_3343_),
    .B(_3339_),
    .C(_3344_),
    .Y(_3345_)
);

AOI21X1 _13967_ (
    .A(_3341_),
    .B(_3342_),
    .C(_3340_),
    .Y(_3346_)
);

AOI21X1 _13968_ (
    .A(_3338_),
    .B(_3335_),
    .C(_3320_),
    .Y(_3347_)
);

AOI21X1 _13969_ (
    .A(_3120_),
    .B(_3122_),
    .C(_3123_),
    .Y(_3348_)
);

NOR3X1 _13970_ (
    .A(_3346_),
    .B(_3348_),
    .C(_3347_),
    .Y(_3349_)
);

OAI21X1 _13971_ (
    .A(_3349_),
    .B(_3345_),
    .C(_3311_),
    .Y(_3351_)
);

INVX1 _13972_ (
    .A(_3070_),
    .Y(_3352_)
);

AOI21X1 _13973_ (
    .A(_3058_),
    .B(_3076_),
    .C(_3352_),
    .Y(_3353_)
);

OAI21X1 _13974_ (
    .A(_3347_),
    .B(_3346_),
    .C(_3348_),
    .Y(_3354_)
);

NAND3X1 _13975_ (
    .A(_3343_),
    .B(_3339_),
    .C(_3344_),
    .Y(_3355_)
);

NAND3X1 _13976_ (
    .A(_3353_),
    .B(_3355_),
    .C(_3354_),
    .Y(_3356_)
);

NAND2X1 _13977_ (
    .A(_3356_),
    .B(_3351_),
    .Y(_3357_)
);

OAI21X1 _13978_ (
    .A(_3127_),
    .B(_3186_),
    .C(_3179_),
    .Y(_3358_)
);

NAND2X1 _13979_ (
    .A(breg_7_bF$buf3),
    .B(areg_12_bF$buf0),
    .Y(_3359_)
);

OAI21X1 _13980_ (
    .A(_2845_),
    .B(_3359_),
    .C(_3106_),
    .Y(_3360_)
);

NAND2X1 _13981_ (
    .A(breg[8]),
    .B(areg_11_bF$buf0),
    .Y(_3362_)
);

INVX1 _13982_ (
    .A(_3362_),
    .Y(_3363_)
);

AND2X2 _13983_ (
    .A(breg_7_bF$buf2),
    .B(areg_12_bF$buf4),
    .Y(_3364_)
);

AND2X2 _13984_ (
    .A(breg_6_bF$buf2),
    .B(areg_13_bF$buf3),
    .Y(_3365_)
);

NAND2X1 _13985_ (
    .A(_3364_),
    .B(_3365_),
    .Y(_3366_)
);

OAI21X1 _13986_ (
    .A(_5453__bF$buf1),
    .B(_549__bF$buf1),
    .C(_3359_),
    .Y(_3367_)
);

NAND3X1 _13987_ (
    .A(_3363_),
    .B(_3367_),
    .C(_3366_),
    .Y(_3368_)
);

OAI21X1 _13988_ (
    .A(_4116__bF$buf1),
    .B(_10869__bF$buf0),
    .C(_3365_),
    .Y(_3369_)
);

OAI21X1 _13989_ (
    .A(_5453__bF$buf0),
    .B(_549__bF$buf0),
    .C(_3364_),
    .Y(_3370_)
);

NAND3X1 _13990_ (
    .A(_3362_),
    .B(_3369_),
    .C(_3370_),
    .Y(_3371_)
);

OAI21X1 _13991_ (
    .A(_3135_),
    .B(_3137_),
    .C(_3132_),
    .Y(_3373_)
);

NAND3X1 _13992_ (
    .A(_3368_),
    .B(_3371_),
    .C(_3373_),
    .Y(_3374_)
);

AOI21X1 _13993_ (
    .A(_3369_),
    .B(_3370_),
    .C(_3362_),
    .Y(_3375_)
);

AOI21X1 _13994_ (
    .A(_3367_),
    .B(_3366_),
    .C(_3363_),
    .Y(_3376_)
);

AOI21X1 _13995_ (
    .A(_3129_),
    .B(_3133_),
    .C(_3136_),
    .Y(_3377_)
);

OAI21X1 _13996_ (
    .A(_3375_),
    .B(_3376_),
    .C(_3377_),
    .Y(_3378_)
);

NAND3X1 _13997_ (
    .A(_3360_),
    .B(_3378_),
    .C(_3374_),
    .Y(_3379_)
);

INVX1 _13998_ (
    .A(_3360_),
    .Y(_3380_)
);

NOR3X1 _13999_ (
    .A(_3376_),
    .B(_3377_),
    .C(_3375_),
    .Y(_3381_)
);

AOI21X1 _14000_ (
    .A(_3368_),
    .B(_3371_),
    .C(_3373_),
    .Y(_3382_)
);

OAI21X1 _14001_ (
    .A(_3381_),
    .B(_3382_),
    .C(_3380_),
    .Y(_3384_)
);

AND2X2 _14002_ (
    .A(_3384_),
    .B(_3379_),
    .Y(_3385_)
);

OAI21X1 _14003_ (
    .A(_3174_),
    .B(_3139_),
    .C(_3167_),
    .Y(_3386_)
);

NOR2X1 _14004_ (
    .A(_4258__bF$buf0),
    .B(_2287__bF$buf1),
    .Y(_3387_)
);

INVX2 _14005_ (
    .A(_3387_),
    .Y(_3388_)
);

INVX1 _14006_ (
    .A(_3130_),
    .Y(_3389_)
);

NAND2X1 _14007_ (
    .A(breg_4_bF$buf1),
    .B(areg_16_bF$buf1),
    .Y(_3390_)
);

INVX2 _14008_ (
    .A(_3390_),
    .Y(_3391_)
);

AOI22X1 _14009_ (
    .A(breg_3_bF$buf2),
    .B(areg_16_bF$buf0),
    .C(breg_4_bF$buf0),
    .D(areg_15_bF$buf4),
    .Y(_3392_)
);

AOI21X1 _14010_ (
    .A(_3389_),
    .B(_3391_),
    .C(_3392_),
    .Y(_3393_)
);

XNOR2X1 _14011_ (
    .A(_3393_),
    .B(_3388_),
    .Y(_3395_)
);

OAI21X1 _14012_ (
    .A(_3161_),
    .B(_3141_),
    .C(_3151_),
    .Y(_3396_)
);

NAND2X1 _14013_ (
    .A(breg_2_bF$buf4),
    .B(areg_17_bF$buf1),
    .Y(_3397_)
);

INVX2 _14014_ (
    .A(_3397_),
    .Y(_3398_)
);

AND2X2 _14015_ (
    .A(breg_1_bF$buf0),
    .B(areg_18_bF$buf2),
    .Y(_3399_)
);

AND2X2 _14016_ (
    .A(breg_0_bF$buf6),
    .B(areg_19_bF$buf5),
    .Y(_3400_)
);

NAND2X1 _14017_ (
    .A(_3399_),
    .B(_3400_),
    .Y(_3401_)
);

INVX8 _14018_ (
    .A(areg_19_bF$buf4),
    .Y(_3402_)
);

NAND2X1 _14019_ (
    .A(breg_1_bF$buf6),
    .B(areg_18_bF$buf1),
    .Y(_3403_)
);

OAI21X1 _14020_ (
    .A(_2551__bF$buf3),
    .B(_3402__bF$buf3),
    .C(_3403_),
    .Y(_3404_)
);

NAND3X1 _14021_ (
    .A(_3398_),
    .B(_3404_),
    .C(_3401_),
    .Y(_3406_)
);

NAND2X1 _14022_ (
    .A(breg_0_bF$buf5),
    .B(areg_19_bF$buf3),
    .Y(_3407_)
);

NOR2X1 _14023_ (
    .A(_3403_),
    .B(_3407_),
    .Y(_3408_)
);

NOR2X1 _14024_ (
    .A(_3399_),
    .B(_3400_),
    .Y(_3409_)
);

OAI21X1 _14025_ (
    .A(_3409_),
    .B(_3408_),
    .C(_3397_),
    .Y(_3410_)
);

NAND3X1 _14026_ (
    .A(_3406_),
    .B(_3396_),
    .C(_3410_),
    .Y(_3411_)
);

AOI21X1 _14027_ (
    .A(_3150_),
    .B(_3153_),
    .C(_3160_),
    .Y(_3412_)
);

OAI21X1 _14028_ (
    .A(_3220_),
    .B(_3146__bF$buf1),
    .C(_3400_),
    .Y(_3413_)
);

OAI21X1 _14029_ (
    .A(_2551__bF$buf2),
    .B(_3402__bF$buf2),
    .C(_3399_),
    .Y(_3414_)
);

AOI21X1 _14030_ (
    .A(_3413_),
    .B(_3414_),
    .C(_3397_),
    .Y(_3415_)
);

AOI21X1 _14031_ (
    .A(_3404_),
    .B(_3401_),
    .C(_3398_),
    .Y(_3417_)
);

OAI21X1 _14032_ (
    .A(_3415_),
    .B(_3417_),
    .C(_3412_),
    .Y(_3418_)
);

NAND3X1 _14033_ (
    .A(_3418_),
    .B(_3411_),
    .C(_3395_),
    .Y(_3419_)
);

XNOR2X1 _14034_ (
    .A(_3393_),
    .B(_3387_),
    .Y(_3420_)
);

OAI21X1 _14035_ (
    .A(_3415_),
    .B(_3417_),
    .C(_3396_),
    .Y(_3421_)
);

NAND3X1 _14036_ (
    .A(_3412_),
    .B(_3406_),
    .C(_3410_),
    .Y(_3422_)
);

NAND3X1 _14037_ (
    .A(_3421_),
    .B(_3422_),
    .C(_3420_),
    .Y(_3423_)
);

NAND3X1 _14038_ (
    .A(_3423_),
    .B(_3419_),
    .C(_3386_),
    .Y(_3424_)
);

AOI21X1 _14039_ (
    .A(_3168_),
    .B(_3166_),
    .C(_3173_),
    .Y(_3425_)
);

AOI21X1 _14040_ (
    .A(_3421_),
    .B(_3422_),
    .C(_3420_),
    .Y(_3426_)
);

AOI21X1 _14041_ (
    .A(_3418_),
    .B(_3411_),
    .C(_3395_),
    .Y(_3428_)
);

OAI21X1 _14042_ (
    .A(_3428_),
    .B(_3426_),
    .C(_3425_),
    .Y(_3429_)
);

NAND3X1 _14043_ (
    .A(_3424_),
    .B(_3429_),
    .C(_3385_),
    .Y(_3430_)
);

NAND2X1 _14044_ (
    .A(_3379_),
    .B(_3384_),
    .Y(_3431_)
);

NOR3X1 _14045_ (
    .A(_3428_),
    .B(_3426_),
    .C(_3425_),
    .Y(_3432_)
);

AOI21X1 _14046_ (
    .A(_3423_),
    .B(_3419_),
    .C(_3386_),
    .Y(_3433_)
);

OAI21X1 _14047_ (
    .A(_3432_),
    .B(_3433_),
    .C(_3431_),
    .Y(_3434_)
);

NAND3X1 _14048_ (
    .A(_3430_),
    .B(_3434_),
    .C(_3358_),
    .Y(_3435_)
);

AOI21X1 _14049_ (
    .A(_3180_),
    .B(_3126_),
    .C(_3185_),
    .Y(_3436_)
);

OAI21X1 _14050_ (
    .A(_3428_),
    .B(_3426_),
    .C(_3386_),
    .Y(_3437_)
);

NAND3X1 _14051_ (
    .A(_3423_),
    .B(_3419_),
    .C(_3425_),
    .Y(_3439_)
);

AOI21X1 _14052_ (
    .A(_3439_),
    .B(_3437_),
    .C(_3431_),
    .Y(_3440_)
);

AOI21X1 _14053_ (
    .A(_3424_),
    .B(_3429_),
    .C(_3385_),
    .Y(_3441_)
);

OAI21X1 _14054_ (
    .A(_3441_),
    .B(_3440_),
    .C(_3436_),
    .Y(_3442_)
);

NAND3X1 _14055_ (
    .A(_3357_),
    .B(_3442_),
    .C(_3435_),
    .Y(_3443_)
);

NAND3X1 _14056_ (
    .A(_3355_),
    .B(_3354_),
    .C(_3311_),
    .Y(_3444_)
);

OAI21X1 _14057_ (
    .A(_3349_),
    .B(_3345_),
    .C(_3353_),
    .Y(_3445_)
);

NAND2X1 _14058_ (
    .A(_3444_),
    .B(_3445_),
    .Y(_3446_)
);

NOR3X1 _14059_ (
    .A(_3440_),
    .B(_3441_),
    .C(_3436_),
    .Y(_3447_)
);

AOI21X1 _14060_ (
    .A(_3430_),
    .B(_3434_),
    .C(_3358_),
    .Y(_3448_)
);

OAI21X1 _14061_ (
    .A(_3448_),
    .B(_3447_),
    .C(_3446_),
    .Y(_3450_)
);

NAND3X1 _14062_ (
    .A(_3443_),
    .B(_3450_),
    .C(_3310_),
    .Y(_3451_)
);

AOI21X1 _14063_ (
    .A(_3191_),
    .B(_3193_),
    .C(_3200_),
    .Y(_3452_)
);

OAI21X1 _14064_ (
    .A(_3440_),
    .B(_3441_),
    .C(_3358_),
    .Y(_3453_)
);

NAND3X1 _14065_ (
    .A(_3430_),
    .B(_3436_),
    .C(_3434_),
    .Y(_3454_)
);

AOI21X1 _14066_ (
    .A(_3454_),
    .B(_3453_),
    .C(_3446_),
    .Y(_3455_)
);

AOI21X1 _14067_ (
    .A(_3442_),
    .B(_3435_),
    .C(_3357_),
    .Y(_3456_)
);

OAI21X1 _14068_ (
    .A(_3456_),
    .B(_3455_),
    .C(_3452_),
    .Y(_3457_)
);

NAND3X1 _14069_ (
    .A(_3457_),
    .B(_3309_),
    .C(_3451_),
    .Y(_3458_)
);

NAND3X1 _14070_ (
    .A(_3249_),
    .B(_3298_),
    .C(_3303_),
    .Y(_3459_)
);

NAND3X1 _14071_ (
    .A(_3305_),
    .B(_3250_),
    .C(_3306_),
    .Y(_3461_)
);

NAND2X1 _14072_ (
    .A(_3459_),
    .B(_3461_),
    .Y(_3462_)
);

NOR3X1 _14073_ (
    .A(_3456_),
    .B(_3455_),
    .C(_3452_),
    .Y(_3463_)
);

AOI21X1 _14074_ (
    .A(_3443_),
    .B(_3450_),
    .C(_3310_),
    .Y(_3464_)
);

OAI21X1 _14075_ (
    .A(_3463_),
    .B(_3464_),
    .C(_3462_),
    .Y(_3465_)
);

NAND3X1 _14076_ (
    .A(_3458_),
    .B(_3465_),
    .C(_3248_),
    .Y(_3466_)
);

NOR3X1 _14077_ (
    .A(_3190_),
    .B(_3194_),
    .C(_3197_),
    .Y(_3467_)
);

AOI21X1 _14078_ (
    .A(_3207_),
    .B(_3210_),
    .C(_3467_),
    .Y(_3468_)
);

OAI21X1 _14079_ (
    .A(_3455_),
    .B(_3456_),
    .C(_3310_),
    .Y(_3469_)
);

NAND3X1 _14080_ (
    .A(_3443_),
    .B(_3450_),
    .C(_3452_),
    .Y(_3470_)
);

AOI21X1 _14081_ (
    .A(_3470_),
    .B(_3469_),
    .C(_3462_),
    .Y(_3472_)
);

AOI21X1 _14082_ (
    .A(_3457_),
    .B(_3451_),
    .C(_3309_),
    .Y(_3473_)
);

OAI21X1 _14083_ (
    .A(_3473_),
    .B(_3472_),
    .C(_3468_),
    .Y(_3474_)
);

NAND3X1 _14084_ (
    .A(_3246_),
    .B(_3474_),
    .C(_3466_),
    .Y(_3475_)
);

INVX2 _14085_ (
    .A(_3246_),
    .Y(_3476_)
);

OAI21X1 _14086_ (
    .A(_3473_),
    .B(_3472_),
    .C(_3248_),
    .Y(_3477_)
);

NAND3X1 _14087_ (
    .A(_3458_),
    .B(_3465_),
    .C(_3468_),
    .Y(_3478_)
);

NAND3X1 _14088_ (
    .A(_3476_),
    .B(_3477_),
    .C(_3478_),
    .Y(_3479_)
);

NAND3X1 _14089_ (
    .A(_3475_),
    .B(_3245_),
    .C(_3479_),
    .Y(_3480_)
);

NOR3X1 _14090_ (
    .A(_3204_),
    .B(_3211_),
    .C(_3214_),
    .Y(_3481_)
);

AOI21X1 _14091_ (
    .A(_2984_),
    .B(_3221_),
    .C(_3481_),
    .Y(_3483_)
);

AOI21X1 _14092_ (
    .A(_3477_),
    .B(_3478_),
    .C(_3476_),
    .Y(_3484_)
);

AOI21X1 _14093_ (
    .A(_3474_),
    .B(_3466_),
    .C(_3246_),
    .Y(_3485_)
);

OAI21X1 _14094_ (
    .A(_3484_),
    .B(_3485_),
    .C(_3483_),
    .Y(_3486_)
);

NAND3X1 _14095_ (
    .A(_3480_),
    .B(_3486_),
    .C(_3243_),
    .Y(_3487_)
);

OAI21X1 _14096_ (
    .A(_3484_),
    .B(_3485_),
    .C(_3245_),
    .Y(_3488_)
);

NAND3X1 _14097_ (
    .A(_3475_),
    .B(_3479_),
    .C(_3483_),
    .Y(_3489_)
);

NAND3X1 _14098_ (
    .A(_3230_),
    .B(_3488_),
    .C(_3489_),
    .Y(_3490_)
);

NAND3X1 _14099_ (
    .A(_3490_),
    .B(_3235_),
    .C(_3487_),
    .Y(_3491_)
);

NAND3X1 _14100_ (
    .A(_3230_),
    .B(_3232_),
    .C(_2981_),
    .Y(_3492_)
);

AOI21X1 _14101_ (
    .A(_3488_),
    .B(_3489_),
    .C(_3230_),
    .Y(_3494_)
);

NOR2X1 _14102_ (
    .A(_3222_),
    .B(_3218_),
    .Y(_3495_)
);

AOI22X1 _14103_ (
    .A(_2983_),
    .B(_3495_),
    .C(_3486_),
    .D(_3480_),
    .Y(_3496_)
);

OAI21X1 _14104_ (
    .A(_3494_),
    .B(_3496_),
    .C(_3492_),
    .Y(_3497_)
);

NAND2X1 _14105_ (
    .A(_3497_),
    .B(_3491_),
    .Y(_3498_)
);

XOR2X1 _14106_ (
    .A(_3242_),
    .B(_3498_),
    .Y(_0_[19])
);

NAND2X1 _14107_ (
    .A(_2341_),
    .B(_2532_),
    .Y(_3499_)
);

NAND3X1 _14108_ (
    .A(_2538_),
    .B(_2745_),
    .C(_3499_),
    .Y(_3500_)
);

AND2X2 _14109_ (
    .A(_2543_),
    .B(_3500_),
    .Y(_3501_)
);

AND2X2 _14110_ (
    .A(_1228_),
    .B(_1282_),
    .Y(_3502_)
);

OAI21X1 _14111_ (
    .A(_3502_),
    .B(_1391_),
    .C(_2537_),
    .Y(_3504_)
);

NAND2X1 _14112_ (
    .A(_1206_),
    .B(_1217_),
    .Y(_3505_)
);

INVX1 _14113_ (
    .A(_1369_),
    .Y(_3506_)
);

AOI22X1 _14114_ (
    .A(_11582_),
    .B(_11625_),
    .C(_3506_),
    .D(_3505_),
    .Y(_3507_)
);

NAND3X1 _14115_ (
    .A(_3507_),
    .B(_2537_),
    .C(_1271_),
    .Y(_3508_)
);

NAND3X1 _14116_ (
    .A(_3501_),
    .B(_3504_),
    .C(_3508_),
    .Y(_3509_)
);

NAND3X1 _14117_ (
    .A(_3491_),
    .B(_3497_),
    .C(_3238_),
    .Y(_3510_)
);

NAND2X1 _14118_ (
    .A(_3491_),
    .B(_3239_),
    .Y(_3511_)
);

NAND2X1 _14119_ (
    .A(_3497_),
    .B(_3511_),
    .Y(_3512_)
);

OAI21X1 _14120_ (
    .A(_3510_),
    .B(_2977_),
    .C(_3512_),
    .Y(_3513_)
);

NOR2X1 _14121_ (
    .A(_3510_),
    .B(_2979_),
    .Y(_3515_)
);

AOI21X1 _14122_ (
    .A(_3509_),
    .B(_3515_),
    .C(_3513_),
    .Y(_3516_)
);

NOR3X1 _14123_ (
    .A(_3484_),
    .B(_3485_),
    .C(_3483_),
    .Y(_3517_)
);

AOI21X1 _14124_ (
    .A(_3458_),
    .B(_3465_),
    .C(_3248_),
    .Y(_3518_)
);

OAI21X1 _14125_ (
    .A(_3518_),
    .B(_3476_),
    .C(_3466_),
    .Y(_3519_)
);

NAND2X1 _14126_ (
    .A(_3298_),
    .B(_3459_),
    .Y(_3520_)
);

INVX2 _14127_ (
    .A(_3520_),
    .Y(_3521_)
);

OAI21X1 _14128_ (
    .A(_3464_),
    .B(_3462_),
    .C(_3451_),
    .Y(_3522_)
);

NAND2X1 _14129_ (
    .A(_3286_),
    .B(_3291_),
    .Y(_3523_)
);

NOR2X1 _14130_ (
    .A(_2990_),
    .B(_3251_),
    .Y(_3524_)
);

INVX4 _14131_ (
    .A(breg_20_bF$buf4),
    .Y(_3526_)
);

NOR2X1 _14132_ (
    .A(_2376__bF$buf0),
    .B(_3526_),
    .Y(_3527_)
);

NAND2X1 _14133_ (
    .A(areg_2_bF$buf0),
    .B(breg_19_bF$buf3),
    .Y(_3528_)
);

INVX8 _14134_ (
    .A(breg_18_bF$buf3),
    .Y(_3529_)
);

OAI21X1 _14135_ (
    .A(_2519__bF$buf3),
    .B(_3529__bF$buf4),
    .C(_3251_),
    .Y(_3530_)
);

OAI21X1 _14136_ (
    .A(_3254_),
    .B(_3528_),
    .C(_3530_),
    .Y(_3531_)
);

XNOR2X1 _14137_ (
    .A(_3531_),
    .B(_3527_),
    .Y(_3532_)
);

NOR2X1 _14138_ (
    .A(_3524_),
    .B(_3532_),
    .Y(_3533_)
);

NAND2X1 _14139_ (
    .A(_3524_),
    .B(_3532_),
    .Y(_3534_)
);

INVX2 _14140_ (
    .A(_3534_),
    .Y(_3535_)
);

NOR2X1 _14141_ (
    .A(_3533_),
    .B(_3535_),
    .Y(_3537_)
);

OAI21X1 _14142_ (
    .A(_3283_),
    .B(_3281_),
    .C(_3273_),
    .Y(_3538_)
);

OAI21X1 _14143_ (
    .A(_2993_),
    .B(_3266_),
    .C(_3265_),
    .Y(_3539_)
);

NAND2X1 _14144_ (
    .A(areg_3_bF$buf4),
    .B(breg_17_bF$buf3),
    .Y(_3540_)
);

INVX1 _14145_ (
    .A(_3540_),
    .Y(_3541_)
);

NAND2X1 _14146_ (
    .A(areg_5_bF$buf2),
    .B(breg_15_bF$buf0),
    .Y(_3542_)
);

OR2X2 _14147_ (
    .A(_3266_),
    .B(_3542_),
    .Y(_3543_)
);

OAI21X1 _14148_ (
    .A(_2825__bF$buf4),
    .B(_2362__bF$buf1),
    .C(_3266_),
    .Y(_3544_)
);

NAND3X1 _14149_ (
    .A(_3541_),
    .B(_3544_),
    .C(_3543_),
    .Y(_3545_)
);

NOR2X1 _14150_ (
    .A(_3266_),
    .B(_3542_),
    .Y(_3546_)
);

AND2X2 _14151_ (
    .A(_3266_),
    .B(_3542_),
    .Y(_3548_)
);

OAI21X1 _14152_ (
    .A(_3548_),
    .B(_3546_),
    .C(_3540_),
    .Y(_3549_)
);

OAI21X1 _14153_ (
    .A(_4434__bF$buf0),
    .B(_2586__bF$buf1),
    .C(_3314_),
    .Y(_3550_)
);

AOI21X1 _14154_ (
    .A(_3312_),
    .B(_3550_),
    .C(_3316_),
    .Y(_3551_)
);

INVX2 _14155_ (
    .A(_3551_),
    .Y(_3552_)
);

NAND3X1 _14156_ (
    .A(_3549_),
    .B(_3545_),
    .C(_3552_),
    .Y(_3553_)
);

NAND2X1 _14157_ (
    .A(areg_5_bF$buf1),
    .B(breg_16_bF$buf0),
    .Y(_3554_)
);

OAI21X1 _14158_ (
    .A(_3262_),
    .B(_3554_),
    .C(_3544_),
    .Y(_3555_)
);

NOR2X1 _14159_ (
    .A(_3540_),
    .B(_3555_),
    .Y(_3556_)
);

AOI21X1 _14160_ (
    .A(_3544_),
    .B(_3543_),
    .C(_3541_),
    .Y(_3557_)
);

OAI21X1 _14161_ (
    .A(_3556_),
    .B(_3557_),
    .C(_3551_),
    .Y(_3559_)
);

NAND3X1 _14162_ (
    .A(_3539_),
    .B(_3553_),
    .C(_3559_),
    .Y(_3560_)
);

NOR2X1 _14163_ (
    .A(_2996_),
    .B(_3262_),
    .Y(_3561_)
);

NOR2X1 _14164_ (
    .A(_3561_),
    .B(_3276_),
    .Y(_3562_)
);

NAND3X1 _14165_ (
    .A(_3551_),
    .B(_3549_),
    .C(_3545_),
    .Y(_3563_)
);

OAI21X1 _14166_ (
    .A(_3556_),
    .B(_3557_),
    .C(_3552_),
    .Y(_3564_)
);

NAND3X1 _14167_ (
    .A(_3562_),
    .B(_3563_),
    .C(_3564_),
    .Y(_3565_)
);

NAND3X1 _14168_ (
    .A(_3560_),
    .B(_3565_),
    .C(_3538_),
    .Y(_3566_)
);

AOI21X1 _14169_ (
    .A(_3260_),
    .B(_3278_),
    .C(_3282_),
    .Y(_3567_)
);

AOI21X1 _14170_ (
    .A(_3563_),
    .B(_3564_),
    .C(_3562_),
    .Y(_3568_)
);

AOI21X1 _14171_ (
    .A(_3553_),
    .B(_3559_),
    .C(_3539_),
    .Y(_3570_)
);

OAI21X1 _14172_ (
    .A(_3568_),
    .B(_3570_),
    .C(_3567_),
    .Y(_3571_)
);

NAND3X1 _14173_ (
    .A(_3537_),
    .B(_3566_),
    .C(_3571_),
    .Y(_3572_)
);

OR2X2 _14174_ (
    .A(_3535_),
    .B(_3533_),
    .Y(_3573_)
);

OAI21X1 _14175_ (
    .A(_3568_),
    .B(_3570_),
    .C(_3538_),
    .Y(_3574_)
);

NAND3X1 _14176_ (
    .A(_3560_),
    .B(_3565_),
    .C(_3567_),
    .Y(_3575_)
);

NAND3X1 _14177_ (
    .A(_3574_),
    .B(_3575_),
    .C(_3573_),
    .Y(_3576_)
);

OAI21X1 _14178_ (
    .A(_3345_),
    .B(_3353_),
    .C(_3355_),
    .Y(_3577_)
);

NAND3X1 _14179_ (
    .A(_3572_),
    .B(_3577_),
    .C(_3576_),
    .Y(_3578_)
);

AOI21X1 _14180_ (
    .A(_3574_),
    .B(_3575_),
    .C(_3573_),
    .Y(_3579_)
);

AOI21X1 _14181_ (
    .A(_3566_),
    .B(_3571_),
    .C(_3537_),
    .Y(_3581_)
);

AOI21X1 _14182_ (
    .A(_3354_),
    .B(_3311_),
    .C(_3349_),
    .Y(_3582_)
);

OAI21X1 _14183_ (
    .A(_3579_),
    .B(_3581_),
    .C(_3582_),
    .Y(_3583_)
);

NAND3X1 _14184_ (
    .A(_3578_),
    .B(_3523_),
    .C(_3583_),
    .Y(_3584_)
);

INVX1 _14185_ (
    .A(_3286_),
    .Y(_3585_)
);

AOI21X1 _14186_ (
    .A(_3257_),
    .B(_3290_),
    .C(_3585_),
    .Y(_3586_)
);

NAND3X1 _14187_ (
    .A(_3572_),
    .B(_3582_),
    .C(_3576_),
    .Y(_3587_)
);

OAI21X1 _14188_ (
    .A(_3579_),
    .B(_3581_),
    .C(_3577_),
    .Y(_3588_)
);

NAND3X1 _14189_ (
    .A(_3586_),
    .B(_3587_),
    .C(_3588_),
    .Y(_3589_)
);

NAND2X1 _14190_ (
    .A(_3589_),
    .B(_3584_),
    .Y(_3590_)
);

AOI21X1 _14191_ (
    .A(_3357_),
    .B(_3442_),
    .C(_3447_),
    .Y(_3592_)
);

NAND2X1 _14192_ (
    .A(_3335_),
    .B(_3339_),
    .Y(_3593_)
);

NOR2X1 _14193_ (
    .A(_3646__bF$buf3),
    .B(_2379_),
    .Y(_3594_)
);

NAND2X1 _14194_ (
    .A(areg_7_bF$buf4),
    .B(breg_13_bF$buf2),
    .Y(_3595_)
);

NAND2X1 _14195_ (
    .A(areg_8_bF$buf3),
    .B(breg_12_bF$buf0),
    .Y(_3596_)
);

XOR2X1 _14196_ (
    .A(_3595_),
    .B(_3596_),
    .Y(_3597_)
);

XNOR2X1 _14197_ (
    .A(_3597_),
    .B(_3594_),
    .Y(_3598_)
);

AOI21X1 _14198_ (
    .A(_3324_),
    .B(_3328_),
    .C(_3332_),
    .Y(_3599_)
);

INVX1 _14199_ (
    .A(_3599_),
    .Y(_3600_)
);

NAND2X1 _14200_ (
    .A(areg_9_bF$buf3),
    .B(breg_11_bF$buf2),
    .Y(_3601_)
);

AND2X2 _14201_ (
    .A(breg_9_bF$buf5),
    .B(areg_11_bF$buf4),
    .Y(_3602_)
);

OAI21X1 _14202_ (
    .A(_7711__bF$buf2),
    .B(_7217__bF$buf2),
    .C(_3602_),
    .Y(_3603_)
);

AND2X2 _14203_ (
    .A(areg_10_bF$buf3),
    .B(breg_10_bF$buf3),
    .Y(_3604_)
);

OAI21X1 _14204_ (
    .A(_6044__bF$buf2),
    .B(_9104__bF$buf1),
    .C(_3604_),
    .Y(_3605_)
);

AOI21X1 _14205_ (
    .A(_3603_),
    .B(_3605_),
    .C(_3601_),
    .Y(_3606_)
);

INVX2 _14206_ (
    .A(_3601_),
    .Y(_3607_)
);

NAND2X1 _14207_ (
    .A(_3604_),
    .B(_3602_),
    .Y(_3608_)
);

OAI21X1 _14208_ (
    .A(_6044__bF$buf1),
    .B(_9104__bF$buf0),
    .C(_3331_),
    .Y(_3609_)
);

AOI21X1 _14209_ (
    .A(_3609_),
    .B(_3608_),
    .C(_3607_),
    .Y(_3610_)
);

OAI21X1 _14210_ (
    .A(_3606_),
    .B(_3610_),
    .C(_3600_),
    .Y(_3611_)
);

NAND3X1 _14211_ (
    .A(_3607_),
    .B(_3609_),
    .C(_3608_),
    .Y(_3614_)
);

AND2X2 _14212_ (
    .A(_3604_),
    .B(_3602_),
    .Y(_3615_)
);

NOR2X1 _14213_ (
    .A(_3604_),
    .B(_3602_),
    .Y(_3616_)
);

OAI21X1 _14214_ (
    .A(_3615_),
    .B(_3616_),
    .C(_3601_),
    .Y(_3617_)
);

NAND3X1 _14215_ (
    .A(_3599_),
    .B(_3614_),
    .C(_3617_),
    .Y(_3618_)
);

AOI21X1 _14216_ (
    .A(_3618_),
    .B(_3611_),
    .C(_3598_),
    .Y(_3619_)
);

INVX1 _14217_ (
    .A(_3594_),
    .Y(_3620_)
);

XNOR2X1 _14218_ (
    .A(_3597_),
    .B(_3620_),
    .Y(_3621_)
);

NAND3X1 _14219_ (
    .A(_3614_),
    .B(_3617_),
    .C(_3600_),
    .Y(_3622_)
);

OAI21X1 _14220_ (
    .A(_3606_),
    .B(_3610_),
    .C(_3599_),
    .Y(_3623_)
);

AOI21X1 _14221_ (
    .A(_3623_),
    .B(_3622_),
    .C(_3621_),
    .Y(_3625_)
);

AOI21X1 _14222_ (
    .A(_3378_),
    .B(_3360_),
    .C(_3381_),
    .Y(_3626_)
);

OAI21X1 _14223_ (
    .A(_3625_),
    .B(_3619_),
    .C(_3626_),
    .Y(_3627_)
);

NAND3X1 _14224_ (
    .A(_3621_),
    .B(_3623_),
    .C(_3622_),
    .Y(_3628_)
);

NAND3X1 _14225_ (
    .A(_3618_),
    .B(_3611_),
    .C(_3598_),
    .Y(_3629_)
);

OAI21X1 _14226_ (
    .A(_3380_),
    .B(_3382_),
    .C(_3374_),
    .Y(_3630_)
);

NAND3X1 _14227_ (
    .A(_3629_),
    .B(_3628_),
    .C(_3630_),
    .Y(_3631_)
);

NAND3X1 _14228_ (
    .A(_3593_),
    .B(_3631_),
    .C(_3627_),
    .Y(_3632_)
);

AND2X2 _14229_ (
    .A(_3339_),
    .B(_3335_),
    .Y(_3633_)
);

AOI21X1 _14230_ (
    .A(_3629_),
    .B(_3628_),
    .C(_3630_),
    .Y(_3634_)
);

NOR3X1 _14231_ (
    .A(_3619_),
    .B(_3626_),
    .C(_3625_),
    .Y(_3636_)
);

OAI21X1 _14232_ (
    .A(_3636_),
    .B(_3634_),
    .C(_3633_),
    .Y(_3637_)
);

NAND2X1 _14233_ (
    .A(_3632_),
    .B(_3637_),
    .Y(_3638_)
);

OAI21X1 _14234_ (
    .A(_3433_),
    .B(_3431_),
    .C(_3424_),
    .Y(_3639_)
);

INVX1 _14235_ (
    .A(_3365_),
    .Y(_3640_)
);

OAI21X1 _14236_ (
    .A(_3359_),
    .B(_3640_),
    .C(_3368_),
    .Y(_3641_)
);

NOR2X1 _14237_ (
    .A(_5420__bF$buf2),
    .B(_10869__bF$buf3),
    .Y(_3642_)
);

AND2X2 _14238_ (
    .A(breg_7_bF$buf1),
    .B(areg_13_bF$buf2),
    .Y(_3643_)
);

AND2X2 _14239_ (
    .A(breg_6_bF$buf1),
    .B(areg_14_bF$buf3),
    .Y(_3644_)
);

NAND2X1 _14240_ (
    .A(_3643_),
    .B(_3644_),
    .Y(_3645_)
);

OAI22X1 _14241_ (
    .A(_5453__bF$buf5),
    .B(_2287__bF$buf0),
    .C(_4116__bF$buf0),
    .D(_549__bF$buf4),
    .Y(_3647_)
);

NAND3X1 _14242_ (
    .A(_3642_),
    .B(_3647_),
    .C(_3645_),
    .Y(_3648_)
);

INVX1 _14243_ (
    .A(_3642_),
    .Y(_3649_)
);

OAI21X1 _14244_ (
    .A(_4116__bF$buf4),
    .B(_549__bF$buf3),
    .C(_3644_),
    .Y(_3650_)
);

OAI21X1 _14245_ (
    .A(_5453__bF$buf4),
    .B(_2287__bF$buf3),
    .C(_3643_),
    .Y(_3651_)
);

NAND3X1 _14246_ (
    .A(_3650_),
    .B(_3651_),
    .C(_3649_),
    .Y(_3652_)
);

OAI22X1 _14247_ (
    .A(_3130_),
    .B(_3390_),
    .C(_3388_),
    .D(_3392_),
    .Y(_3653_)
);

NAND3X1 _14248_ (
    .A(_3648_),
    .B(_3652_),
    .C(_3653_),
    .Y(_3654_)
);

AOI21X1 _14249_ (
    .A(_3650_),
    .B(_3651_),
    .C(_3649_),
    .Y(_3655_)
);

AOI21X1 _14250_ (
    .A(_3647_),
    .B(_3645_),
    .C(_3642_),
    .Y(_3656_)
);

INVX1 _14251_ (
    .A(_3392_),
    .Y(_3658_)
);

AOI22X1 _14252_ (
    .A(_3389_),
    .B(_3391_),
    .C(_3658_),
    .D(_3387_),
    .Y(_3659_)
);

OAI21X1 _14253_ (
    .A(_3655_),
    .B(_3656_),
    .C(_3659_),
    .Y(_3660_)
);

NAND3X1 _14254_ (
    .A(_3641_),
    .B(_3660_),
    .C(_3654_),
    .Y(_3661_)
);

INVX2 _14255_ (
    .A(_3641_),
    .Y(_3662_)
);

NOR3X1 _14256_ (
    .A(_3656_),
    .B(_3659_),
    .C(_3655_),
    .Y(_3663_)
);

AOI21X1 _14257_ (
    .A(_3648_),
    .B(_3652_),
    .C(_3653_),
    .Y(_3664_)
);

OAI21X1 _14258_ (
    .A(_3663_),
    .B(_3664_),
    .C(_3662_),
    .Y(_3665_)
);

NAND2X1 _14259_ (
    .A(_3661_),
    .B(_3665_),
    .Y(_3666_)
);

AOI21X1 _14260_ (
    .A(_3406_),
    .B(_3410_),
    .C(_3396_),
    .Y(_3667_)
);

OAI21X1 _14261_ (
    .A(_3667_),
    .B(_3420_),
    .C(_3411_),
    .Y(_3669_)
);

NOR2X1 _14262_ (
    .A(_4258__bF$buf3),
    .B(_2465__bF$buf2),
    .Y(_3670_)
);

AND2X2 _14263_ (
    .A(breg_3_bF$buf1),
    .B(areg_16_bF$buf5),
    .Y(_3671_)
);

NAND2X1 _14264_ (
    .A(breg_4_bF$buf5),
    .B(areg_17_bF$buf0),
    .Y(_3672_)
);

INVX2 _14265_ (
    .A(_3672_),
    .Y(_3673_)
);

AOI22X1 _14266_ (
    .A(breg_3_bF$buf0),
    .B(areg_17_bF$buf5),
    .C(breg_4_bF$buf4),
    .D(areg_16_bF$buf4),
    .Y(_3674_)
);

AOI21X1 _14267_ (
    .A(_3671_),
    .B(_3673_),
    .C(_3674_),
    .Y(_3675_)
);

XNOR2X1 _14268_ (
    .A(_3675_),
    .B(_3670_),
    .Y(_3676_)
);

OAI21X1 _14269_ (
    .A(_3409_),
    .B(_3397_),
    .C(_3401_),
    .Y(_3677_)
);

NAND2X1 _14270_ (
    .A(breg_2_bF$buf3),
    .B(areg_18_bF$buf0),
    .Y(_3678_)
);

NAND2X1 _14271_ (
    .A(breg_1_bF$buf5),
    .B(areg_20_bF$buf4),
    .Y(_3680_)
);

NOR2X1 _14272_ (
    .A(_3407_),
    .B(_3680_),
    .Y(_3681_)
);

AOI22X1 _14273_ (
    .A(breg_0_bF$buf4),
    .B(areg_20_bF$buf3),
    .C(breg_1_bF$buf4),
    .D(areg_19_bF$buf2),
    .Y(_3682_)
);

NOR3X1 _14274_ (
    .A(_3678_),
    .B(_3682_),
    .C(_3681_),
    .Y(_3683_)
);

INVX2 _14275_ (
    .A(_3678_),
    .Y(_3684_)
);

AND2X2 _14276_ (
    .A(breg_1_bF$buf3),
    .B(areg_20_bF$buf2),
    .Y(_3685_)
);

NAND2X1 _14277_ (
    .A(_3400_),
    .B(_3685_),
    .Y(_3686_)
);

INVX2 _14278_ (
    .A(_3682_),
    .Y(_3687_)
);

AOI21X1 _14279_ (
    .A(_3687_),
    .B(_3686_),
    .C(_3684_),
    .Y(_3688_)
);

OAI21X1 _14280_ (
    .A(_3688_),
    .B(_3683_),
    .C(_3677_),
    .Y(_3689_)
);

AOI21X1 _14281_ (
    .A(_3398_),
    .B(_3404_),
    .C(_3408_),
    .Y(_3691_)
);

NAND3X1 _14282_ (
    .A(_3684_),
    .B(_3687_),
    .C(_3686_),
    .Y(_3692_)
);

OAI21X1 _14283_ (
    .A(_3681_),
    .B(_3682_),
    .C(_3678_),
    .Y(_3693_)
);

NAND3X1 _14284_ (
    .A(_3691_),
    .B(_3693_),
    .C(_3692_),
    .Y(_3694_)
);

AOI21X1 _14285_ (
    .A(_3694_),
    .B(_3689_),
    .C(_3676_),
    .Y(_3695_)
);

XOR2X1 _14286_ (
    .A(_3675_),
    .B(_3670_),
    .Y(_3696_)
);

NAND3X1 _14287_ (
    .A(_3693_),
    .B(_3692_),
    .C(_3677_),
    .Y(_3697_)
);

OAI21X1 _14288_ (
    .A(_3688_),
    .B(_3683_),
    .C(_3691_),
    .Y(_3698_)
);

AOI21X1 _14289_ (
    .A(_3698_),
    .B(_3697_),
    .C(_3696_),
    .Y(_3699_)
);

OAI21X1 _14290_ (
    .A(_3699_),
    .B(_3695_),
    .C(_3669_),
    .Y(_3700_)
);

NOR3X1 _14291_ (
    .A(_3417_),
    .B(_3412_),
    .C(_3415_),
    .Y(_3702_)
);

AOI21X1 _14292_ (
    .A(_3418_),
    .B(_3395_),
    .C(_3702_),
    .Y(_3703_)
);

NAND3X1 _14293_ (
    .A(_3698_),
    .B(_3697_),
    .C(_3696_),
    .Y(_3704_)
);

NAND3X1 _14294_ (
    .A(_3694_),
    .B(_3689_),
    .C(_3676_),
    .Y(_3705_)
);

NAND3X1 _14295_ (
    .A(_3704_),
    .B(_3705_),
    .C(_3703_),
    .Y(_3706_)
);

AOI21X1 _14296_ (
    .A(_3706_),
    .B(_3700_),
    .C(_3666_),
    .Y(_3707_)
);

NAND3X1 _14297_ (
    .A(_3660_),
    .B(_3654_),
    .C(_3662_),
    .Y(_3708_)
);

OAI21X1 _14298_ (
    .A(_3663_),
    .B(_3664_),
    .C(_3641_),
    .Y(_3709_)
);

NAND2X1 _14299_ (
    .A(_3708_),
    .B(_3709_),
    .Y(_3710_)
);

NAND3X1 _14300_ (
    .A(_3704_),
    .B(_3705_),
    .C(_3669_),
    .Y(_3711_)
);

OAI21X1 _14301_ (
    .A(_3699_),
    .B(_3695_),
    .C(_3703_),
    .Y(_3713_)
);

AOI21X1 _14302_ (
    .A(_3711_),
    .B(_3713_),
    .C(_3710_),
    .Y(_3714_)
);

OAI21X1 _14303_ (
    .A(_3714_),
    .B(_3707_),
    .C(_3639_),
    .Y(_3715_)
);

AOI21X1 _14304_ (
    .A(_3429_),
    .B(_3385_),
    .C(_3432_),
    .Y(_3716_)
);

NAND3X1 _14305_ (
    .A(_3711_),
    .B(_3710_),
    .C(_3713_),
    .Y(_3717_)
);

NAND3X1 _14306_ (
    .A(_3706_),
    .B(_3666_),
    .C(_3700_),
    .Y(_3718_)
);

NAND3X1 _14307_ (
    .A(_3717_),
    .B(_3718_),
    .C(_3716_),
    .Y(_3719_)
);

AOI21X1 _14308_ (
    .A(_3715_),
    .B(_3719_),
    .C(_3638_),
    .Y(_3720_)
);

OAI21X1 _14309_ (
    .A(_3636_),
    .B(_3634_),
    .C(_3593_),
    .Y(_3721_)
);

NAND3X1 _14310_ (
    .A(_3631_),
    .B(_3633_),
    .C(_3627_),
    .Y(_3722_)
);

NAND2X1 _14311_ (
    .A(_3722_),
    .B(_3721_),
    .Y(_3724_)
);

NAND3X1 _14312_ (
    .A(_3639_),
    .B(_3717_),
    .C(_3718_),
    .Y(_3725_)
);

OAI21X1 _14313_ (
    .A(_3714_),
    .B(_3707_),
    .C(_3716_),
    .Y(_3726_)
);

AOI21X1 _14314_ (
    .A(_3725_),
    .B(_3726_),
    .C(_3724_),
    .Y(_3727_)
);

NOR3X1 _14315_ (
    .A(_3720_),
    .B(_3727_),
    .C(_3592_),
    .Y(_3728_)
);

OAI21X1 _14316_ (
    .A(_3448_),
    .B(_3446_),
    .C(_3435_),
    .Y(_3729_)
);

NAND3X1 _14317_ (
    .A(_3725_),
    .B(_3726_),
    .C(_3724_),
    .Y(_3730_)
);

NOR3X1 _14318_ (
    .A(_3707_),
    .B(_3714_),
    .C(_3716_),
    .Y(_3731_)
);

AOI21X1 _14319_ (
    .A(_3718_),
    .B(_3717_),
    .C(_3639_),
    .Y(_3732_)
);

OAI21X1 _14320_ (
    .A(_3731_),
    .B(_3732_),
    .C(_3638_),
    .Y(_3733_)
);

AOI21X1 _14321_ (
    .A(_3730_),
    .B(_3733_),
    .C(_3729_),
    .Y(_3735_)
);

NOR3X1 _14322_ (
    .A(_3728_),
    .B(_3590_),
    .C(_3735_),
    .Y(_3736_)
);

NAND3X1 _14323_ (
    .A(_3586_),
    .B(_3578_),
    .C(_3583_),
    .Y(_3737_)
);

NAND3X1 _14324_ (
    .A(_3587_),
    .B(_3523_),
    .C(_3588_),
    .Y(_3738_)
);

NAND2X1 _14325_ (
    .A(_3737_),
    .B(_3738_),
    .Y(_3739_)
);

NAND3X1 _14326_ (
    .A(_3730_),
    .B(_3733_),
    .C(_3729_),
    .Y(_3740_)
);

OAI21X1 _14327_ (
    .A(_3720_),
    .B(_3727_),
    .C(_3592_),
    .Y(_3741_)
);

AOI21X1 _14328_ (
    .A(_3741_),
    .B(_3740_),
    .C(_3739_),
    .Y(_3742_)
);

OAI21X1 _14329_ (
    .A(_3736_),
    .B(_3742_),
    .C(_3522_),
    .Y(_3743_)
);

AOI21X1 _14330_ (
    .A(_3457_),
    .B(_3309_),
    .C(_3463_),
    .Y(_3744_)
);

NAND3X1 _14331_ (
    .A(_3741_),
    .B(_3739_),
    .C(_3740_),
    .Y(_3746_)
);

OAI21X1 _14332_ (
    .A(_3735_),
    .B(_3728_),
    .C(_3590_),
    .Y(_3747_)
);

NAND3X1 _14333_ (
    .A(_3746_),
    .B(_3747_),
    .C(_3744_),
    .Y(_3748_)
);

AOI21X1 _14334_ (
    .A(_3743_),
    .B(_3748_),
    .C(_3521_),
    .Y(_3749_)
);

NAND3X1 _14335_ (
    .A(_3746_),
    .B(_3747_),
    .C(_3522_),
    .Y(_3750_)
);

OAI21X1 _14336_ (
    .A(_3736_),
    .B(_3742_),
    .C(_3744_),
    .Y(_3751_)
);

AOI21X1 _14337_ (
    .A(_3751_),
    .B(_3750_),
    .C(_3520_),
    .Y(_3752_)
);

OAI21X1 _14338_ (
    .A(_3752_),
    .B(_3749_),
    .C(_3519_),
    .Y(_3753_)
);

NOR3X1 _14339_ (
    .A(_3473_),
    .B(_3472_),
    .C(_3468_),
    .Y(_3754_)
);

AOI21X1 _14340_ (
    .A(_3246_),
    .B(_3474_),
    .C(_3754_),
    .Y(_3755_)
);

NAND3X1 _14341_ (
    .A(_3520_),
    .B(_3751_),
    .C(_3750_),
    .Y(_3757_)
);

NOR3X1 _14342_ (
    .A(_3736_),
    .B(_3742_),
    .C(_3744_),
    .Y(_3758_)
);

AOI21X1 _14343_ (
    .A(_3746_),
    .B(_3747_),
    .C(_3522_),
    .Y(_3759_)
);

OAI21X1 _14344_ (
    .A(_3758_),
    .B(_3759_),
    .C(_3521_),
    .Y(_3760_)
);

NAND3X1 _14345_ (
    .A(_3757_),
    .B(_3760_),
    .C(_3755_),
    .Y(_3761_)
);

AOI21X1 _14346_ (
    .A(_3753_),
    .B(_3761_),
    .C(_3517_),
    .Y(_3762_)
);

NAND3X1 _14347_ (
    .A(_3757_),
    .B(_3519_),
    .C(_3760_),
    .Y(_3763_)
);

OAI21X1 _14348_ (
    .A(_3752_),
    .B(_3749_),
    .C(_3755_),
    .Y(_3764_)
);

AOI21X1 _14349_ (
    .A(_3764_),
    .B(_3763_),
    .C(_3480_),
    .Y(_3765_)
);

OAI21X1 _14350_ (
    .A(_3762_),
    .B(_3765_),
    .C(_3487_),
    .Y(_3766_)
);

AOI21X1 _14351_ (
    .A(_3753_),
    .B(_3761_),
    .C(_3480_),
    .Y(_3767_)
);

AOI21X1 _14352_ (
    .A(_3763_),
    .B(_3764_),
    .C(_3517_),
    .Y(_3768_)
);

OAI21X1 _14353_ (
    .A(_3768_),
    .B(_3767_),
    .C(_3494_),
    .Y(_3769_)
);

NAND2X1 _14354_ (
    .A(_3766_),
    .B(_3769_),
    .Y(_3770_)
);

XNOR2X1 _14355_ (
    .A(_3516_),
    .B(_3770_),
    .Y(_0_[20])
);

OAI21X1 _14356_ (
    .A(_3762_),
    .B(_3765_),
    .C(_3494_),
    .Y(_3771_)
);

INVX1 _14357_ (
    .A(_3770_),
    .Y(_3772_)
);

OAI21X1 _14358_ (
    .A(_3516_),
    .B(_3772_),
    .C(_3771_),
    .Y(_3773_)
);

NOR2X1 _14359_ (
    .A(_3749_),
    .B(_3752_),
    .Y(_3774_)
);

OAI21X1 _14360_ (
    .A(_3759_),
    .B(_3521_),
    .C(_3750_),
    .Y(_3775_)
);

NAND2X1 _14361_ (
    .A(_3578_),
    .B(_3584_),
    .Y(_3777_)
);

XNOR2X1 _14362_ (
    .A(_3777_),
    .B(_3535_),
    .Y(_3778_)
);

AOI21X1 _14363_ (
    .A(_3739_),
    .B(_3741_),
    .C(_3728_),
    .Y(_3779_)
);

NAND2X1 _14364_ (
    .A(_3566_),
    .B(_3572_),
    .Y(_3780_)
);

INVX8 _14365_ (
    .A(breg_21_bF$buf4),
    .Y(_3781_)
);

NOR2X1 _14366_ (
    .A(_2376__bF$buf3),
    .B(_3781__bF$buf3),
    .Y(_3782_)
);

INVX2 _14367_ (
    .A(_3782_),
    .Y(_3783_)
);

NOR2X1 _14368_ (
    .A(_3254_),
    .B(_3528_),
    .Y(_3784_)
);

AOI21X1 _14369_ (
    .A(_3527_),
    .B(_3530_),
    .C(_3784_),
    .Y(_3785_)
);

INVX1 _14370_ (
    .A(_3785_),
    .Y(_3786_)
);

NAND2X1 _14371_ (
    .A(areg_1_bF$buf0),
    .B(breg_20_bF$buf3),
    .Y(_3789_)
);

NAND2X1 _14372_ (
    .A(areg_3_bF$buf3),
    .B(breg_18_bF$buf2),
    .Y(_3790_)
);

NOR2X1 _14373_ (
    .A(_3528_),
    .B(_3790_),
    .Y(_3791_)
);

AND2X2 _14374_ (
    .A(_3528_),
    .B(_3790_),
    .Y(_3792_)
);

OAI21X1 _14375_ (
    .A(_3792_),
    .B(_3791_),
    .C(_3789_),
    .Y(_3793_)
);

INVX1 _14376_ (
    .A(_3789_),
    .Y(_3794_)
);

OR2X2 _14377_ (
    .A(_3528_),
    .B(_3790_),
    .Y(_3795_)
);

OAI21X1 _14378_ (
    .A(_2519__bF$buf2),
    .B(_3253__bF$buf2),
    .C(_3790_),
    .Y(_3796_)
);

NAND3X1 _14379_ (
    .A(_3794_),
    .B(_3796_),
    .C(_3795_),
    .Y(_3797_)
);

AOI21X1 _14380_ (
    .A(_3793_),
    .B(_3797_),
    .C(_3786_),
    .Y(_3798_)
);

NAND2X1 _14381_ (
    .A(_3793_),
    .B(_3797_),
    .Y(_3800_)
);

NOR2X1 _14382_ (
    .A(_3785_),
    .B(_3800_),
    .Y(_3801_)
);

OAI21X1 _14383_ (
    .A(_3801_),
    .B(_3798_),
    .C(_3783_),
    .Y(_3802_)
);

NAND2X1 _14384_ (
    .A(_3785_),
    .B(_3800_),
    .Y(_3803_)
);

NAND3X1 _14385_ (
    .A(_3793_),
    .B(_3797_),
    .C(_3786_),
    .Y(_3804_)
);

NAND3X1 _14386_ (
    .A(_3782_),
    .B(_3804_),
    .C(_3803_),
    .Y(_3805_)
);

AND2X2 _14387_ (
    .A(_3802_),
    .B(_3805_),
    .Y(_3806_)
);

AOI21X1 _14388_ (
    .A(_3549_),
    .B(_3545_),
    .C(_3552_),
    .Y(_3807_)
);

OAI21X1 _14389_ (
    .A(_3562_),
    .B(_3807_),
    .C(_3553_),
    .Y(_3808_)
);

OAI21X1 _14390_ (
    .A(_3548_),
    .B(_3540_),
    .C(_3543_),
    .Y(_3809_)
);

NOR2X1 _14391_ (
    .A(_2562__bF$buf3),
    .B(_2763_),
    .Y(_3811_)
);

AND2X2 _14392_ (
    .A(areg_5_bF$buf0),
    .B(breg_16_bF$buf5),
    .Y(_3812_)
);

AND2X2 _14393_ (
    .A(areg_6_bF$buf2),
    .B(breg_15_bF$buf5),
    .Y(_3813_)
);

NAND2X1 _14394_ (
    .A(_3812_),
    .B(_3813_),
    .Y(_3814_)
);

OAI21X1 _14395_ (
    .A(_3646__bF$buf2),
    .B(_2362__bF$buf0),
    .C(_3554_),
    .Y(_3815_)
);

NAND3X1 _14396_ (
    .A(_3811_),
    .B(_3815_),
    .C(_3814_),
    .Y(_3816_)
);

NAND2X1 _14397_ (
    .A(areg_6_bF$buf1),
    .B(breg_16_bF$buf4),
    .Y(_3817_)
);

OAI21X1 _14398_ (
    .A(_3542_),
    .B(_3817_),
    .C(_3815_),
    .Y(_3818_)
);

OAI21X1 _14399_ (
    .A(_2562__bF$buf2),
    .B(_2763_),
    .C(_3818_),
    .Y(_3819_)
);

NOR2X1 _14400_ (
    .A(_3595_),
    .B(_3596_),
    .Y(_3820_)
);

OAI21X1 _14401_ (
    .A(_5190__bF$buf2),
    .B(_2586__bF$buf0),
    .C(_3595_),
    .Y(_3822_)
);

AOI21X1 _14402_ (
    .A(_3594_),
    .B(_3822_),
    .C(_3820_),
    .Y(_3823_)
);

INVX2 _14403_ (
    .A(_3823_),
    .Y(_3824_)
);

NAND3X1 _14404_ (
    .A(_3816_),
    .B(_3819_),
    .C(_3824_),
    .Y(_3825_)
);

INVX1 _14405_ (
    .A(_3811_),
    .Y(_3826_)
);

OAI21X1 _14406_ (
    .A(_2825__bF$buf3),
    .B(_2560__bF$buf3),
    .C(_3813_),
    .Y(_3827_)
);

OAI21X1 _14407_ (
    .A(_3646__bF$buf1),
    .B(_2362__bF$buf5),
    .C(_3812_),
    .Y(_3828_)
);

AOI21X1 _14408_ (
    .A(_3827_),
    .B(_3828_),
    .C(_3826_),
    .Y(_3829_)
);

AOI21X1 _14409_ (
    .A(_3815_),
    .B(_3814_),
    .C(_3811_),
    .Y(_3830_)
);

OAI21X1 _14410_ (
    .A(_3829_),
    .B(_3830_),
    .C(_3823_),
    .Y(_3831_)
);

NAND3X1 _14411_ (
    .A(_3809_),
    .B(_3831_),
    .C(_3825_),
    .Y(_3833_)
);

INVX2 _14412_ (
    .A(_3809_),
    .Y(_3834_)
);

NOR3X1 _14413_ (
    .A(_3830_),
    .B(_3823_),
    .C(_3829_),
    .Y(_3835_)
);

AOI21X1 _14414_ (
    .A(_3816_),
    .B(_3819_),
    .C(_3824_),
    .Y(_3836_)
);

OAI21X1 _14415_ (
    .A(_3836_),
    .B(_3835_),
    .C(_3834_),
    .Y(_3837_)
);

NAND3X1 _14416_ (
    .A(_3833_),
    .B(_3808_),
    .C(_3837_),
    .Y(_3838_)
);

NAND2X1 _14417_ (
    .A(_3549_),
    .B(_3545_),
    .Y(_3839_)
);

NOR2X1 _14418_ (
    .A(_3551_),
    .B(_3839_),
    .Y(_3840_)
);

AOI21X1 _14419_ (
    .A(_3539_),
    .B(_3559_),
    .C(_3840_),
    .Y(_3841_)
);

NAND3X1 _14420_ (
    .A(_3816_),
    .B(_3823_),
    .C(_3819_),
    .Y(_3842_)
);

OAI21X1 _14421_ (
    .A(_3829_),
    .B(_3830_),
    .C(_3824_),
    .Y(_3844_)
);

AOI21X1 _14422_ (
    .A(_3844_),
    .B(_3842_),
    .C(_3834_),
    .Y(_3845_)
);

AOI21X1 _14423_ (
    .A(_3831_),
    .B(_3825_),
    .C(_3809_),
    .Y(_3846_)
);

OAI21X1 _14424_ (
    .A(_3846_),
    .B(_3845_),
    .C(_3841_),
    .Y(_3847_)
);

NAND3X1 _14425_ (
    .A(_3838_),
    .B(_3847_),
    .C(_3806_),
    .Y(_3848_)
);

NAND2X1 _14426_ (
    .A(_3805_),
    .B(_3802_),
    .Y(_3849_)
);

OAI21X1 _14427_ (
    .A(_3846_),
    .B(_3845_),
    .C(_3808_),
    .Y(_3850_)
);

NAND3X1 _14428_ (
    .A(_3833_),
    .B(_3837_),
    .C(_3841_),
    .Y(_3851_)
);

NAND3X1 _14429_ (
    .A(_3850_),
    .B(_3849_),
    .C(_3851_),
    .Y(_3852_)
);

OAI21X1 _14430_ (
    .A(_3633_),
    .B(_3634_),
    .C(_3631_),
    .Y(_3853_)
);

NAND3X1 _14431_ (
    .A(_3852_),
    .B(_3853_),
    .C(_3848_),
    .Y(_3855_)
);

AOI21X1 _14432_ (
    .A(_3850_),
    .B(_3851_),
    .C(_3849_),
    .Y(_3856_)
);

AOI22X1 _14433_ (
    .A(_3802_),
    .B(_3805_),
    .C(_3847_),
    .D(_3838_),
    .Y(_3857_)
);

AOI21X1 _14434_ (
    .A(_3593_),
    .B(_3627_),
    .C(_3636_),
    .Y(_3858_)
);

OAI21X1 _14435_ (
    .A(_3856_),
    .B(_3857_),
    .C(_3858_),
    .Y(_3859_)
);

NAND3X1 _14436_ (
    .A(_3780_),
    .B(_3859_),
    .C(_3855_),
    .Y(_3860_)
);

AND2X2 _14437_ (
    .A(_3572_),
    .B(_3566_),
    .Y(_3861_)
);

NAND3X1 _14438_ (
    .A(_3852_),
    .B(_3858_),
    .C(_3848_),
    .Y(_3862_)
);

OAI21X1 _14439_ (
    .A(_3856_),
    .B(_3857_),
    .C(_3853_),
    .Y(_3863_)
);

NAND3X1 _14440_ (
    .A(_3861_),
    .B(_3863_),
    .C(_3862_),
    .Y(_3864_)
);

NAND2X1 _14441_ (
    .A(_3860_),
    .B(_3864_),
    .Y(_3866_)
);

OAI21X1 _14442_ (
    .A(_3638_),
    .B(_3732_),
    .C(_3725_),
    .Y(_3867_)
);

NAND2X1 _14443_ (
    .A(_3622_),
    .B(_3628_),
    .Y(_3868_)
);

NOR2X1 _14444_ (
    .A(_4434__bF$buf3),
    .B(_2379_),
    .Y(_3869_)
);

NAND2X1 _14445_ (
    .A(areg_8_bF$buf2),
    .B(breg_13_bF$buf1),
    .Y(_3870_)
);

NAND2X1 _14446_ (
    .A(areg_9_bF$buf2),
    .B(breg_12_bF$buf4),
    .Y(_3871_)
);

XOR2X1 _14447_ (
    .A(_3870_),
    .B(_3871_),
    .Y(_3872_)
);

XNOR2X1 _14448_ (
    .A(_3872_),
    .B(_3869_),
    .Y(_3873_)
);

OAI21X1 _14449_ (
    .A(_3616_),
    .B(_3601_),
    .C(_3608_),
    .Y(_3874_)
);

NAND2X1 _14450_ (
    .A(areg_10_bF$buf2),
    .B(breg_11_bF$buf1),
    .Y(_3875_)
);

AND2X2 _14451_ (
    .A(breg_9_bF$buf4),
    .B(areg_12_bF$buf3),
    .Y(_3877_)
);

OAI21X1 _14452_ (
    .A(_7217__bF$buf1),
    .B(_9104__bF$buf3),
    .C(_3877_),
    .Y(_3878_)
);

AND2X2 _14453_ (
    .A(breg_10_bF$buf2),
    .B(areg_11_bF$buf3),
    .Y(_3879_)
);

OAI21X1 _14454_ (
    .A(_6044__bF$buf0),
    .B(_10869__bF$buf2),
    .C(_3879_),
    .Y(_3880_)
);

AOI21X1 _14455_ (
    .A(_3878_),
    .B(_3880_),
    .C(_3875_),
    .Y(_3881_)
);

INVX2 _14456_ (
    .A(_3875_),
    .Y(_3882_)
);

NAND2X1 _14457_ (
    .A(_3879_),
    .B(_3877_),
    .Y(_3883_)
);

OAI22X1 _14458_ (
    .A(_6044__bF$buf5),
    .B(_10869__bF$buf1),
    .C(_7217__bF$buf0),
    .D(_9104__bF$buf2),
    .Y(_3884_)
);

AOI21X1 _14459_ (
    .A(_3884_),
    .B(_3883_),
    .C(_3882_),
    .Y(_3885_)
);

OAI21X1 _14460_ (
    .A(_3881_),
    .B(_3885_),
    .C(_3874_),
    .Y(_3886_)
);

AOI21X1 _14461_ (
    .A(_3607_),
    .B(_3609_),
    .C(_3615_),
    .Y(_3888_)
);

NAND3X1 _14462_ (
    .A(_3882_),
    .B(_3884_),
    .C(_3883_),
    .Y(_3889_)
);

AND2X2 _14463_ (
    .A(_3879_),
    .B(_3877_),
    .Y(_3890_)
);

NOR2X1 _14464_ (
    .A(_3879_),
    .B(_3877_),
    .Y(_3891_)
);

OAI21X1 _14465_ (
    .A(_3890_),
    .B(_3891_),
    .C(_3875_),
    .Y(_3892_)
);

NAND3X1 _14466_ (
    .A(_3888_),
    .B(_3889_),
    .C(_3892_),
    .Y(_3893_)
);

AOI21X1 _14467_ (
    .A(_3886_),
    .B(_3893_),
    .C(_3873_),
    .Y(_3894_)
);

INVX1 _14468_ (
    .A(_3869_),
    .Y(_3895_)
);

XNOR2X1 _14469_ (
    .A(_3872_),
    .B(_3895_),
    .Y(_3896_)
);

NAND3X1 _14470_ (
    .A(_3889_),
    .B(_3874_),
    .C(_3892_),
    .Y(_3897_)
);

OAI21X1 _14471_ (
    .A(_3881_),
    .B(_3885_),
    .C(_3888_),
    .Y(_3899_)
);

AOI21X1 _14472_ (
    .A(_3899_),
    .B(_3897_),
    .C(_3896_),
    .Y(_3900_)
);

AOI21X1 _14473_ (
    .A(_3641_),
    .B(_3660_),
    .C(_3663_),
    .Y(_3901_)
);

OAI21X1 _14474_ (
    .A(_3894_),
    .B(_3900_),
    .C(_3901_),
    .Y(_3902_)
);

NAND3X1 _14475_ (
    .A(_3897_),
    .B(_3899_),
    .C(_3896_),
    .Y(_3903_)
);

NAND3X1 _14476_ (
    .A(_3886_),
    .B(_3893_),
    .C(_3873_),
    .Y(_3904_)
);

OAI21X1 _14477_ (
    .A(_3662_),
    .B(_3664_),
    .C(_3654_),
    .Y(_3905_)
);

NAND3X1 _14478_ (
    .A(_3903_),
    .B(_3904_),
    .C(_3905_),
    .Y(_3906_)
);

NAND3X1 _14479_ (
    .A(_3868_),
    .B(_3902_),
    .C(_3906_),
    .Y(_3907_)
);

AND2X2 _14480_ (
    .A(_3628_),
    .B(_3622_),
    .Y(_3908_)
);

AOI21X1 _14481_ (
    .A(_3903_),
    .B(_3904_),
    .C(_3905_),
    .Y(_3910_)
);

NOR3X1 _14482_ (
    .A(_3894_),
    .B(_3900_),
    .C(_3901_),
    .Y(_3911_)
);

OAI21X1 _14483_ (
    .A(_3911_),
    .B(_3910_),
    .C(_3908_),
    .Y(_3912_)
);

NAND2X1 _14484_ (
    .A(_3907_),
    .B(_3912_),
    .Y(_3913_)
);

AOI21X1 _14485_ (
    .A(_3705_),
    .B(_3704_),
    .C(_3669_),
    .Y(_3914_)
);

OAI21X1 _14486_ (
    .A(_3666_),
    .B(_3914_),
    .C(_3711_),
    .Y(_3915_)
);

NAND2X1 _14487_ (
    .A(breg_7_bF$buf0),
    .B(areg_14_bF$buf2),
    .Y(_3916_)
);

OAI21X1 _14488_ (
    .A(_3640_),
    .B(_3916_),
    .C(_3648_),
    .Y(_3917_)
);

NOR2X1 _14489_ (
    .A(_5420__bF$buf1),
    .B(_549__bF$buf2),
    .Y(_3918_)
);

AND2X2 _14490_ (
    .A(breg_7_bF$buf5),
    .B(areg_14_bF$buf1),
    .Y(_3919_)
);

AND2X2 _14491_ (
    .A(breg_6_bF$buf0),
    .B(areg_15_bF$buf3),
    .Y(_3921_)
);

NAND2X1 _14492_ (
    .A(_3919_),
    .B(_3921_),
    .Y(_3922_)
);

OAI21X1 _14493_ (
    .A(_5453__bF$buf3),
    .B(_2465__bF$buf1),
    .C(_3916_),
    .Y(_3923_)
);

NAND3X1 _14494_ (
    .A(_3918_),
    .B(_3923_),
    .C(_3922_),
    .Y(_3924_)
);

INVX1 _14495_ (
    .A(_3918_),
    .Y(_3925_)
);

OAI21X1 _14496_ (
    .A(_4116__bF$buf3),
    .B(_2287__bF$buf2),
    .C(_3921_),
    .Y(_3926_)
);

OAI21X1 _14497_ (
    .A(_5453__bF$buf2),
    .B(_2465__bF$buf0),
    .C(_3919_),
    .Y(_3927_)
);

NAND3X1 _14498_ (
    .A(_3926_),
    .B(_3927_),
    .C(_3925_),
    .Y(_3928_)
);

INVX1 _14499_ (
    .A(_3670_),
    .Y(_3929_)
);

AND2X2 _14500_ (
    .A(breg_3_bF$buf5),
    .B(areg_17_bF$buf4),
    .Y(_3930_)
);

NAND2X1 _14501_ (
    .A(_3930_),
    .B(_3391_),
    .Y(_3932_)
);

OAI21X1 _14502_ (
    .A(_3929_),
    .B(_3674_),
    .C(_3932_),
    .Y(_3933_)
);

NAND3X1 _14503_ (
    .A(_3924_),
    .B(_3928_),
    .C(_3933_),
    .Y(_3934_)
);

AOI21X1 _14504_ (
    .A(_3926_),
    .B(_3927_),
    .C(_3925_),
    .Y(_3935_)
);

AOI21X1 _14505_ (
    .A(_3923_),
    .B(_3922_),
    .C(_3918_),
    .Y(_3936_)
);

INVX1 _14506_ (
    .A(_3674_),
    .Y(_3937_)
);

AOI22X1 _14507_ (
    .A(_3671_),
    .B(_3673_),
    .C(_3937_),
    .D(_3670_),
    .Y(_3938_)
);

OAI21X1 _14508_ (
    .A(_3935_),
    .B(_3936_),
    .C(_3938_),
    .Y(_3939_)
);

NAND3X1 _14509_ (
    .A(_3917_),
    .B(_3939_),
    .C(_3934_),
    .Y(_3940_)
);

INVX2 _14510_ (
    .A(_3917_),
    .Y(_3941_)
);

NOR3X1 _14511_ (
    .A(_3936_),
    .B(_3938_),
    .C(_3935_),
    .Y(_3943_)
);

AOI21X1 _14512_ (
    .A(_3924_),
    .B(_3928_),
    .C(_3933_),
    .Y(_3944_)
);

OAI21X1 _14513_ (
    .A(_3943_),
    .B(_3944_),
    .C(_3941_),
    .Y(_3945_)
);

NAND2X1 _14514_ (
    .A(_3940_),
    .B(_3945_),
    .Y(_3946_)
);

AOI21X1 _14515_ (
    .A(_3693_),
    .B(_3692_),
    .C(_3677_),
    .Y(_3947_)
);

OAI21X1 _14516_ (
    .A(_3676_),
    .B(_3947_),
    .C(_3697_),
    .Y(_3948_)
);

NOR2X1 _14517_ (
    .A(_4258__bF$buf2),
    .B(_2669__bF$buf2),
    .Y(_3949_)
);

NAND2X1 _14518_ (
    .A(breg_4_bF$buf3),
    .B(areg_18_bF$buf5),
    .Y(_3950_)
);

INVX1 _14519_ (
    .A(_3950_),
    .Y(_3951_)
);

AOI22X1 _14520_ (
    .A(breg_3_bF$buf4),
    .B(areg_18_bF$buf4),
    .C(breg_4_bF$buf2),
    .D(areg_17_bF$buf3),
    .Y(_3952_)
);

AOI21X1 _14521_ (
    .A(_3930_),
    .B(_3951_),
    .C(_3952_),
    .Y(_3954_)
);

XNOR2X1 _14522_ (
    .A(_3954_),
    .B(_3949_),
    .Y(_3955_)
);

OAI21X1 _14523_ (
    .A(_3678_),
    .B(_3682_),
    .C(_3686_),
    .Y(_3956_)
);

NAND2X1 _14524_ (
    .A(breg_2_bF$buf2),
    .B(areg_19_bF$buf1),
    .Y(_3957_)
);

INVX8 _14525_ (
    .A(areg_20_bF$buf1),
    .Y(_3958_)
);

AND2X2 _14526_ (
    .A(breg_0_bF$buf3),
    .B(areg_21_bF$buf4),
    .Y(_3959_)
);

OAI21X1 _14527_ (
    .A(_3220_),
    .B(_3958__bF$buf3),
    .C(_3959_),
    .Y(_3960_)
);

INVX8 _14528_ (
    .A(areg_21_bF$buf3),
    .Y(_3961_)
);

OAI21X1 _14529_ (
    .A(_2551__bF$buf1),
    .B(_3961__bF$buf4),
    .C(_3685_),
    .Y(_3962_)
);

AOI21X1 _14530_ (
    .A(_3960_),
    .B(_3962_),
    .C(_3957_),
    .Y(_3963_)
);

INVX2 _14531_ (
    .A(_3957_),
    .Y(_3965_)
);

NAND2X1 _14532_ (
    .A(_3685_),
    .B(_3959_),
    .Y(_3966_)
);

OAI21X1 _14533_ (
    .A(_2551__bF$buf0),
    .B(_3961__bF$buf3),
    .C(_3680_),
    .Y(_3967_)
);

AOI21X1 _14534_ (
    .A(_3967_),
    .B(_3966_),
    .C(_3965_),
    .Y(_3968_)
);

OAI21X1 _14535_ (
    .A(_3963_),
    .B(_3968_),
    .C(_3956_),
    .Y(_3969_)
);

AOI21X1 _14536_ (
    .A(_3684_),
    .B(_3687_),
    .C(_3681_),
    .Y(_3970_)
);

NAND3X1 _14537_ (
    .A(_3965_),
    .B(_3967_),
    .C(_3966_),
    .Y(_3971_)
);

NAND2X1 _14538_ (
    .A(breg_0_bF$buf2),
    .B(areg_21_bF$buf2),
    .Y(_3972_)
);

NOR2X1 _14539_ (
    .A(_3680_),
    .B(_3972_),
    .Y(_3973_)
);

NOR2X1 _14540_ (
    .A(_3685_),
    .B(_3959_),
    .Y(_3974_)
);

OAI21X1 _14541_ (
    .A(_3974_),
    .B(_3973_),
    .C(_3957_),
    .Y(_3976_)
);

NAND3X1 _14542_ (
    .A(_3970_),
    .B(_3971_),
    .C(_3976_),
    .Y(_3977_)
);

AOI21X1 _14543_ (
    .A(_3969_),
    .B(_3977_),
    .C(_3955_),
    .Y(_3978_)
);

XOR2X1 _14544_ (
    .A(_3954_),
    .B(_3949_),
    .Y(_3979_)
);

NAND3X1 _14545_ (
    .A(_3956_),
    .B(_3971_),
    .C(_3976_),
    .Y(_3980_)
);

OAI21X1 _14546_ (
    .A(_3963_),
    .B(_3968_),
    .C(_3970_),
    .Y(_3981_)
);

AOI21X1 _14547_ (
    .A(_3981_),
    .B(_3980_),
    .C(_3979_),
    .Y(_3982_)
);

OAI21X1 _14548_ (
    .A(_3978_),
    .B(_3982_),
    .C(_3948_),
    .Y(_3983_)
);

NOR3X1 _14549_ (
    .A(_3683_),
    .B(_3691_),
    .C(_3688_),
    .Y(_3984_)
);

AOI21X1 _14550_ (
    .A(_3696_),
    .B(_3698_),
    .C(_3984_),
    .Y(_3985_)
);

NAND3X1 _14551_ (
    .A(_3981_),
    .B(_3980_),
    .C(_3979_),
    .Y(_3987_)
);

NAND3X1 _14552_ (
    .A(_3969_),
    .B(_3977_),
    .C(_3955_),
    .Y(_3988_)
);

NAND3X1 _14553_ (
    .A(_3988_),
    .B(_3987_),
    .C(_3985_),
    .Y(_3989_)
);

AOI21X1 _14554_ (
    .A(_3989_),
    .B(_3983_),
    .C(_3946_),
    .Y(_3990_)
);

NAND3X1 _14555_ (
    .A(_3934_),
    .B(_3939_),
    .C(_3941_),
    .Y(_3991_)
);

OAI21X1 _14556_ (
    .A(_3943_),
    .B(_3944_),
    .C(_3917_),
    .Y(_3992_)
);

NAND2X1 _14557_ (
    .A(_3991_),
    .B(_3992_),
    .Y(_3993_)
);

NAND3X1 _14558_ (
    .A(_3987_),
    .B(_3988_),
    .C(_3948_),
    .Y(_3994_)
);

OAI21X1 _14559_ (
    .A(_3978_),
    .B(_3982_),
    .C(_3985_),
    .Y(_3995_)
);

AOI21X1 _14560_ (
    .A(_3994_),
    .B(_3995_),
    .C(_3993_),
    .Y(_3996_)
);

OAI21X1 _14561_ (
    .A(_3990_),
    .B(_3996_),
    .C(_3915_),
    .Y(_3998_)
);

NOR3X1 _14562_ (
    .A(_3699_),
    .B(_3695_),
    .C(_3703_),
    .Y(_3999_)
);

AOI21X1 _14563_ (
    .A(_3710_),
    .B(_3713_),
    .C(_3999_),
    .Y(_4000_)
);

NAND3X1 _14564_ (
    .A(_3994_),
    .B(_3993_),
    .C(_3995_),
    .Y(_4001_)
);

NAND3X1 _14565_ (
    .A(_3989_),
    .B(_3946_),
    .C(_3983_),
    .Y(_4002_)
);

NAND3X1 _14566_ (
    .A(_4001_),
    .B(_4002_),
    .C(_4000_),
    .Y(_4003_)
);

AOI21X1 _14567_ (
    .A(_4003_),
    .B(_3998_),
    .C(_3913_),
    .Y(_4004_)
);

OAI21X1 _14568_ (
    .A(_3911_),
    .B(_3910_),
    .C(_3868_),
    .Y(_4005_)
);

NAND3X1 _14569_ (
    .A(_3902_),
    .B(_3906_),
    .C(_3908_),
    .Y(_4006_)
);

NAND2X1 _14570_ (
    .A(_4006_),
    .B(_4005_),
    .Y(_4007_)
);

NAND3X1 _14571_ (
    .A(_4001_),
    .B(_3915_),
    .C(_4002_),
    .Y(_4009_)
);

OAI21X1 _14572_ (
    .A(_3990_),
    .B(_3996_),
    .C(_4000_),
    .Y(_4010_)
);

AOI21X1 _14573_ (
    .A(_4009_),
    .B(_4010_),
    .C(_4007_),
    .Y(_4011_)
);

OAI21X1 _14574_ (
    .A(_4004_),
    .B(_4011_),
    .C(_3867_),
    .Y(_4012_)
);

AOI21X1 _14575_ (
    .A(_3724_),
    .B(_3726_),
    .C(_3731_),
    .Y(_4013_)
);

NAND3X1 _14576_ (
    .A(_4009_),
    .B(_4010_),
    .C(_4007_),
    .Y(_4014_)
);

NAND3X1 _14577_ (
    .A(_4003_),
    .B(_3998_),
    .C(_3913_),
    .Y(_4015_)
);

NAND3X1 _14578_ (
    .A(_4014_),
    .B(_4015_),
    .C(_4013_),
    .Y(_4016_)
);

AOI21X1 _14579_ (
    .A(_4012_),
    .B(_4016_),
    .C(_3866_),
    .Y(_4017_)
);

NAND3X1 _14580_ (
    .A(_3861_),
    .B(_3859_),
    .C(_3855_),
    .Y(_4018_)
);

NAND3X1 _14581_ (
    .A(_3780_),
    .B(_3863_),
    .C(_3862_),
    .Y(_4020_)
);

NAND2X1 _14582_ (
    .A(_4020_),
    .B(_4018_),
    .Y(_4021_)
);

NAND3X1 _14583_ (
    .A(_4014_),
    .B(_4015_),
    .C(_3867_),
    .Y(_4022_)
);

OAI21X1 _14584_ (
    .A(_4004_),
    .B(_4011_),
    .C(_4013_),
    .Y(_4023_)
);

AOI21X1 _14585_ (
    .A(_4022_),
    .B(_4023_),
    .C(_4021_),
    .Y(_4024_)
);

NOR3X1 _14586_ (
    .A(_4017_),
    .B(_4024_),
    .C(_3779_),
    .Y(_4025_)
);

OAI21X1 _14587_ (
    .A(_3735_),
    .B(_3590_),
    .C(_3740_),
    .Y(_4026_)
);

NAND3X1 _14588_ (
    .A(_4022_),
    .B(_4023_),
    .C(_4021_),
    .Y(_4027_)
);

NAND3X1 _14589_ (
    .A(_4012_),
    .B(_4016_),
    .C(_3866_),
    .Y(_4028_)
);

AOI21X1 _14590_ (
    .A(_4027_),
    .B(_4028_),
    .C(_4026_),
    .Y(_4029_)
);

NOR3X1 _14591_ (
    .A(_4029_),
    .B(_3778_),
    .C(_4025_),
    .Y(_4031_)
);

XNOR2X1 _14592_ (
    .A(_3777_),
    .B(_3534_),
    .Y(_4032_)
);

NAND3X1 _14593_ (
    .A(_4027_),
    .B(_4028_),
    .C(_4026_),
    .Y(_4033_)
);

OAI21X1 _14594_ (
    .A(_4017_),
    .B(_4024_),
    .C(_3779_),
    .Y(_4034_)
);

AOI21X1 _14595_ (
    .A(_4034_),
    .B(_4033_),
    .C(_4032_),
    .Y(_4035_)
);

OAI21X1 _14596_ (
    .A(_4031_),
    .B(_4035_),
    .C(_3775_),
    .Y(_4036_)
);

AOI21X1 _14597_ (
    .A(_3520_),
    .B(_3751_),
    .C(_3758_),
    .Y(_4037_)
);

NAND3X1 _14598_ (
    .A(_4032_),
    .B(_4034_),
    .C(_4033_),
    .Y(_4038_)
);

OAI21X1 _14599_ (
    .A(_4025_),
    .B(_4029_),
    .C(_3778_),
    .Y(_4039_)
);

NAND3X1 _14600_ (
    .A(_4038_),
    .B(_4039_),
    .C(_4037_),
    .Y(_4040_)
);

AOI22X1 _14601_ (
    .A(_3519_),
    .B(_3774_),
    .C(_4040_),
    .D(_4036_),
    .Y(_4041_)
);

NAND3X1 _14602_ (
    .A(_4038_),
    .B(_4039_),
    .C(_3775_),
    .Y(_4042_)
);

OAI21X1 _14603_ (
    .A(_4031_),
    .B(_4035_),
    .C(_4037_),
    .Y(_4043_)
);

AOI21X1 _14604_ (
    .A(_4042_),
    .B(_4043_),
    .C(_3763_),
    .Y(_4044_)
);

OAI21X1 _14605_ (
    .A(_4041_),
    .B(_4044_),
    .C(_3767_),
    .Y(_4045_)
);

NAND3X1 _14606_ (
    .A(_3763_),
    .B(_3764_),
    .C(_3517_),
    .Y(_4046_)
);

AOI21X1 _14607_ (
    .A(_4036_),
    .B(_4040_),
    .C(_3763_),
    .Y(_4047_)
);

AOI22X1 _14608_ (
    .A(_3774_),
    .B(_3519_),
    .C(_4043_),
    .D(_4042_),
    .Y(_4048_)
);

OAI21X1 _14609_ (
    .A(_4047_),
    .B(_4048_),
    .C(_4046_),
    .Y(_4049_)
);

NAND2X1 _14610_ (
    .A(_4045_),
    .B(_4049_),
    .Y(_4050_)
);

XNOR2X1 _14611_ (
    .A(_3773_),
    .B(_4050_),
    .Y(_0_[21])
);

OAI21X1 _14612_ (
    .A(_4050_),
    .B(_3771_),
    .C(_4045_),
    .Y(_4052_)
);

INVX1 _14613_ (
    .A(_4052_),
    .Y(_4053_)
);

NAND3X1 _14614_ (
    .A(_4045_),
    .B(_4049_),
    .C(_3770_),
    .Y(_4054_)
);

OAI21X1 _14615_ (
    .A(_3516_),
    .B(_4054_),
    .C(_4053_),
    .Y(_4055_)
);

INVX1 _14616_ (
    .A(_4042_),
    .Y(_4056_)
);

NAND2X1 _14617_ (
    .A(_3535_),
    .B(_3777_),
    .Y(_4057_)
);

INVX2 _14618_ (
    .A(_4057_),
    .Y(_4058_)
);

OAI21X1 _14619_ (
    .A(_4029_),
    .B(_3778_),
    .C(_4033_),
    .Y(_4059_)
);

OAI21X1 _14620_ (
    .A(_3798_),
    .B(_3783_),
    .C(_3804_),
    .Y(_4060_)
);

NAND2X1 _14621_ (
    .A(_3855_),
    .B(_3860_),
    .Y(_4062_)
);

XOR2X1 _14622_ (
    .A(_4062_),
    .B(_4060_),
    .Y(_4063_)
);

AOI21X1 _14623_ (
    .A(_4014_),
    .B(_4015_),
    .C(_3867_),
    .Y(_4064_)
);

OAI21X1 _14624_ (
    .A(_3866_),
    .B(_4064_),
    .C(_4022_),
    .Y(_4065_)
);

NOR2X1 _14625_ (
    .A(_3845_),
    .B(_3846_),
    .Y(_4066_)
);

AOI21X1 _14626_ (
    .A(_3808_),
    .B(_4066_),
    .C(_3856_),
    .Y(_4067_)
);

NAND2X1 _14627_ (
    .A(areg_1_bF$buf4),
    .B(breg_22_bF$buf4),
    .Y(_4068_)
);

INVX2 _14628_ (
    .A(breg_22_bF$buf3),
    .Y(_4069_)
);

OAI22X1 _14629_ (
    .A(_2661_),
    .B(_3781__bF$buf2),
    .C(_2376__bF$buf2),
    .D(_4069_),
    .Y(_4070_)
);

OAI21X1 _14630_ (
    .A(_3783_),
    .B(_4068_),
    .C(_4070_),
    .Y(_4071_)
);

AOI21X1 _14631_ (
    .A(_3794_),
    .B(_3796_),
    .C(_3791_),
    .Y(_4073_)
);

INVX1 _14632_ (
    .A(_4073_),
    .Y(_4074_)
);

NAND2X1 _14633_ (
    .A(areg_2_bF$buf4),
    .B(breg_20_bF$buf2),
    .Y(_4075_)
);

NAND2X1 _14634_ (
    .A(areg_4_bF$buf0),
    .B(breg_19_bF$buf2),
    .Y(_4076_)
);

NOR2X1 _14635_ (
    .A(_3790_),
    .B(_4076_),
    .Y(_4077_)
);

NAND2X1 _14636_ (
    .A(areg_3_bF$buf2),
    .B(breg_19_bF$buf1),
    .Y(_4078_)
);

NAND2X1 _14637_ (
    .A(areg_4_bF$buf4),
    .B(breg_18_bF$buf1),
    .Y(_4079_)
);

AND2X2 _14638_ (
    .A(_4078_),
    .B(_4079_),
    .Y(_4080_)
);

OAI21X1 _14639_ (
    .A(_4080_),
    .B(_4077_),
    .C(_4075_),
    .Y(_4081_)
);

INVX2 _14640_ (
    .A(_4075_),
    .Y(_4082_)
);

OR2X2 _14641_ (
    .A(_4078_),
    .B(_4079_),
    .Y(_4084_)
);

OAI21X1 _14642_ (
    .A(_2562__bF$buf1),
    .B(_3529__bF$buf3),
    .C(_4078_),
    .Y(_4085_)
);

NAND3X1 _14643_ (
    .A(_4082_),
    .B(_4085_),
    .C(_4084_),
    .Y(_4086_)
);

AOI21X1 _14644_ (
    .A(_4081_),
    .B(_4086_),
    .C(_4074_),
    .Y(_4087_)
);

AOI21X1 _14645_ (
    .A(_4085_),
    .B(_4084_),
    .C(_4082_),
    .Y(_4088_)
);

NOR3X1 _14646_ (
    .A(_4075_),
    .B(_4077_),
    .C(_4080_),
    .Y(_4089_)
);

NOR3X1 _14647_ (
    .A(_4088_),
    .B(_4073_),
    .C(_4089_),
    .Y(_4090_)
);

OAI21X1 _14648_ (
    .A(_4087_),
    .B(_4090_),
    .C(_4071_),
    .Y(_4091_)
);

INVX1 _14649_ (
    .A(_4071_),
    .Y(_4092_)
);

OAI21X1 _14650_ (
    .A(_4089_),
    .B(_4088_),
    .C(_4073_),
    .Y(_4093_)
);

NAND3X1 _14651_ (
    .A(_4081_),
    .B(_4086_),
    .C(_4074_),
    .Y(_4095_)
);

NAND3X1 _14652_ (
    .A(_4092_),
    .B(_4093_),
    .C(_4095_),
    .Y(_4096_)
);

AND2X2 _14653_ (
    .A(_4091_),
    .B(_4096_),
    .Y(_4097_)
);

OAI21X1 _14654_ (
    .A(_3836_),
    .B(_3834_),
    .C(_3825_),
    .Y(_4098_)
);

OAI21X1 _14655_ (
    .A(_3818_),
    .B(_3826_),
    .C(_3814_),
    .Y(_4099_)
);

NOR2X1 _14656_ (
    .A(_2825__bF$buf2),
    .B(_2763_),
    .Y(_4100_)
);

AND2X2 _14657_ (
    .A(areg_6_bF$buf0),
    .B(breg_16_bF$buf3),
    .Y(_4101_)
);

AND2X2 _14658_ (
    .A(areg_7_bF$buf3),
    .B(breg_15_bF$buf4),
    .Y(_4102_)
);

NAND2X1 _14659_ (
    .A(_4101_),
    .B(_4102_),
    .Y(_4103_)
);

OAI21X1 _14660_ (
    .A(_4434__bF$buf2),
    .B(_2362__bF$buf4),
    .C(_3817_),
    .Y(_4104_)
);

NAND3X1 _14661_ (
    .A(_4100_),
    .B(_4104_),
    .C(_4103_),
    .Y(_4106_)
);

NAND2X1 _14662_ (
    .A(_4104_),
    .B(_4103_),
    .Y(_4107_)
);

OAI21X1 _14663_ (
    .A(_2825__bF$buf1),
    .B(_2763_),
    .C(_4107_),
    .Y(_4108_)
);

NOR2X1 _14664_ (
    .A(_3870_),
    .B(_3871_),
    .Y(_4109_)
);

OAI21X1 _14665_ (
    .A(_6582__bF$buf1),
    .B(_2586__bF$buf4),
    .C(_3870_),
    .Y(_4110_)
);

AOI21X1 _14666_ (
    .A(_3869_),
    .B(_4110_),
    .C(_4109_),
    .Y(_4111_)
);

INVX2 _14667_ (
    .A(_4111_),
    .Y(_4112_)
);

NAND3X1 _14668_ (
    .A(_4106_),
    .B(_4112_),
    .C(_4108_),
    .Y(_4113_)
);

INVX1 _14669_ (
    .A(_4100_),
    .Y(_4114_)
);

OAI21X1 _14670_ (
    .A(_3646__bF$buf0),
    .B(_2560__bF$buf2),
    .C(_4102_),
    .Y(_4115_)
);

OAI21X1 _14671_ (
    .A(_4434__bF$buf1),
    .B(_2362__bF$buf3),
    .C(_4101_),
    .Y(_4117_)
);

AOI21X1 _14672_ (
    .A(_4115_),
    .B(_4117_),
    .C(_4114_),
    .Y(_4118_)
);

AOI21X1 _14673_ (
    .A(_4104_),
    .B(_4103_),
    .C(_4100_),
    .Y(_4119_)
);

OAI21X1 _14674_ (
    .A(_4118_),
    .B(_4119_),
    .C(_4111_),
    .Y(_4120_)
);

NAND3X1 _14675_ (
    .A(_4099_),
    .B(_4120_),
    .C(_4113_),
    .Y(_4121_)
);

INVX2 _14676_ (
    .A(_4099_),
    .Y(_4122_)
);

NOR3X1 _14677_ (
    .A(_4119_),
    .B(_4111_),
    .C(_4118_),
    .Y(_4123_)
);

AOI21X1 _14678_ (
    .A(_4106_),
    .B(_4108_),
    .C(_4112_),
    .Y(_4124_)
);

OAI21X1 _14679_ (
    .A(_4124_),
    .B(_4123_),
    .C(_4122_),
    .Y(_4125_)
);

NAND3X1 _14680_ (
    .A(_4098_),
    .B(_4121_),
    .C(_4125_),
    .Y(_4126_)
);

AOI21X1 _14681_ (
    .A(_3831_),
    .B(_3809_),
    .C(_3835_),
    .Y(_4128_)
);

NAND3X1 _14682_ (
    .A(_4106_),
    .B(_4111_),
    .C(_4108_),
    .Y(_4129_)
);

OAI21X1 _14683_ (
    .A(_4118_),
    .B(_4119_),
    .C(_4112_),
    .Y(_4130_)
);

AOI21X1 _14684_ (
    .A(_4130_),
    .B(_4129_),
    .C(_4122_),
    .Y(_4131_)
);

AOI21X1 _14685_ (
    .A(_4120_),
    .B(_4113_),
    .C(_4099_),
    .Y(_4132_)
);

OAI21X1 _14686_ (
    .A(_4131_),
    .B(_4132_),
    .C(_4128_),
    .Y(_4133_)
);

NAND3X1 _14687_ (
    .A(_4097_),
    .B(_4126_),
    .C(_4133_),
    .Y(_4134_)
);

NAND2X1 _14688_ (
    .A(_4096_),
    .B(_4091_),
    .Y(_4135_)
);

OAI21X1 _14689_ (
    .A(_4131_),
    .B(_4132_),
    .C(_4098_),
    .Y(_4136_)
);

NAND3X1 _14690_ (
    .A(_4128_),
    .B(_4121_),
    .C(_4125_),
    .Y(_4137_)
);

NAND3X1 _14691_ (
    .A(_4135_),
    .B(_4137_),
    .C(_4136_),
    .Y(_4139_)
);

OAI21X1 _14692_ (
    .A(_3908_),
    .B(_3910_),
    .C(_3906_),
    .Y(_4140_)
);

NAND3X1 _14693_ (
    .A(_4140_),
    .B(_4134_),
    .C(_4139_),
    .Y(_4141_)
);

AOI21X1 _14694_ (
    .A(_4137_),
    .B(_4136_),
    .C(_4135_),
    .Y(_4142_)
);

AOI21X1 _14695_ (
    .A(_4126_),
    .B(_4133_),
    .C(_4097_),
    .Y(_4143_)
);

AOI21X1 _14696_ (
    .A(_3868_),
    .B(_3902_),
    .C(_3911_),
    .Y(_4144_)
);

OAI21X1 _14697_ (
    .A(_4143_),
    .B(_4142_),
    .C(_4144_),
    .Y(_4145_)
);

NAND3X1 _14698_ (
    .A(_4067_),
    .B(_4141_),
    .C(_4145_),
    .Y(_4146_)
);

NAND2X1 _14699_ (
    .A(_3838_),
    .B(_3848_),
    .Y(_4147_)
);

NAND3X1 _14700_ (
    .A(_4144_),
    .B(_4134_),
    .C(_4139_),
    .Y(_4148_)
);

OAI21X1 _14701_ (
    .A(_4143_),
    .B(_4142_),
    .C(_4140_),
    .Y(_4150_)
);

NAND3X1 _14702_ (
    .A(_4147_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4151_)
);

NAND2X1 _14703_ (
    .A(_4146_),
    .B(_4151_),
    .Y(_4152_)
);

AOI21X1 _14704_ (
    .A(_4001_),
    .B(_4002_),
    .C(_3915_),
    .Y(_4153_)
);

OAI21X1 _14705_ (
    .A(_3913_),
    .B(_4153_),
    .C(_4009_),
    .Y(_4154_)
);

NAND2X1 _14706_ (
    .A(_3897_),
    .B(_3903_),
    .Y(_4155_)
);

NOR2X1 _14707_ (
    .A(_5190__bF$buf1),
    .B(_2379_),
    .Y(_4156_)
);

INVX1 _14708_ (
    .A(_4156_),
    .Y(_4157_)
);

NAND2X1 _14709_ (
    .A(areg_9_bF$buf1),
    .B(breg_13_bF$buf0),
    .Y(_4158_)
);

NAND2X1 _14710_ (
    .A(areg_10_bF$buf1),
    .B(breg_12_bF$buf3),
    .Y(_4159_)
);

XOR2X1 _14711_ (
    .A(_4158_),
    .B(_4159_),
    .Y(_4161_)
);

XNOR2X1 _14712_ (
    .A(_4161_),
    .B(_4157_),
    .Y(_4162_)
);

OAI21X1 _14713_ (
    .A(_3891_),
    .B(_3875_),
    .C(_3883_),
    .Y(_4163_)
);

NAND2X1 _14714_ (
    .A(areg_11_bF$buf2),
    .B(breg_11_bF$buf0),
    .Y(_4164_)
);

INVX2 _14715_ (
    .A(_4164_),
    .Y(_4165_)
);

AND2X2 _14716_ (
    .A(breg_10_bF$buf1),
    .B(areg_12_bF$buf2),
    .Y(_4166_)
);

AND2X2 _14717_ (
    .A(breg_9_bF$buf3),
    .B(areg_13_bF$buf1),
    .Y(_4167_)
);

NAND2X1 _14718_ (
    .A(_4166_),
    .B(_4167_),
    .Y(_4168_)
);

OAI22X1 _14719_ (
    .A(_6044__bF$buf4),
    .B(_549__bF$buf1),
    .C(_7217__bF$buf4),
    .D(_10869__bF$buf0),
    .Y(_4169_)
);

NAND3X1 _14720_ (
    .A(_4165_),
    .B(_4169_),
    .C(_4168_),
    .Y(_4170_)
);

AND2X2 _14721_ (
    .A(_4166_),
    .B(_4167_),
    .Y(_4172_)
);

NOR2X1 _14722_ (
    .A(_4166_),
    .B(_4167_),
    .Y(_4173_)
);

OAI21X1 _14723_ (
    .A(_4172_),
    .B(_4173_),
    .C(_4164_),
    .Y(_4174_)
);

NAND3X1 _14724_ (
    .A(_4170_),
    .B(_4163_),
    .C(_4174_),
    .Y(_4175_)
);

AOI21X1 _14725_ (
    .A(_3882_),
    .B(_3884_),
    .C(_3890_),
    .Y(_4176_)
);

OAI21X1 _14726_ (
    .A(_7217__bF$buf3),
    .B(_10869__bF$buf3),
    .C(_4167_),
    .Y(_4177_)
);

OAI21X1 _14727_ (
    .A(_6044__bF$buf3),
    .B(_549__bF$buf0),
    .C(_4166_),
    .Y(_4178_)
);

AOI21X1 _14728_ (
    .A(_4177_),
    .B(_4178_),
    .C(_4164_),
    .Y(_4179_)
);

AOI21X1 _14729_ (
    .A(_4169_),
    .B(_4168_),
    .C(_4165_),
    .Y(_4180_)
);

OAI21X1 _14730_ (
    .A(_4179_),
    .B(_4180_),
    .C(_4176_),
    .Y(_4181_)
);

NAND3X1 _14731_ (
    .A(_4175_),
    .B(_4181_),
    .C(_4162_),
    .Y(_4183_)
);

XNOR2X1 _14732_ (
    .A(_4161_),
    .B(_4156_),
    .Y(_4184_)
);

OAI21X1 _14733_ (
    .A(_4179_),
    .B(_4180_),
    .C(_4163_),
    .Y(_4185_)
);

NAND3X1 _14734_ (
    .A(_4176_),
    .B(_4170_),
    .C(_4174_),
    .Y(_4186_)
);

NAND3X1 _14735_ (
    .A(_4185_),
    .B(_4186_),
    .C(_4184_),
    .Y(_4187_)
);

OAI21X1 _14736_ (
    .A(_3941_),
    .B(_3944_),
    .C(_3934_),
    .Y(_4188_)
);

AOI21X1 _14737_ (
    .A(_4183_),
    .B(_4187_),
    .C(_4188_),
    .Y(_4189_)
);

AOI21X1 _14738_ (
    .A(_4185_),
    .B(_4186_),
    .C(_4184_),
    .Y(_4190_)
);

AOI21X1 _14739_ (
    .A(_4181_),
    .B(_4175_),
    .C(_4162_),
    .Y(_4191_)
);

AOI21X1 _14740_ (
    .A(_3917_),
    .B(_3939_),
    .C(_3943_),
    .Y(_4192_)
);

NOR3X1 _14741_ (
    .A(_4190_),
    .B(_4191_),
    .C(_4192_),
    .Y(_4194_)
);

OAI21X1 _14742_ (
    .A(_4194_),
    .B(_4189_),
    .C(_4155_),
    .Y(_4195_)
);

AND2X2 _14743_ (
    .A(_3903_),
    .B(_3897_),
    .Y(_4196_)
);

OAI21X1 _14744_ (
    .A(_4190_),
    .B(_4191_),
    .C(_4192_),
    .Y(_4197_)
);

NAND3X1 _14745_ (
    .A(_4183_),
    .B(_4187_),
    .C(_4188_),
    .Y(_4198_)
);

NAND3X1 _14746_ (
    .A(_4196_),
    .B(_4197_),
    .C(_4198_),
    .Y(_4199_)
);

NAND2X1 _14747_ (
    .A(_4199_),
    .B(_4195_),
    .Y(_4200_)
);

AOI21X1 _14748_ (
    .A(_3988_),
    .B(_3987_),
    .C(_3948_),
    .Y(_4201_)
);

OAI21X1 _14749_ (
    .A(_3946_),
    .B(_4201_),
    .C(_3994_),
    .Y(_4202_)
);

INVX1 _14750_ (
    .A(_3921_),
    .Y(_4203_)
);

OAI21X1 _14751_ (
    .A(_3916_),
    .B(_4203_),
    .C(_3924_),
    .Y(_4205_)
);

INVX2 _14752_ (
    .A(_4205_),
    .Y(_4206_)
);

NAND2X1 _14753_ (
    .A(breg[8]),
    .B(areg_14_bF$buf0),
    .Y(_4207_)
);

INVX1 _14754_ (
    .A(_4207_),
    .Y(_4208_)
);

AND2X2 _14755_ (
    .A(breg_7_bF$buf4),
    .B(areg_15_bF$buf2),
    .Y(_4209_)
);

AND2X2 _14756_ (
    .A(breg_6_bF$buf5),
    .B(areg_16_bF$buf3),
    .Y(_4210_)
);

NAND2X1 _14757_ (
    .A(_4209_),
    .B(_4210_),
    .Y(_4211_)
);

OAI22X1 _14758_ (
    .A(_5453__bF$buf1),
    .B(_2669__bF$buf1),
    .C(_4116__bF$buf2),
    .D(_2465__bF$buf4),
    .Y(_4212_)
);

NAND3X1 _14759_ (
    .A(_4208_),
    .B(_4212_),
    .C(_4211_),
    .Y(_4213_)
);

OAI21X1 _14760_ (
    .A(_4116__bF$buf1),
    .B(_2465__bF$buf3),
    .C(_4210_),
    .Y(_4214_)
);

OAI21X1 _14761_ (
    .A(_5453__bF$buf0),
    .B(_2669__bF$buf0),
    .C(_4209_),
    .Y(_4216_)
);

NAND3X1 _14762_ (
    .A(_4207_),
    .B(_4214_),
    .C(_4216_),
    .Y(_4217_)
);

INVX1 _14763_ (
    .A(_3949_),
    .Y(_4218_)
);

AND2X2 _14764_ (
    .A(breg_3_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_4219_)
);

NAND2X1 _14765_ (
    .A(_4219_),
    .B(_3673_),
    .Y(_4220_)
);

OAI21X1 _14766_ (
    .A(_4218_),
    .B(_3952_),
    .C(_4220_),
    .Y(_4221_)
);

NAND3X1 _14767_ (
    .A(_4213_),
    .B(_4217_),
    .C(_4221_),
    .Y(_4222_)
);

AOI21X1 _14768_ (
    .A(_4214_),
    .B(_4216_),
    .C(_4207_),
    .Y(_4223_)
);

AOI21X1 _14769_ (
    .A(_4212_),
    .B(_4211_),
    .C(_4208_),
    .Y(_4224_)
);

INVX1 _14770_ (
    .A(_3952_),
    .Y(_4225_)
);

AOI22X1 _14771_ (
    .A(_3930_),
    .B(_3951_),
    .C(_4225_),
    .D(_3949_),
    .Y(_4227_)
);

OAI21X1 _14772_ (
    .A(_4223_),
    .B(_4224_),
    .C(_4227_),
    .Y(_4228_)
);

NAND3X1 _14773_ (
    .A(_4222_),
    .B(_4228_),
    .C(_4206_),
    .Y(_4229_)
);

NOR3X1 _14774_ (
    .A(_4224_),
    .B(_4227_),
    .C(_4223_),
    .Y(_4230_)
);

AOI21X1 _14775_ (
    .A(_4213_),
    .B(_4217_),
    .C(_4221_),
    .Y(_4231_)
);

OAI21X1 _14776_ (
    .A(_4230_),
    .B(_4231_),
    .C(_4205_),
    .Y(_4232_)
);

NAND2X1 _14777_ (
    .A(_4232_),
    .B(_4229_),
    .Y(_4233_)
);

AOI21X1 _14778_ (
    .A(_3971_),
    .B(_3976_),
    .C(_3956_),
    .Y(_4234_)
);

OAI21X1 _14779_ (
    .A(_4234_),
    .B(_3955_),
    .C(_3980_),
    .Y(_4235_)
);

NAND2X1 _14780_ (
    .A(breg_5_bF$buf1),
    .B(areg_17_bF$buf2),
    .Y(_4236_)
);

AND2X2 _14781_ (
    .A(breg_4_bF$buf1),
    .B(areg_19_bF$buf0),
    .Y(_4238_)
);

AOI22X1 _14782_ (
    .A(breg_3_bF$buf2),
    .B(areg_19_bF$buf5),
    .C(breg_4_bF$buf0),
    .D(areg_18_bF$buf2),
    .Y(_4239_)
);

AOI21X1 _14783_ (
    .A(_4219_),
    .B(_4238_),
    .C(_4239_),
    .Y(_4240_)
);

XNOR2X1 _14784_ (
    .A(_4240_),
    .B(_4236_),
    .Y(_4241_)
);

OAI21X1 _14785_ (
    .A(_3974_),
    .B(_3957_),
    .C(_3966_),
    .Y(_4242_)
);

NAND2X1 _14786_ (
    .A(breg_2_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_4243_)
);

INVX2 _14787_ (
    .A(_4243_),
    .Y(_4244_)
);

AND2X2 _14788_ (
    .A(breg_1_bF$buf2),
    .B(areg_22_bF$buf4),
    .Y(_4245_)
);

NAND2X1 _14789_ (
    .A(_3959_),
    .B(_4245_),
    .Y(_4246_)
);

AOI22X1 _14790_ (
    .A(breg_0_bF$buf1),
    .B(areg_22_bF$buf3),
    .C(breg_1_bF$buf1),
    .D(areg_21_bF$buf1),
    .Y(_4247_)
);

INVX2 _14791_ (
    .A(_4247_),
    .Y(_4248_)
);

NAND3X1 _14792_ (
    .A(_4244_),
    .B(_4248_),
    .C(_4246_),
    .Y(_4249_)
);

NAND2X1 _14793_ (
    .A(breg_1_bF$buf0),
    .B(areg_22_bF$buf2),
    .Y(_4250_)
);

NOR2X1 _14794_ (
    .A(_3972_),
    .B(_4250_),
    .Y(_4251_)
);

OAI21X1 _14795_ (
    .A(_4251_),
    .B(_4247_),
    .C(_4243_),
    .Y(_4252_)
);

NAND3X1 _14796_ (
    .A(_4252_),
    .B(_4249_),
    .C(_4242_),
    .Y(_4253_)
);

AOI21X1 _14797_ (
    .A(_3965_),
    .B(_3967_),
    .C(_3973_),
    .Y(_4254_)
);

NOR3X1 _14798_ (
    .A(_4243_),
    .B(_4247_),
    .C(_4251_),
    .Y(_4255_)
);

AOI21X1 _14799_ (
    .A(_4248_),
    .B(_4246_),
    .C(_4244_),
    .Y(_4256_)
);

OAI21X1 _14800_ (
    .A(_4256_),
    .B(_4255_),
    .C(_4254_),
    .Y(_4257_)
);

NAND3X1 _14801_ (
    .A(_4241_),
    .B(_4257_),
    .C(_4253_),
    .Y(_4260_)
);

INVX2 _14802_ (
    .A(_4236_),
    .Y(_4261_)
);

XNOR2X1 _14803_ (
    .A(_4240_),
    .B(_4261_),
    .Y(_4262_)
);

OAI21X1 _14804_ (
    .A(_4256_),
    .B(_4255_),
    .C(_4242_),
    .Y(_4263_)
);

NAND3X1 _14805_ (
    .A(_4254_),
    .B(_4252_),
    .C(_4249_),
    .Y(_4264_)
);

NAND3X1 _14806_ (
    .A(_4262_),
    .B(_4264_),
    .C(_4263_),
    .Y(_4265_)
);

NAND3X1 _14807_ (
    .A(_4260_),
    .B(_4265_),
    .C(_4235_),
    .Y(_4266_)
);

NOR3X1 _14808_ (
    .A(_3968_),
    .B(_3970_),
    .C(_3963_),
    .Y(_4267_)
);

AOI21X1 _14809_ (
    .A(_3981_),
    .B(_3979_),
    .C(_4267_),
    .Y(_4268_)
);

AOI21X1 _14810_ (
    .A(_4264_),
    .B(_4263_),
    .C(_4262_),
    .Y(_4269_)
);

AOI21X1 _14811_ (
    .A(_4257_),
    .B(_4253_),
    .C(_4241_),
    .Y(_4271_)
);

OAI21X1 _14812_ (
    .A(_4271_),
    .B(_4269_),
    .C(_4268_),
    .Y(_4272_)
);

NAND3X1 _14813_ (
    .A(_4233_),
    .B(_4266_),
    .C(_4272_),
    .Y(_4273_)
);

NAND3X1 _14814_ (
    .A(_4205_),
    .B(_4228_),
    .C(_4222_),
    .Y(_4274_)
);

OAI21X1 _14815_ (
    .A(_4230_),
    .B(_4231_),
    .C(_4206_),
    .Y(_4275_)
);

NAND2X1 _14816_ (
    .A(_4274_),
    .B(_4275_),
    .Y(_4276_)
);

OAI21X1 _14817_ (
    .A(_4271_),
    .B(_4269_),
    .C(_4235_),
    .Y(_4277_)
);

NAND3X1 _14818_ (
    .A(_4260_),
    .B(_4265_),
    .C(_4268_),
    .Y(_4278_)
);

NAND3X1 _14819_ (
    .A(_4276_),
    .B(_4278_),
    .C(_4277_),
    .Y(_4279_)
);

NAND3X1 _14820_ (
    .A(_4279_),
    .B(_4273_),
    .C(_4202_),
    .Y(_4280_)
);

NOR3X1 _14821_ (
    .A(_3978_),
    .B(_3982_),
    .C(_3985_),
    .Y(_4282_)
);

AOI21X1 _14822_ (
    .A(_3993_),
    .B(_3995_),
    .C(_4282_),
    .Y(_4283_)
);

AOI21X1 _14823_ (
    .A(_4278_),
    .B(_4277_),
    .C(_4276_),
    .Y(_4284_)
);

AOI21X1 _14824_ (
    .A(_4266_),
    .B(_4272_),
    .C(_4233_),
    .Y(_4285_)
);

OAI21X1 _14825_ (
    .A(_4284_),
    .B(_4285_),
    .C(_4283_),
    .Y(_4286_)
);

NAND3X1 _14826_ (
    .A(_4280_),
    .B(_4286_),
    .C(_4200_),
    .Y(_4287_)
);

NAND3X1 _14827_ (
    .A(_4155_),
    .B(_4197_),
    .C(_4198_),
    .Y(_4288_)
);

OAI21X1 _14828_ (
    .A(_4194_),
    .B(_4189_),
    .C(_4196_),
    .Y(_4289_)
);

NAND2X1 _14829_ (
    .A(_4288_),
    .B(_4289_),
    .Y(_4290_)
);

OAI21X1 _14830_ (
    .A(_4284_),
    .B(_4285_),
    .C(_4202_),
    .Y(_4291_)
);

NAND3X1 _14831_ (
    .A(_4273_),
    .B(_4279_),
    .C(_4283_),
    .Y(_4293_)
);

NAND3X1 _14832_ (
    .A(_4291_),
    .B(_4293_),
    .C(_4290_),
    .Y(_4294_)
);

NAND3X1 _14833_ (
    .A(_4287_),
    .B(_4294_),
    .C(_4154_),
    .Y(_4295_)
);

NOR3X1 _14834_ (
    .A(_3990_),
    .B(_3996_),
    .C(_4000_),
    .Y(_4296_)
);

AOI21X1 _14835_ (
    .A(_4007_),
    .B(_4010_),
    .C(_4296_),
    .Y(_4297_)
);

AOI21X1 _14836_ (
    .A(_4291_),
    .B(_4293_),
    .C(_4290_),
    .Y(_4298_)
);

AOI21X1 _14837_ (
    .A(_4280_),
    .B(_4286_),
    .C(_4200_),
    .Y(_4299_)
);

OAI21X1 _14838_ (
    .A(_4298_),
    .B(_4299_),
    .C(_4297_),
    .Y(_4300_)
);

NAND3X1 _14839_ (
    .A(_4295_),
    .B(_4300_),
    .C(_4152_),
    .Y(_4301_)
);

NAND3X1 _14840_ (
    .A(_4147_),
    .B(_4141_),
    .C(_4145_),
    .Y(_4302_)
);

NAND3X1 _14841_ (
    .A(_4067_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4304_)
);

NAND2X1 _14842_ (
    .A(_4302_),
    .B(_4304_),
    .Y(_4305_)
);

OAI21X1 _14843_ (
    .A(_4298_),
    .B(_4299_),
    .C(_4154_),
    .Y(_4306_)
);

NAND3X1 _14844_ (
    .A(_4287_),
    .B(_4294_),
    .C(_4297_),
    .Y(_4307_)
);

NAND3X1 _14845_ (
    .A(_4307_),
    .B(_4306_),
    .C(_4305_),
    .Y(_4308_)
);

NAND3X1 _14846_ (
    .A(_4301_),
    .B(_4308_),
    .C(_4065_),
    .Y(_4309_)
);

NOR3X1 _14847_ (
    .A(_4004_),
    .B(_4011_),
    .C(_4013_),
    .Y(_4310_)
);

AOI21X1 _14848_ (
    .A(_4021_),
    .B(_4023_),
    .C(_4310_),
    .Y(_4311_)
);

AOI21X1 _14849_ (
    .A(_4306_),
    .B(_4307_),
    .C(_4305_),
    .Y(_4312_)
);

AOI21X1 _14850_ (
    .A(_4295_),
    .B(_4300_),
    .C(_4152_),
    .Y(_4313_)
);

OAI21X1 _14851_ (
    .A(_4312_),
    .B(_4313_),
    .C(_4311_),
    .Y(_4315_)
);

NAND3X1 _14852_ (
    .A(_4063_),
    .B(_4309_),
    .C(_4315_),
    .Y(_4316_)
);

XNOR2X1 _14853_ (
    .A(_4062_),
    .B(_4060_),
    .Y(_4317_)
);

OAI21X1 _14854_ (
    .A(_4312_),
    .B(_4313_),
    .C(_4065_),
    .Y(_4318_)
);

NAND3X1 _14855_ (
    .A(_4301_),
    .B(_4308_),
    .C(_4311_),
    .Y(_4319_)
);

NAND3X1 _14856_ (
    .A(_4317_),
    .B(_4318_),
    .C(_4319_),
    .Y(_4320_)
);

NAND3X1 _14857_ (
    .A(_4316_),
    .B(_4320_),
    .C(_4059_),
    .Y(_4321_)
);

AOI21X1 _14858_ (
    .A(_4032_),
    .B(_4034_),
    .C(_4025_),
    .Y(_4322_)
);

AOI21X1 _14859_ (
    .A(_4318_),
    .B(_4319_),
    .C(_4317_),
    .Y(_4323_)
);

AOI21X1 _14860_ (
    .A(_4309_),
    .B(_4315_),
    .C(_4063_),
    .Y(_4324_)
);

OAI21X1 _14861_ (
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4326_)
);

NAND3X1 _14862_ (
    .A(_4058_),
    .B(_4326_),
    .C(_4321_),
    .Y(_4327_)
);

OAI21X1 _14863_ (
    .A(_4323_),
    .B(_4324_),
    .C(_4059_),
    .Y(_4328_)
);

NAND3X1 _14864_ (
    .A(_4316_),
    .B(_4320_),
    .C(_4322_),
    .Y(_4329_)
);

NAND3X1 _14865_ (
    .A(_4057_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4330_)
);

NAND3X1 _14866_ (
    .A(_4327_),
    .B(_4056_),
    .C(_4330_),
    .Y(_4331_)
);

NAND3X1 _14867_ (
    .A(_4057_),
    .B(_4326_),
    .C(_4321_),
    .Y(_4332_)
);

NAND3X1 _14868_ (
    .A(_4058_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4333_)
);

NAND3X1 _14869_ (
    .A(_4042_),
    .B(_4332_),
    .C(_4333_),
    .Y(_4334_)
);

NAND3X1 _14870_ (
    .A(_4047_),
    .B(_4334_),
    .C(_4331_),
    .Y(_4335_)
);

NOR3X1 _14871_ (
    .A(_3749_),
    .B(_3752_),
    .C(_3755_),
    .Y(_4337_)
);

NAND3X1 _14872_ (
    .A(_4042_),
    .B(_4043_),
    .C(_4337_),
    .Y(_4338_)
);

AOI21X1 _14873_ (
    .A(_4332_),
    .B(_4333_),
    .C(_4042_),
    .Y(_4339_)
);

AOI21X1 _14874_ (
    .A(_4327_),
    .B(_4330_),
    .C(_4056_),
    .Y(_4340_)
);

OAI21X1 _14875_ (
    .A(_4339_),
    .B(_4340_),
    .C(_4338_),
    .Y(_4341_)
);

NAND2X1 _14876_ (
    .A(_4335_),
    .B(_4341_),
    .Y(_4342_)
);

XNOR2X1 _14877_ (
    .A(_4055_),
    .B(_4342_),
    .Y(_0_[22])
);

AND2X2 _14878_ (
    .A(_4341_),
    .B(_4335_),
    .Y(_4343_)
);

NAND2X1 _14879_ (
    .A(_4343_),
    .B(_4055_),
    .Y(_4344_)
);

NAND2X1 _14880_ (
    .A(_4335_),
    .B(_4344_),
    .Y(_4345_)
);

AOI21X1 _14881_ (
    .A(_4316_),
    .B(_4320_),
    .C(_4059_),
    .Y(_4347_)
);

OAI21X1 _14882_ (
    .A(_4347_),
    .B(_4057_),
    .C(_4321_),
    .Y(_4348_)
);

NAND2X1 _14883_ (
    .A(_4060_),
    .B(_4062_),
    .Y(_4349_)
);

INVX2 _14884_ (
    .A(_4349_),
    .Y(_4350_)
);

AOI21X1 _14885_ (
    .A(_4301_),
    .B(_4308_),
    .C(_4065_),
    .Y(_4351_)
);

OAI21X1 _14886_ (
    .A(_4351_),
    .B(_4317_),
    .C(_4309_),
    .Y(_4352_)
);

OR2X2 _14887_ (
    .A(_3783_),
    .B(_4068_),
    .Y(_4353_)
);

NOR2X1 _14888_ (
    .A(_4353_),
    .B(_4095_),
    .Y(_4354_)
);

AND2X2 _14889_ (
    .A(_4095_),
    .B(_4353_),
    .Y(_4355_)
);

AOI21X1 _14890_ (
    .A(_4096_),
    .B(_4355_),
    .C(_4354_),
    .Y(_4356_)
);

NAND2X1 _14891_ (
    .A(_4141_),
    .B(_4302_),
    .Y(_4358_)
);

XOR2X1 _14892_ (
    .A(_4358_),
    .B(_4356_),
    .Y(_4359_)
);

AOI21X1 _14893_ (
    .A(_4287_),
    .B(_4294_),
    .C(_4154_),
    .Y(_4360_)
);

OAI21X1 _14894_ (
    .A(_4305_),
    .B(_4360_),
    .C(_4295_),
    .Y(_4361_)
);

AND2X2 _14895_ (
    .A(_4134_),
    .B(_4126_),
    .Y(_4362_)
);

NAND2X1 _14896_ (
    .A(areg[0]),
    .B(breg_23_bF$buf3),
    .Y(_4363_)
);

NAND2X1 _14897_ (
    .A(areg_2_bF$buf3),
    .B(breg_21_bF$buf3),
    .Y(_4364_)
);

XOR2X1 _14898_ (
    .A(_4068_),
    .B(_4364_),
    .Y(_4365_)
);

XNOR2X1 _14899_ (
    .A(_4365_),
    .B(_4363_),
    .Y(_4366_)
);

INVX1 _14900_ (
    .A(_4366_),
    .Y(_4367_)
);

AOI21X1 _14901_ (
    .A(_4082_),
    .B(_4085_),
    .C(_4077_),
    .Y(_4369_)
);

NAND2X1 _14902_ (
    .A(areg_3_bF$buf1),
    .B(breg_20_bF$buf1),
    .Y(_4370_)
);

NAND2X1 _14903_ (
    .A(areg_5_bF$buf4),
    .B(breg_18_bF$buf0),
    .Y(_4371_)
);

NOR2X1 _14904_ (
    .A(_4076_),
    .B(_4371_),
    .Y(_4372_)
);

AND2X2 _14905_ (
    .A(_4076_),
    .B(_4371_),
    .Y(_4373_)
);

NOR3X1 _14906_ (
    .A(_4370_),
    .B(_4372_),
    .C(_4373_),
    .Y(_4374_)
);

INVX2 _14907_ (
    .A(_4370_),
    .Y(_4375_)
);

OR2X2 _14908_ (
    .A(_4076_),
    .B(_4371_),
    .Y(_4376_)
);

OAI21X1 _14909_ (
    .A(_2825__bF$buf0),
    .B(_3529__bF$buf2),
    .C(_4076_),
    .Y(_4377_)
);

AOI21X1 _14910_ (
    .A(_4377_),
    .B(_4376_),
    .C(_4375_),
    .Y(_4378_)
);

OAI21X1 _14911_ (
    .A(_4374_),
    .B(_4378_),
    .C(_4369_),
    .Y(_4380_)
);

OAI21X1 _14912_ (
    .A(_4080_),
    .B(_4075_),
    .C(_4084_),
    .Y(_4381_)
);

NAND3X1 _14913_ (
    .A(_4375_),
    .B(_4377_),
    .C(_4376_),
    .Y(_4382_)
);

OAI21X1 _14914_ (
    .A(_4373_),
    .B(_4372_),
    .C(_4370_),
    .Y(_4383_)
);

NAND3X1 _14915_ (
    .A(_4381_),
    .B(_4383_),
    .C(_4382_),
    .Y(_4384_)
);

NAND2X1 _14916_ (
    .A(_4384_),
    .B(_4380_),
    .Y(_4385_)
);

NAND2X1 _14917_ (
    .A(_4385_),
    .B(_4367_),
    .Y(_4386_)
);

NAND3X1 _14918_ (
    .A(_4380_),
    .B(_4384_),
    .C(_4366_),
    .Y(_4387_)
);

AND2X2 _14919_ (
    .A(_4386_),
    .B(_4387_),
    .Y(_4388_)
);

OAI21X1 _14920_ (
    .A(_4124_),
    .B(_4122_),
    .C(_4113_),
    .Y(_4389_)
);

OAI21X1 _14921_ (
    .A(_4107_),
    .B(_4114_),
    .C(_4103_),
    .Y(_4391_)
);

NAND2X1 _14922_ (
    .A(areg_6_bF$buf4),
    .B(breg_17_bF$buf2),
    .Y(_4392_)
);

INVX1 _14923_ (
    .A(_4392_),
    .Y(_4393_)
);

AND2X2 _14924_ (
    .A(areg_7_bF$buf2),
    .B(breg_16_bF$buf2),
    .Y(_4394_)
);

AND2X2 _14925_ (
    .A(areg_8_bF$buf1),
    .B(breg_15_bF$buf3),
    .Y(_4395_)
);

NAND2X1 _14926_ (
    .A(_4394_),
    .B(_4395_),
    .Y(_4396_)
);

NAND2X1 _14927_ (
    .A(areg_7_bF$buf1),
    .B(breg_16_bF$buf1),
    .Y(_4397_)
);

OAI21X1 _14928_ (
    .A(_5190__bF$buf0),
    .B(_2362__bF$buf2),
    .C(_4397_),
    .Y(_4398_)
);

NAND3X1 _14929_ (
    .A(_4393_),
    .B(_4398_),
    .C(_4396_),
    .Y(_4399_)
);

NAND2X1 _14930_ (
    .A(areg_8_bF$buf0),
    .B(breg_15_bF$buf2),
    .Y(_4400_)
);

NOR2X1 _14931_ (
    .A(_4397_),
    .B(_4400_),
    .Y(_4402_)
);

NOR2X1 _14932_ (
    .A(_4394_),
    .B(_4395_),
    .Y(_4403_)
);

OAI21X1 _14933_ (
    .A(_4403_),
    .B(_4402_),
    .C(_4392_),
    .Y(_4404_)
);

NOR2X1 _14934_ (
    .A(_4158_),
    .B(_4159_),
    .Y(_4405_)
);

OAI21X1 _14935_ (
    .A(_7711__bF$buf1),
    .B(_2586__bF$buf3),
    .C(_4158_),
    .Y(_4406_)
);

AOI21X1 _14936_ (
    .A(_4156_),
    .B(_4406_),
    .C(_4405_),
    .Y(_4407_)
);

INVX2 _14937_ (
    .A(_4407_),
    .Y(_4408_)
);

NAND3X1 _14938_ (
    .A(_4399_),
    .B(_4404_),
    .C(_4408_),
    .Y(_4409_)
);

NOR3X1 _14939_ (
    .A(_4392_),
    .B(_4402_),
    .C(_4403_),
    .Y(_4410_)
);

AOI21X1 _14940_ (
    .A(_4398_),
    .B(_4396_),
    .C(_4393_),
    .Y(_4411_)
);

OAI21X1 _14941_ (
    .A(_4410_),
    .B(_4411_),
    .C(_4407_),
    .Y(_4413_)
);

NAND3X1 _14942_ (
    .A(_4391_),
    .B(_4413_),
    .C(_4409_),
    .Y(_4414_)
);

INVX2 _14943_ (
    .A(_4391_),
    .Y(_4415_)
);

NOR3X1 _14944_ (
    .A(_4411_),
    .B(_4407_),
    .C(_4410_),
    .Y(_4416_)
);

AOI21X1 _14945_ (
    .A(_4399_),
    .B(_4404_),
    .C(_4408_),
    .Y(_4417_)
);

OAI21X1 _14946_ (
    .A(_4416_),
    .B(_4417_),
    .C(_4415_),
    .Y(_4418_)
);

NAND3X1 _14947_ (
    .A(_4414_),
    .B(_4418_),
    .C(_4389_),
    .Y(_4419_)
);

AOI21X1 _14948_ (
    .A(_4099_),
    .B(_4120_),
    .C(_4123_),
    .Y(_4420_)
);

NAND3X1 _14949_ (
    .A(_4399_),
    .B(_4407_),
    .C(_4404_),
    .Y(_4421_)
);

OAI21X1 _14950_ (
    .A(_4410_),
    .B(_4411_),
    .C(_4408_),
    .Y(_4422_)
);

AOI21X1 _14951_ (
    .A(_4421_),
    .B(_4422_),
    .C(_4415_),
    .Y(_4424_)
);

AOI21X1 _14952_ (
    .A(_4413_),
    .B(_4409_),
    .C(_4391_),
    .Y(_4425_)
);

OAI21X1 _14953_ (
    .A(_4425_),
    .B(_4424_),
    .C(_4420_),
    .Y(_4426_)
);

NAND3X1 _14954_ (
    .A(_4419_),
    .B(_4426_),
    .C(_4388_),
    .Y(_4427_)
);

NAND2X1 _14955_ (
    .A(_4387_),
    .B(_4386_),
    .Y(_4428_)
);

OAI21X1 _14956_ (
    .A(_4425_),
    .B(_4424_),
    .C(_4389_),
    .Y(_4429_)
);

NAND3X1 _14957_ (
    .A(_4420_),
    .B(_4414_),
    .C(_4418_),
    .Y(_4430_)
);

NAND3X1 _14958_ (
    .A(_4430_),
    .B(_4429_),
    .C(_4428_),
    .Y(_4431_)
);

OAI21X1 _14959_ (
    .A(_4189_),
    .B(_4196_),
    .C(_4198_),
    .Y(_4432_)
);

NAND3X1 _14960_ (
    .A(_4431_),
    .B(_4432_),
    .C(_4427_),
    .Y(_4433_)
);

AOI21X1 _14961_ (
    .A(_4430_),
    .B(_4429_),
    .C(_4428_),
    .Y(_4435_)
);

AOI21X1 _14962_ (
    .A(_4419_),
    .B(_4426_),
    .C(_4388_),
    .Y(_4436_)
);

AOI21X1 _14963_ (
    .A(_4155_),
    .B(_4197_),
    .C(_4194_),
    .Y(_4437_)
);

OAI21X1 _14964_ (
    .A(_4436_),
    .B(_4435_),
    .C(_4437_),
    .Y(_4438_)
);

NAND3X1 _14965_ (
    .A(_4362_),
    .B(_4433_),
    .C(_4438_),
    .Y(_4439_)
);

NAND2X1 _14966_ (
    .A(_4126_),
    .B(_4134_),
    .Y(_4440_)
);

NAND3X1 _14967_ (
    .A(_4431_),
    .B(_4437_),
    .C(_4427_),
    .Y(_4441_)
);

OAI21X1 _14968_ (
    .A(_4436_),
    .B(_4435_),
    .C(_4432_),
    .Y(_4442_)
);

NAND3X1 _14969_ (
    .A(_4440_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4443_)
);

NAND2X1 _14970_ (
    .A(_4439_),
    .B(_4443_),
    .Y(_4444_)
);

AOI21X1 _14971_ (
    .A(_4279_),
    .B(_4273_),
    .C(_4202_),
    .Y(_4446_)
);

OAI21X1 _14972_ (
    .A(_4290_),
    .B(_4446_),
    .C(_4280_),
    .Y(_4447_)
);

NAND2X1 _14973_ (
    .A(_4175_),
    .B(_4183_),
    .Y(_4448_)
);

NAND2X1 _14974_ (
    .A(areg_9_bF$buf0),
    .B(breg_14_bF$buf3),
    .Y(_4449_)
);

NAND2X1 _14975_ (
    .A(areg_10_bF$buf0),
    .B(breg_13_bF$buf4),
    .Y(_4450_)
);

NAND2X1 _14976_ (
    .A(areg_11_bF$buf1),
    .B(breg_12_bF$buf2),
    .Y(_4451_)
);

XOR2X1 _14977_ (
    .A(_4450_),
    .B(_4451_),
    .Y(_4452_)
);

XNOR2X1 _14978_ (
    .A(_4452_),
    .B(_4449_),
    .Y(_4453_)
);

OAI21X1 _14979_ (
    .A(_4173_),
    .B(_4164_),
    .C(_4168_),
    .Y(_4454_)
);

NAND2X1 _14980_ (
    .A(breg_11_bF$buf4),
    .B(areg_12_bF$buf1),
    .Y(_4455_)
);

INVX2 _14981_ (
    .A(_4455_),
    .Y(_4456_)
);

AND2X2 _14982_ (
    .A(breg_10_bF$buf0),
    .B(areg_13_bF$buf0),
    .Y(_4457_)
);

AND2X2 _14983_ (
    .A(breg_9_bF$buf2),
    .B(areg_14_bF$buf4),
    .Y(_4458_)
);

NAND2X1 _14984_ (
    .A(_4457_),
    .B(_4458_),
    .Y(_4459_)
);

NAND2X1 _14985_ (
    .A(breg_10_bF$buf5),
    .B(areg_13_bF$buf4),
    .Y(_4460_)
);

OAI21X1 _14986_ (
    .A(_6044__bF$buf2),
    .B(_2287__bF$buf1),
    .C(_4460_),
    .Y(_4461_)
);

NAND3X1 _14987_ (
    .A(_4456_),
    .B(_4461_),
    .C(_4459_),
    .Y(_4462_)
);

NAND2X1 _14988_ (
    .A(breg_9_bF$buf1),
    .B(areg_14_bF$buf3),
    .Y(_4463_)
);

NOR2X1 _14989_ (
    .A(_4460_),
    .B(_4463_),
    .Y(_4464_)
);

NOR2X1 _14990_ (
    .A(_4457_),
    .B(_4458_),
    .Y(_4465_)
);

OAI21X1 _14991_ (
    .A(_4465_),
    .B(_4464_),
    .C(_4455_),
    .Y(_4467_)
);

NAND3X1 _14992_ (
    .A(_4462_),
    .B(_4454_),
    .C(_4467_),
    .Y(_4468_)
);

AOI21X1 _14993_ (
    .A(_4165_),
    .B(_4169_),
    .C(_4172_),
    .Y(_4469_)
);

OAI21X1 _14994_ (
    .A(_7217__bF$buf2),
    .B(_549__bF$buf4),
    .C(_4458_),
    .Y(_4470_)
);

OAI21X1 _14995_ (
    .A(_6044__bF$buf1),
    .B(_2287__bF$buf0),
    .C(_4457_),
    .Y(_4471_)
);

AOI21X1 _14996_ (
    .A(_4470_),
    .B(_4471_),
    .C(_4455_),
    .Y(_4472_)
);

AOI21X1 _14997_ (
    .A(_4461_),
    .B(_4459_),
    .C(_4456_),
    .Y(_4473_)
);

OAI21X1 _14998_ (
    .A(_4472_),
    .B(_4473_),
    .C(_4469_),
    .Y(_4474_)
);

NAND3X1 _14999_ (
    .A(_4468_),
    .B(_4474_),
    .C(_4453_),
    .Y(_4475_)
);

INVX2 _15000_ (
    .A(_4449_),
    .Y(_4476_)
);

XNOR2X1 _15001_ (
    .A(_4452_),
    .B(_4476_),
    .Y(_4479_)
);

OAI21X1 _15002_ (
    .A(_4472_),
    .B(_4473_),
    .C(_4454_),
    .Y(_4480_)
);

NAND3X1 _15003_ (
    .A(_4462_),
    .B(_4467_),
    .C(_4469_),
    .Y(_4481_)
);

NAND3X1 _15004_ (
    .A(_4480_),
    .B(_4481_),
    .C(_4479_),
    .Y(_4482_)
);

OAI21X1 _15005_ (
    .A(_4206_),
    .B(_4231_),
    .C(_4222_),
    .Y(_4483_)
);

AOI21X1 _15006_ (
    .A(_4475_),
    .B(_4482_),
    .C(_4483_),
    .Y(_4484_)
);

AOI21X1 _15007_ (
    .A(_4480_),
    .B(_4481_),
    .C(_4479_),
    .Y(_4485_)
);

AOI21X1 _15008_ (
    .A(_4468_),
    .B(_4474_),
    .C(_4453_),
    .Y(_4486_)
);

AOI21X1 _15009_ (
    .A(_4205_),
    .B(_4228_),
    .C(_4230_),
    .Y(_4487_)
);

NOR3X1 _15010_ (
    .A(_4486_),
    .B(_4487_),
    .C(_4485_),
    .Y(_4488_)
);

OAI21X1 _15011_ (
    .A(_4488_),
    .B(_4484_),
    .C(_4448_),
    .Y(_4490_)
);

AND2X2 _15012_ (
    .A(_4183_),
    .B(_4175_),
    .Y(_4491_)
);

OAI21X1 _15013_ (
    .A(_4485_),
    .B(_4486_),
    .C(_4487_),
    .Y(_4492_)
);

NAND3X1 _15014_ (
    .A(_4475_),
    .B(_4482_),
    .C(_4483_),
    .Y(_4493_)
);

NAND3X1 _15015_ (
    .A(_4491_),
    .B(_4492_),
    .C(_4493_),
    .Y(_4494_)
);

NAND2X1 _15016_ (
    .A(_4494_),
    .B(_4490_),
    .Y(_4495_)
);

AOI21X1 _15017_ (
    .A(_4260_),
    .B(_4265_),
    .C(_4235_),
    .Y(_4496_)
);

OAI21X1 _15018_ (
    .A(_4496_),
    .B(_4276_),
    .C(_4266_),
    .Y(_4497_)
);

NAND2X1 _15019_ (
    .A(breg_7_bF$buf3),
    .B(areg_16_bF$buf2),
    .Y(_4498_)
);

OAI21X1 _15020_ (
    .A(_4203_),
    .B(_4498_),
    .C(_4213_),
    .Y(_4499_)
);

INVX2 _15021_ (
    .A(_4499_),
    .Y(_4501_)
);

NOR2X1 _15022_ (
    .A(_5420__bF$buf0),
    .B(_2465__bF$buf2),
    .Y(_4502_)
);

AND2X2 _15023_ (
    .A(breg_7_bF$buf2),
    .B(areg_16_bF$buf1),
    .Y(_4503_)
);

AND2X2 _15024_ (
    .A(breg_6_bF$buf4),
    .B(areg_17_bF$buf1),
    .Y(_4504_)
);

NAND2X1 _15025_ (
    .A(_4503_),
    .B(_4504_),
    .Y(_4505_)
);

OAI21X1 _15026_ (
    .A(_5453__bF$buf5),
    .B(_2884__bF$buf1),
    .C(_4498_),
    .Y(_4506_)
);

NAND3X1 _15027_ (
    .A(_4502_),
    .B(_4506_),
    .C(_4505_),
    .Y(_4507_)
);

INVX1 _15028_ (
    .A(_4502_),
    .Y(_4508_)
);

OAI21X1 _15029_ (
    .A(_4116__bF$buf0),
    .B(_2669__bF$buf3),
    .C(_4504_),
    .Y(_4509_)
);

OAI21X1 _15030_ (
    .A(_5453__bF$buf4),
    .B(_2884__bF$buf0),
    .C(_4503_),
    .Y(_4510_)
);

NAND3X1 _15031_ (
    .A(_4509_),
    .B(_4510_),
    .C(_4508_),
    .Y(_4512_)
);

NAND2X1 _15032_ (
    .A(_4219_),
    .B(_4238_),
    .Y(_4513_)
);

OAI21X1 _15033_ (
    .A(_4236_),
    .B(_4239_),
    .C(_4513_),
    .Y(_4514_)
);

NAND3X1 _15034_ (
    .A(_4514_),
    .B(_4507_),
    .C(_4512_),
    .Y(_4515_)
);

AOI21X1 _15035_ (
    .A(_4509_),
    .B(_4510_),
    .C(_4508_),
    .Y(_4516_)
);

AOI21X1 _15036_ (
    .A(_4506_),
    .B(_4505_),
    .C(_4502_),
    .Y(_4517_)
);

INVX1 _15037_ (
    .A(_4239_),
    .Y(_4518_)
);

AOI22X1 _15038_ (
    .A(_4219_),
    .B(_4238_),
    .C(_4518_),
    .D(_4261_),
    .Y(_4519_)
);

OAI21X1 _15039_ (
    .A(_4516_),
    .B(_4517_),
    .C(_4519_),
    .Y(_4520_)
);

NAND3X1 _15040_ (
    .A(_4515_),
    .B(_4520_),
    .C(_4501_),
    .Y(_4521_)
);

NOR3X1 _15041_ (
    .A(_4517_),
    .B(_4519_),
    .C(_4516_),
    .Y(_4523_)
);

AOI21X1 _15042_ (
    .A(_4507_),
    .B(_4512_),
    .C(_4514_),
    .Y(_4524_)
);

OAI21X1 _15043_ (
    .A(_4523_),
    .B(_4524_),
    .C(_4499_),
    .Y(_4525_)
);

NAND2X1 _15044_ (
    .A(_4521_),
    .B(_4525_),
    .Y(_4526_)
);

AOI21X1 _15045_ (
    .A(_4252_),
    .B(_4249_),
    .C(_4242_),
    .Y(_4527_)
);

OAI21X1 _15046_ (
    .A(_4527_),
    .B(_4262_),
    .C(_4253_),
    .Y(_4528_)
);

NOR2X1 _15047_ (
    .A(_4258__bF$buf1),
    .B(_3146__bF$buf0),
    .Y(_4529_)
);

AND2X2 _15048_ (
    .A(breg_3_bF$buf1),
    .B(areg_19_bF$buf4),
    .Y(_4530_)
);

AND2X2 _15049_ (
    .A(breg_4_bF$buf5),
    .B(areg_20_bF$buf4),
    .Y(_4531_)
);

AOI22X1 _15050_ (
    .A(breg_3_bF$buf0),
    .B(areg_20_bF$buf3),
    .C(breg_4_bF$buf4),
    .D(areg_19_bF$buf3),
    .Y(_4532_)
);

AOI21X1 _15051_ (
    .A(_4530_),
    .B(_4531_),
    .C(_4532_),
    .Y(_4534_)
);

XOR2X1 _15052_ (
    .A(_4534_),
    .B(_4529_),
    .Y(_4535_)
);

OAI21X1 _15053_ (
    .A(_4243_),
    .B(_4247_),
    .C(_4246_),
    .Y(_4536_)
);

NAND2X1 _15054_ (
    .A(breg_2_bF$buf0),
    .B(areg_21_bF$buf0),
    .Y(_4537_)
);

INVX2 _15055_ (
    .A(_4537_),
    .Y(_4538_)
);

AND2X2 _15056_ (
    .A(breg_0_bF$buf0),
    .B(areg_23_bF$buf4),
    .Y(_4539_)
);

NAND2X1 _15057_ (
    .A(_4245_),
    .B(_4539_),
    .Y(_4540_)
);

INVX8 _15058_ (
    .A(areg_23_bF$buf3),
    .Y(_4541_)
);

OAI21X1 _15059_ (
    .A(_2551__bF$buf3),
    .B(_4541__bF$buf4),
    .C(_4250_),
    .Y(_4542_)
);

NAND3X1 _15060_ (
    .A(_4538_),
    .B(_4542_),
    .C(_4540_),
    .Y(_4543_)
);

NAND2X1 _15061_ (
    .A(breg_0_bF$buf6),
    .B(areg_23_bF$buf2),
    .Y(_4545_)
);

NOR2X1 _15062_ (
    .A(_4250_),
    .B(_4545_),
    .Y(_4546_)
);

NOR2X1 _15063_ (
    .A(_4245_),
    .B(_4539_),
    .Y(_4547_)
);

OAI21X1 _15064_ (
    .A(_4547_),
    .B(_4546_),
    .C(_4537_),
    .Y(_4548_)
);

NAND3X1 _15065_ (
    .A(_4536_),
    .B(_4543_),
    .C(_4548_),
    .Y(_4549_)
);

AOI21X1 _15066_ (
    .A(_4244_),
    .B(_4248_),
    .C(_4251_),
    .Y(_4550_)
);

INVX8 _15067_ (
    .A(areg_22_bF$buf1),
    .Y(_4551_)
);

OAI21X1 _15068_ (
    .A(_3220_),
    .B(_4551__bF$buf4),
    .C(_4539_),
    .Y(_4552_)
);

OAI21X1 _15069_ (
    .A(_2551__bF$buf2),
    .B(_4541__bF$buf3),
    .C(_4245_),
    .Y(_4553_)
);

AOI21X1 _15070_ (
    .A(_4552_),
    .B(_4553_),
    .C(_4537_),
    .Y(_4554_)
);

AOI21X1 _15071_ (
    .A(_4542_),
    .B(_4540_),
    .C(_4538_),
    .Y(_4556_)
);

OAI21X1 _15072_ (
    .A(_4554_),
    .B(_4556_),
    .C(_4550_),
    .Y(_4557_)
);

NAND3X1 _15073_ (
    .A(_4535_),
    .B(_4557_),
    .C(_4549_),
    .Y(_4558_)
);

XNOR2X1 _15074_ (
    .A(_4534_),
    .B(_4529_),
    .Y(_4559_)
);

OAI21X1 _15075_ (
    .A(_4554_),
    .B(_4556_),
    .C(_4536_),
    .Y(_4560_)
);

NAND3X1 _15076_ (
    .A(_4550_),
    .B(_4543_),
    .C(_4548_),
    .Y(_4561_)
);

NAND3X1 _15077_ (
    .A(_4559_),
    .B(_4560_),
    .C(_4561_),
    .Y(_4562_)
);

NAND3X1 _15078_ (
    .A(_4558_),
    .B(_4528_),
    .C(_4562_),
    .Y(_4563_)
);

NOR3X1 _15079_ (
    .A(_4255_),
    .B(_4254_),
    .C(_4256_),
    .Y(_4564_)
);

AOI21X1 _15080_ (
    .A(_4241_),
    .B(_4257_),
    .C(_4564_),
    .Y(_4565_)
);

AOI21X1 _15081_ (
    .A(_4560_),
    .B(_4561_),
    .C(_4559_),
    .Y(_4567_)
);

AOI21X1 _15082_ (
    .A(_4557_),
    .B(_4549_),
    .C(_4535_),
    .Y(_4568_)
);

OAI21X1 _15083_ (
    .A(_4567_),
    .B(_4568_),
    .C(_4565_),
    .Y(_4569_)
);

NAND3X1 _15084_ (
    .A(_4563_),
    .B(_4526_),
    .C(_4569_),
    .Y(_4570_)
);

NAND3X1 _15085_ (
    .A(_4499_),
    .B(_4515_),
    .C(_4520_),
    .Y(_4571_)
);

OAI21X1 _15086_ (
    .A(_4523_),
    .B(_4524_),
    .C(_4501_),
    .Y(_4572_)
);

NAND2X1 _15087_ (
    .A(_4571_),
    .B(_4572_),
    .Y(_4573_)
);

OAI21X1 _15088_ (
    .A(_4567_),
    .B(_4568_),
    .C(_4528_),
    .Y(_4574_)
);

NAND3X1 _15089_ (
    .A(_4558_),
    .B(_4562_),
    .C(_4565_),
    .Y(_4575_)
);

NAND3X1 _15090_ (
    .A(_4575_),
    .B(_4573_),
    .C(_4574_),
    .Y(_4576_)
);

NAND3X1 _15091_ (
    .A(_4497_),
    .B(_4570_),
    .C(_4576_),
    .Y(_4578_)
);

NOR3X1 _15092_ (
    .A(_4271_),
    .B(_4269_),
    .C(_4268_),
    .Y(_4579_)
);

AOI21X1 _15093_ (
    .A(_4233_),
    .B(_4272_),
    .C(_4579_),
    .Y(_4580_)
);

AOI21X1 _15094_ (
    .A(_4575_),
    .B(_4574_),
    .C(_4573_),
    .Y(_4581_)
);

AOI21X1 _15095_ (
    .A(_4563_),
    .B(_4569_),
    .C(_4526_),
    .Y(_4582_)
);

OAI21X1 _15096_ (
    .A(_4581_),
    .B(_4582_),
    .C(_4580_),
    .Y(_4583_)
);

NAND3X1 _15097_ (
    .A(_4578_),
    .B(_4583_),
    .C(_4495_),
    .Y(_4584_)
);

NAND3X1 _15098_ (
    .A(_4448_),
    .B(_4492_),
    .C(_4493_),
    .Y(_4585_)
);

OAI21X1 _15099_ (
    .A(_4488_),
    .B(_4484_),
    .C(_4491_),
    .Y(_4586_)
);

NAND2X1 _15100_ (
    .A(_4585_),
    .B(_4586_),
    .Y(_4587_)
);

OAI21X1 _15101_ (
    .A(_4581_),
    .B(_4582_),
    .C(_4497_),
    .Y(_4589_)
);

NAND3X1 _15102_ (
    .A(_4570_),
    .B(_4576_),
    .C(_4580_),
    .Y(_4590_)
);

NAND3X1 _15103_ (
    .A(_4590_),
    .B(_4589_),
    .C(_4587_),
    .Y(_4591_)
);

NAND3X1 _15104_ (
    .A(_4584_),
    .B(_4591_),
    .C(_4447_),
    .Y(_4592_)
);

NOR3X1 _15105_ (
    .A(_4284_),
    .B(_4285_),
    .C(_4283_),
    .Y(_4593_)
);

AOI21X1 _15106_ (
    .A(_4200_),
    .B(_4286_),
    .C(_4593_),
    .Y(_4594_)
);

AOI21X1 _15107_ (
    .A(_4590_),
    .B(_4589_),
    .C(_4587_),
    .Y(_4595_)
);

AOI21X1 _15108_ (
    .A(_4578_),
    .B(_4583_),
    .C(_4495_),
    .Y(_4596_)
);

OAI21X1 _15109_ (
    .A(_4595_),
    .B(_4596_),
    .C(_4594_),
    .Y(_4597_)
);

NAND3X1 _15110_ (
    .A(_4592_),
    .B(_4597_),
    .C(_4444_),
    .Y(_4598_)
);

NAND3X1 _15111_ (
    .A(_4440_),
    .B(_4433_),
    .C(_4438_),
    .Y(_4600_)
);

NAND3X1 _15112_ (
    .A(_4362_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4601_)
);

NAND2X1 _15113_ (
    .A(_4600_),
    .B(_4601_),
    .Y(_4602_)
);

OAI21X1 _15114_ (
    .A(_4595_),
    .B(_4596_),
    .C(_4447_),
    .Y(_4603_)
);

NAND3X1 _15115_ (
    .A(_4584_),
    .B(_4591_),
    .C(_4594_),
    .Y(_4604_)
);

NAND3X1 _15116_ (
    .A(_4604_),
    .B(_4603_),
    .C(_4602_),
    .Y(_4605_)
);

NAND3X1 _15117_ (
    .A(_4598_),
    .B(_4605_),
    .C(_4361_),
    .Y(_4606_)
);

NOR3X1 _15118_ (
    .A(_4298_),
    .B(_4299_),
    .C(_4297_),
    .Y(_4607_)
);

AOI21X1 _15119_ (
    .A(_4300_),
    .B(_4152_),
    .C(_4607_),
    .Y(_4608_)
);

AOI21X1 _15120_ (
    .A(_4604_),
    .B(_4603_),
    .C(_4602_),
    .Y(_4609_)
);

AOI21X1 _15121_ (
    .A(_4592_),
    .B(_4597_),
    .C(_4444_),
    .Y(_4611_)
);

OAI21X1 _15122_ (
    .A(_4609_),
    .B(_4611_),
    .C(_4608_),
    .Y(_4612_)
);

NAND3X1 _15123_ (
    .A(_4359_),
    .B(_4606_),
    .C(_4612_),
    .Y(_4613_)
);

XNOR2X1 _15124_ (
    .A(_4358_),
    .B(_4356_),
    .Y(_4614_)
);

OAI21X1 _15125_ (
    .A(_4609_),
    .B(_4611_),
    .C(_4361_),
    .Y(_4615_)
);

NAND3X1 _15126_ (
    .A(_4598_),
    .B(_4605_),
    .C(_4608_),
    .Y(_4616_)
);

NAND3X1 _15127_ (
    .A(_4614_),
    .B(_4616_),
    .C(_4615_),
    .Y(_4617_)
);

NAND3X1 _15128_ (
    .A(_4613_),
    .B(_4617_),
    .C(_4352_),
    .Y(_4618_)
);

NOR3X1 _15129_ (
    .A(_4312_),
    .B(_4313_),
    .C(_4311_),
    .Y(_4619_)
);

AOI21X1 _15130_ (
    .A(_4063_),
    .B(_4315_),
    .C(_4619_),
    .Y(_4620_)
);

AOI21X1 _15131_ (
    .A(_4616_),
    .B(_4615_),
    .C(_4614_),
    .Y(_4622_)
);

AOI21X1 _15132_ (
    .A(_4606_),
    .B(_4612_),
    .C(_4359_),
    .Y(_4623_)
);

OAI21X1 _15133_ (
    .A(_4622_),
    .B(_4623_),
    .C(_4620_),
    .Y(_4624_)
);

NAND3X1 _15134_ (
    .A(_4350_),
    .B(_4618_),
    .C(_4624_),
    .Y(_4625_)
);

OAI21X1 _15135_ (
    .A(_4622_),
    .B(_4623_),
    .C(_4352_),
    .Y(_4626_)
);

NAND3X1 _15136_ (
    .A(_4613_),
    .B(_4617_),
    .C(_4620_),
    .Y(_4627_)
);

NAND3X1 _15137_ (
    .A(_4349_),
    .B(_4627_),
    .C(_4626_),
    .Y(_4628_)
);

NAND3X1 _15138_ (
    .A(_4625_),
    .B(_4628_),
    .C(_4348_),
    .Y(_4629_)
);

NOR3X1 _15139_ (
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4630_)
);

AOI21X1 _15140_ (
    .A(_4058_),
    .B(_4326_),
    .C(_4630_),
    .Y(_4631_)
);

AOI21X1 _15141_ (
    .A(_4627_),
    .B(_4626_),
    .C(_4349_),
    .Y(_4633_)
);

AOI21X1 _15142_ (
    .A(_4618_),
    .B(_4624_),
    .C(_4350_),
    .Y(_4634_)
);

OAI21X1 _15143_ (
    .A(_4633_),
    .B(_4634_),
    .C(_4631_),
    .Y(_4635_)
);

NAND3X1 _15144_ (
    .A(_4339_),
    .B(_4629_),
    .C(_4635_),
    .Y(_4636_)
);

OAI21X1 _15145_ (
    .A(_4633_),
    .B(_4634_),
    .C(_4348_),
    .Y(_4637_)
);

NAND3X1 _15146_ (
    .A(_4625_),
    .B(_4628_),
    .C(_4631_),
    .Y(_4638_)
);

NAND3X1 _15147_ (
    .A(_4331_),
    .B(_4638_),
    .C(_4637_),
    .Y(_4639_)
);

NAND2X1 _15148_ (
    .A(_4636_),
    .B(_4639_),
    .Y(_4640_)
);

XNOR2X1 _15149_ (
    .A(_4345_),
    .B(_4640_),
    .Y(_0_[23])
);

NOR3X1 _15150_ (
    .A(_4342_),
    .B(_4640_),
    .C(_4054_),
    .Y(_4641_)
);

NAND2X1 _15151_ (
    .A(_3513_),
    .B(_4641_),
    .Y(_4643_)
);

NOR2X1 _15152_ (
    .A(_4342_),
    .B(_4640_),
    .Y(_4644_)
);

OAI21X1 _15153_ (
    .A(_4640_),
    .B(_4335_),
    .C(_4636_),
    .Y(_4645_)
);

AOI21X1 _15154_ (
    .A(_4052_),
    .B(_4644_),
    .C(_4645_),
    .Y(_4646_)
);

NAND3X1 _15155_ (
    .A(_3509_),
    .B(_3515_),
    .C(_4641_),
    .Y(_4647_)
);

NAND3X1 _15156_ (
    .A(_4643_),
    .B(_4646_),
    .C(_4647_),
    .Y(_4648_)
);

NOR3X1 _15157_ (
    .A(_4633_),
    .B(_4634_),
    .C(_4631_),
    .Y(_4649_)
);

AOI21X1 _15158_ (
    .A(_4613_),
    .B(_4617_),
    .C(_4352_),
    .Y(_4650_)
);

OAI21X1 _15159_ (
    .A(_4650_),
    .B(_4349_),
    .C(_4618_),
    .Y(_4651_)
);

NAND2X1 _15160_ (
    .A(_4356_),
    .B(_4358_),
    .Y(_4652_)
);

INVX2 _15161_ (
    .A(_4652_),
    .Y(_4654_)
);

AOI21X1 _15162_ (
    .A(_4598_),
    .B(_4605_),
    .C(_4361_),
    .Y(_4655_)
);

OAI21X1 _15163_ (
    .A(_4655_),
    .B(_4614_),
    .C(_4606_),
    .Y(_4656_)
);

OAI21X1 _15164_ (
    .A(_4367_),
    .B(_4385_),
    .C(_4384_),
    .Y(_4657_)
);

NAND2X1 _15165_ (
    .A(areg[0]),
    .B(breg_24_bF$buf5),
    .Y(_4658_)
);

INVX1 _15166_ (
    .A(_4658_),
    .Y(_4659_)
);

NAND3X1 _15167_ (
    .A(areg[0]),
    .B(breg_23_bF$buf2),
    .C(_4365_),
    .Y(_4660_)
);

OAI21X1 _15168_ (
    .A(_4068_),
    .B(_4364_),
    .C(_4660_),
    .Y(_4661_)
);

AND2X2 _15169_ (
    .A(_4661_),
    .B(_4659_),
    .Y(_4662_)
);

NOR2X1 _15170_ (
    .A(_4659_),
    .B(_4661_),
    .Y(_4663_)
);

NOR2X1 _15171_ (
    .A(_4663_),
    .B(_4662_),
    .Y(_4665_)
);

XNOR2X1 _15172_ (
    .A(_4665_),
    .B(_4657_),
    .Y(_4666_)
);

OAI21X1 _15173_ (
    .A(_4353_),
    .B(_4095_),
    .C(_4666_),
    .Y(_4667_)
);

INVX1 _15174_ (
    .A(_4354_),
    .Y(_4668_)
);

NOR2X1 _15175_ (
    .A(_4668_),
    .B(_4666_),
    .Y(_4669_)
);

INVX1 _15176_ (
    .A(_4669_),
    .Y(_4670_)
);

NAND2X1 _15177_ (
    .A(_4667_),
    .B(_4670_),
    .Y(_4671_)
);

NAND2X1 _15178_ (
    .A(_4433_),
    .B(_4600_),
    .Y(_4672_)
);

XNOR2X1 _15179_ (
    .A(_4672_),
    .B(_4671_),
    .Y(_4673_)
);

AOI21X1 _15180_ (
    .A(_4584_),
    .B(_4591_),
    .C(_4447_),
    .Y(_4674_)
);

OAI21X1 _15181_ (
    .A(_4602_),
    .B(_4674_),
    .C(_4592_),
    .Y(_4676_)
);

NAND2X1 _15182_ (
    .A(_4419_),
    .B(_4427_),
    .Y(_4677_)
);

NAND2X1 _15183_ (
    .A(areg_1_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_4678_)
);

NAND2X1 _15184_ (
    .A(areg_3_bF$buf0),
    .B(breg_22_bF$buf2),
    .Y(_4679_)
);

NOR2X1 _15185_ (
    .A(_4364_),
    .B(_4679_),
    .Y(_4680_)
);

AOI22X1 _15186_ (
    .A(areg_3_bF$buf4),
    .B(breg_21_bF$buf2),
    .C(areg_2_bF$buf2),
    .D(breg_22_bF$buf1),
    .Y(_4681_)
);

NOR2X1 _15187_ (
    .A(_4681_),
    .B(_4680_),
    .Y(_4682_)
);

XNOR2X1 _15188_ (
    .A(_4682_),
    .B(_4678_),
    .Y(_4683_)
);

AOI21X1 _15189_ (
    .A(_4375_),
    .B(_4377_),
    .C(_4372_),
    .Y(_4684_)
);

INVX2 _15190_ (
    .A(_4684_),
    .Y(_4685_)
);

NOR2X1 _15191_ (
    .A(_2562__bF$buf0),
    .B(_3526_),
    .Y(_4687_)
);

NAND2X1 _15192_ (
    .A(areg_5_bF$buf3),
    .B(breg_19_bF$buf0),
    .Y(_4688_)
);

NAND2X1 _15193_ (
    .A(areg_6_bF$buf3),
    .B(breg_18_bF$buf5),
    .Y(_4689_)
);

NOR2X1 _15194_ (
    .A(_4688_),
    .B(_4689_),
    .Y(_4690_)
);

INVX1 _15195_ (
    .A(_4690_),
    .Y(_4691_)
);

OAI21X1 _15196_ (
    .A(_3646__bF$buf3),
    .B(_3529__bF$buf1),
    .C(_4688_),
    .Y(_4692_)
);

NAND3X1 _15197_ (
    .A(_4687_),
    .B(_4692_),
    .C(_4691_),
    .Y(_4693_)
);

NAND2X1 _15198_ (
    .A(areg_6_bF$buf2),
    .B(breg_19_bF$buf5),
    .Y(_4694_)
);

OAI21X1 _15199_ (
    .A(_4371_),
    .B(_4694_),
    .C(_4692_),
    .Y(_4695_)
);

OAI21X1 _15200_ (
    .A(_2562__bF$buf4),
    .B(_3526_),
    .C(_4695_),
    .Y(_4696_)
);

NAND3X1 _15201_ (
    .A(_4693_),
    .B(_4696_),
    .C(_4685_),
    .Y(_4698_)
);

INVX1 _15202_ (
    .A(_4687_),
    .Y(_4699_)
);

NOR2X1 _15203_ (
    .A(_4699_),
    .B(_4695_),
    .Y(_4700_)
);

AOI21X1 _15204_ (
    .A(_4692_),
    .B(_4691_),
    .C(_4687_),
    .Y(_4701_)
);

OAI21X1 _15205_ (
    .A(_4700_),
    .B(_4701_),
    .C(_4684_),
    .Y(_4702_)
);

NAND3X1 _15206_ (
    .A(_4683_),
    .B(_4698_),
    .C(_4702_),
    .Y(_4703_)
);

XOR2X1 _15207_ (
    .A(_4682_),
    .B(_4678_),
    .Y(_4704_)
);

OAI21X1 _15208_ (
    .A(_4700_),
    .B(_4701_),
    .C(_4685_),
    .Y(_4705_)
);

NAND3X1 _15209_ (
    .A(_4684_),
    .B(_4693_),
    .C(_4696_),
    .Y(_4706_)
);

NAND3X1 _15210_ (
    .A(_4704_),
    .B(_4706_),
    .C(_4705_),
    .Y(_4707_)
);

AND2X2 _15211_ (
    .A(_4703_),
    .B(_4707_),
    .Y(_4709_)
);

OAI21X1 _15212_ (
    .A(_4415_),
    .B(_4417_),
    .C(_4409_),
    .Y(_4710_)
);

OAI21X1 _15213_ (
    .A(_4403_),
    .B(_4392_),
    .C(_4396_),
    .Y(_4711_)
);

NAND2X1 _15214_ (
    .A(areg_7_bF$buf0),
    .B(breg_17_bF$buf1),
    .Y(_4712_)
);

INVX1 _15215_ (
    .A(_4712_),
    .Y(_4713_)
);

AND2X2 _15216_ (
    .A(areg_8_bF$buf4),
    .B(breg_16_bF$buf0),
    .Y(_4714_)
);

AND2X2 _15217_ (
    .A(areg_9_bF$buf4),
    .B(breg_15_bF$buf1),
    .Y(_4715_)
);

NAND2X1 _15218_ (
    .A(_4714_),
    .B(_4715_),
    .Y(_4716_)
);

OAI22X1 _15219_ (
    .A(_5190__bF$buf3),
    .B(_2560__bF$buf1),
    .C(_6582__bF$buf0),
    .D(_2362__bF$buf1),
    .Y(_4717_)
);

NAND3X1 _15220_ (
    .A(_4713_),
    .B(_4717_),
    .C(_4716_),
    .Y(_4718_)
);

OAI21X1 _15221_ (
    .A(_5190__bF$buf2),
    .B(_2560__bF$buf0),
    .C(_4715_),
    .Y(_4720_)
);

OAI21X1 _15222_ (
    .A(_6582__bF$buf3),
    .B(_2362__bF$buf0),
    .C(_4714_),
    .Y(_4721_)
);

NAND3X1 _15223_ (
    .A(_4712_),
    .B(_4720_),
    .C(_4721_),
    .Y(_4722_)
);

NAND2X1 _15224_ (
    .A(areg_11_bF$buf0),
    .B(breg_13_bF$buf3),
    .Y(_4723_)
);

AND2X2 _15225_ (
    .A(_4450_),
    .B(_4451_),
    .Y(_4724_)
);

OAI22X1 _15226_ (
    .A(_4159_),
    .B(_4723_),
    .C(_4724_),
    .D(_4449_),
    .Y(_4725_)
);

NAND3X1 _15227_ (
    .A(_4718_),
    .B(_4722_),
    .C(_4725_),
    .Y(_4726_)
);

AOI21X1 _15228_ (
    .A(_4720_),
    .B(_4721_),
    .C(_4712_),
    .Y(_4727_)
);

AOI21X1 _15229_ (
    .A(_4717_),
    .B(_4716_),
    .C(_4713_),
    .Y(_4728_)
);

NOR2X1 _15230_ (
    .A(_4450_),
    .B(_4451_),
    .Y(_4729_)
);

OAI21X1 _15231_ (
    .A(_9104__bF$buf1),
    .B(_2586__bF$buf2),
    .C(_4450_),
    .Y(_4731_)
);

AOI21X1 _15232_ (
    .A(_4476_),
    .B(_4731_),
    .C(_4729_),
    .Y(_4732_)
);

OAI21X1 _15233_ (
    .A(_4727_),
    .B(_4728_),
    .C(_4732_),
    .Y(_4733_)
);

NAND3X1 _15234_ (
    .A(_4711_),
    .B(_4726_),
    .C(_4733_),
    .Y(_4734_)
);

INVX2 _15235_ (
    .A(_4711_),
    .Y(_4735_)
);

NOR3X1 _15236_ (
    .A(_4728_),
    .B(_4732_),
    .C(_4727_),
    .Y(_4736_)
);

AOI21X1 _15237_ (
    .A(_4718_),
    .B(_4722_),
    .C(_4725_),
    .Y(_4737_)
);

OAI21X1 _15238_ (
    .A(_4736_),
    .B(_4737_),
    .C(_4735_),
    .Y(_4738_)
);

NAND3X1 _15239_ (
    .A(_4734_),
    .B(_4738_),
    .C(_4710_),
    .Y(_4739_)
);

AOI21X1 _15240_ (
    .A(_4391_),
    .B(_4413_),
    .C(_4416_),
    .Y(_4740_)
);

NAND3X1 _15241_ (
    .A(_4732_),
    .B(_4718_),
    .C(_4722_),
    .Y(_4742_)
);

OAI21X1 _15242_ (
    .A(_4727_),
    .B(_4728_),
    .C(_4725_),
    .Y(_4743_)
);

AOI21X1 _15243_ (
    .A(_4742_),
    .B(_4743_),
    .C(_4735_),
    .Y(_4744_)
);

AOI21X1 _15244_ (
    .A(_4726_),
    .B(_4733_),
    .C(_4711_),
    .Y(_4745_)
);

OAI21X1 _15245_ (
    .A(_4744_),
    .B(_4745_),
    .C(_4740_),
    .Y(_4746_)
);

NAND3X1 _15246_ (
    .A(_4739_),
    .B(_4746_),
    .C(_4709_),
    .Y(_4747_)
);

NAND2X1 _15247_ (
    .A(_4703_),
    .B(_4707_),
    .Y(_4748_)
);

OAI21X1 _15248_ (
    .A(_4744_),
    .B(_4745_),
    .C(_4710_),
    .Y(_4749_)
);

NAND3X1 _15249_ (
    .A(_4734_),
    .B(_4738_),
    .C(_4740_),
    .Y(_4750_)
);

NAND3X1 _15250_ (
    .A(_4749_),
    .B(_4750_),
    .C(_4748_),
    .Y(_4751_)
);

OAI21X1 _15251_ (
    .A(_4484_),
    .B(_4491_),
    .C(_4493_),
    .Y(_4753_)
);

AOI21X1 _15252_ (
    .A(_4751_),
    .B(_4747_),
    .C(_4753_),
    .Y(_4754_)
);

AOI21X1 _15253_ (
    .A(_4749_),
    .B(_4750_),
    .C(_4748_),
    .Y(_4755_)
);

AOI21X1 _15254_ (
    .A(_4739_),
    .B(_4746_),
    .C(_4709_),
    .Y(_4756_)
);

AOI21X1 _15255_ (
    .A(_4448_),
    .B(_4492_),
    .C(_4488_),
    .Y(_4757_)
);

NOR3X1 _15256_ (
    .A(_4757_),
    .B(_4755_),
    .C(_4756_),
    .Y(_4758_)
);

OAI21X1 _15257_ (
    .A(_4758_),
    .B(_4754_),
    .C(_4677_),
    .Y(_4759_)
);

NOR2X1 _15258_ (
    .A(_4424_),
    .B(_4425_),
    .Y(_4760_)
);

AOI21X1 _15259_ (
    .A(_4389_),
    .B(_4760_),
    .C(_4435_),
    .Y(_4761_)
);

OAI21X1 _15260_ (
    .A(_4756_),
    .B(_4755_),
    .C(_4757_),
    .Y(_4762_)
);

NAND3X1 _15261_ (
    .A(_4751_),
    .B(_4753_),
    .C(_4747_),
    .Y(_4764_)
);

NAND3X1 _15262_ (
    .A(_4761_),
    .B(_4764_),
    .C(_4762_),
    .Y(_4765_)
);

NAND2X1 _15263_ (
    .A(_4765_),
    .B(_4759_),
    .Y(_4766_)
);

AOI21X1 _15264_ (
    .A(_4570_),
    .B(_4576_),
    .C(_4497_),
    .Y(_4767_)
);

OAI21X1 _15265_ (
    .A(_4587_),
    .B(_4767_),
    .C(_4578_),
    .Y(_4768_)
);

NAND2X1 _15266_ (
    .A(_4468_),
    .B(_4475_),
    .Y(_4769_)
);

NAND2X1 _15267_ (
    .A(areg_10_bF$buf4),
    .B(breg_14_bF$buf2),
    .Y(_4770_)
);

NAND2X1 _15268_ (
    .A(areg_12_bF$buf0),
    .B(breg_12_bF$buf1),
    .Y(_4771_)
);

XOR2X1 _15269_ (
    .A(_4723_),
    .B(_4771_),
    .Y(_4772_)
);

XNOR2X1 _15270_ (
    .A(_4772_),
    .B(_4770_),
    .Y(_4773_)
);

OAI21X1 _15271_ (
    .A(_4465_),
    .B(_4455_),
    .C(_4459_),
    .Y(_4775_)
);

NAND2X1 _15272_ (
    .A(breg_11_bF$buf3),
    .B(areg_13_bF$buf3),
    .Y(_4776_)
);

INVX2 _15273_ (
    .A(_4776_),
    .Y(_4777_)
);

AND2X2 _15274_ (
    .A(breg_10_bF$buf4),
    .B(areg_14_bF$buf2),
    .Y(_4778_)
);

AND2X2 _15275_ (
    .A(breg_9_bF$buf0),
    .B(areg_15_bF$buf1),
    .Y(_4779_)
);

NAND2X1 _15276_ (
    .A(_4778_),
    .B(_4779_),
    .Y(_4780_)
);

OAI22X1 _15277_ (
    .A(_6044__bF$buf0),
    .B(_2465__bF$buf1),
    .C(_7217__bF$buf1),
    .D(_2287__bF$buf3),
    .Y(_4781_)
);

NAND3X1 _15278_ (
    .A(_4777_),
    .B(_4781_),
    .C(_4780_),
    .Y(_4782_)
);

NAND2X1 _15279_ (
    .A(breg_10_bF$buf3),
    .B(areg_15_bF$buf0),
    .Y(_4783_)
);

NOR2X1 _15280_ (
    .A(_4463_),
    .B(_4783_),
    .Y(_4784_)
);

NOR2X1 _15281_ (
    .A(_4778_),
    .B(_4779_),
    .Y(_4786_)
);

OAI21X1 _15282_ (
    .A(_4786_),
    .B(_4784_),
    .C(_4776_),
    .Y(_4787_)
);

NAND3X1 _15283_ (
    .A(_4782_),
    .B(_4775_),
    .C(_4787_),
    .Y(_4788_)
);

AOI21X1 _15284_ (
    .A(_4456_),
    .B(_4461_),
    .C(_4464_),
    .Y(_4789_)
);

NOR3X1 _15285_ (
    .A(_4776_),
    .B(_4784_),
    .C(_4786_),
    .Y(_4790_)
);

AOI21X1 _15286_ (
    .A(_4781_),
    .B(_4780_),
    .C(_4777_),
    .Y(_4791_)
);

OAI21X1 _15287_ (
    .A(_4790_),
    .B(_4791_),
    .C(_4789_),
    .Y(_4792_)
);

NAND3X1 _15288_ (
    .A(_4788_),
    .B(_4792_),
    .C(_4773_),
    .Y(_4793_)
);

INVX2 _15289_ (
    .A(_4770_),
    .Y(_4794_)
);

XNOR2X1 _15290_ (
    .A(_4772_),
    .B(_4794_),
    .Y(_4795_)
);

OAI21X1 _15291_ (
    .A(_4790_),
    .B(_4791_),
    .C(_4775_),
    .Y(_4797_)
);

NAND3X1 _15292_ (
    .A(_4789_),
    .B(_4782_),
    .C(_4787_),
    .Y(_4798_)
);

NAND3X1 _15293_ (
    .A(_4798_),
    .B(_4797_),
    .C(_4795_),
    .Y(_4799_)
);

OAI21X1 _15294_ (
    .A(_4501_),
    .B(_4524_),
    .C(_4515_),
    .Y(_4800_)
);

AOI21X1 _15295_ (
    .A(_4793_),
    .B(_4799_),
    .C(_4800_),
    .Y(_4801_)
);

AOI21X1 _15296_ (
    .A(_4798_),
    .B(_4797_),
    .C(_4795_),
    .Y(_4802_)
);

AOI21X1 _15297_ (
    .A(_4788_),
    .B(_4792_),
    .C(_4773_),
    .Y(_4803_)
);

AOI21X1 _15298_ (
    .A(_4499_),
    .B(_4520_),
    .C(_4523_),
    .Y(_4804_)
);

NOR3X1 _15299_ (
    .A(_4803_),
    .B(_4804_),
    .C(_4802_),
    .Y(_4805_)
);

OAI21X1 _15300_ (
    .A(_4805_),
    .B(_4801_),
    .C(_4769_),
    .Y(_4806_)
);

AND2X2 _15301_ (
    .A(_4475_),
    .B(_4468_),
    .Y(_4808_)
);

OAI21X1 _15302_ (
    .A(_4802_),
    .B(_4803_),
    .C(_4804_),
    .Y(_4809_)
);

NAND3X1 _15303_ (
    .A(_4793_),
    .B(_4799_),
    .C(_4800_),
    .Y(_4810_)
);

NAND3X1 _15304_ (
    .A(_4808_),
    .B(_4810_),
    .C(_4809_),
    .Y(_4811_)
);

NAND2X1 _15305_ (
    .A(_4811_),
    .B(_4806_),
    .Y(_4812_)
);

AOI21X1 _15306_ (
    .A(_4558_),
    .B(_4562_),
    .C(_4528_),
    .Y(_4813_)
);

OAI21X1 _15307_ (
    .A(_4573_),
    .B(_4813_),
    .C(_4563_),
    .Y(_4814_)
);

INVX1 _15308_ (
    .A(_4504_),
    .Y(_4815_)
);

OAI21X1 _15309_ (
    .A(_4498_),
    .B(_4815_),
    .C(_4507_),
    .Y(_4816_)
);

INVX2 _15310_ (
    .A(_4816_),
    .Y(_4817_)
);

NOR2X1 _15311_ (
    .A(_5420__bF$buf3),
    .B(_2669__bF$buf2),
    .Y(_4819_)
);

AND2X2 _15312_ (
    .A(breg_7_bF$buf1),
    .B(areg_17_bF$buf0),
    .Y(_4820_)
);

AND2X2 _15313_ (
    .A(breg_6_bF$buf3),
    .B(areg_18_bF$buf1),
    .Y(_4821_)
);

NAND2X1 _15314_ (
    .A(_4820_),
    .B(_4821_),
    .Y(_4822_)
);

OAI22X1 _15315_ (
    .A(_5453__bF$buf3),
    .B(_3146__bF$buf3),
    .C(_4116__bF$buf4),
    .D(_2884__bF$buf3),
    .Y(_4823_)
);

NAND3X1 _15316_ (
    .A(_4819_),
    .B(_4823_),
    .C(_4822_),
    .Y(_4824_)
);

INVX1 _15317_ (
    .A(_4819_),
    .Y(_4825_)
);

OAI21X1 _15318_ (
    .A(_4116__bF$buf3),
    .B(_2884__bF$buf2),
    .C(_4821_),
    .Y(_4826_)
);

OAI21X1 _15319_ (
    .A(_5453__bF$buf2),
    .B(_3146__bF$buf2),
    .C(_4820_),
    .Y(_4827_)
);

NAND3X1 _15320_ (
    .A(_4826_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4828_)
);

INVX1 _15321_ (
    .A(_4529_),
    .Y(_4830_)
);

AND2X2 _15322_ (
    .A(breg_3_bF$buf5),
    .B(areg_20_bF$buf2),
    .Y(_4831_)
);

NAND2X1 _15323_ (
    .A(_4238_),
    .B(_4831_),
    .Y(_4832_)
);

OAI21X1 _15324_ (
    .A(_4830_),
    .B(_4532_),
    .C(_4832_),
    .Y(_4833_)
);

NAND3X1 _15325_ (
    .A(_4824_),
    .B(_4828_),
    .C(_4833_),
    .Y(_4834_)
);

AOI21X1 _15326_ (
    .A(_4826_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4835_)
);

AOI21X1 _15327_ (
    .A(_4823_),
    .B(_4822_),
    .C(_4819_),
    .Y(_4836_)
);

INVX1 _15328_ (
    .A(_4532_),
    .Y(_4837_)
);

AOI22X1 _15329_ (
    .A(_4530_),
    .B(_4531_),
    .C(_4837_),
    .D(_4529_),
    .Y(_4838_)
);

OAI21X1 _15330_ (
    .A(_4835_),
    .B(_4836_),
    .C(_4838_),
    .Y(_4839_)
);

NAND3X1 _15331_ (
    .A(_4834_),
    .B(_4839_),
    .C(_4817_),
    .Y(_4841_)
);

NOR3X1 _15332_ (
    .A(_4836_),
    .B(_4838_),
    .C(_4835_),
    .Y(_4842_)
);

AOI21X1 _15333_ (
    .A(_4824_),
    .B(_4828_),
    .C(_4833_),
    .Y(_4843_)
);

OAI21X1 _15334_ (
    .A(_4842_),
    .B(_4843_),
    .C(_4816_),
    .Y(_4844_)
);

NAND2X1 _15335_ (
    .A(_4841_),
    .B(_4844_),
    .Y(_4845_)
);

AOI21X1 _15336_ (
    .A(_4543_),
    .B(_4548_),
    .C(_4536_),
    .Y(_4846_)
);

OAI21X1 _15337_ (
    .A(_4846_),
    .B(_4559_),
    .C(_4549_),
    .Y(_4847_)
);

NAND2X1 _15338_ (
    .A(breg_5_bF$buf0),
    .B(areg_19_bF$buf2),
    .Y(_4848_)
);

AND2X2 _15339_ (
    .A(breg_4_bF$buf3),
    .B(areg_21_bF$buf4),
    .Y(_4849_)
);

AOI22X1 _15340_ (
    .A(breg_3_bF$buf4),
    .B(areg_21_bF$buf3),
    .C(breg_4_bF$buf2),
    .D(areg_20_bF$buf1),
    .Y(_4850_)
);

AOI21X1 _15341_ (
    .A(_4831_),
    .B(_4849_),
    .C(_4850_),
    .Y(_4852_)
);

XNOR2X1 _15342_ (
    .A(_4852_),
    .B(_4848_),
    .Y(_4853_)
);

OAI21X1 _15343_ (
    .A(_4547_),
    .B(_4537_),
    .C(_4540_),
    .Y(_4854_)
);

NAND2X1 _15344_ (
    .A(breg_2_bF$buf4),
    .B(areg_22_bF$buf0),
    .Y(_4855_)
);

INVX2 _15345_ (
    .A(_4855_),
    .Y(_4856_)
);

AND2X2 _15346_ (
    .A(breg_1_bF$buf6),
    .B(areg_24_bF$buf4),
    .Y(_4857_)
);

NAND2X1 _15347_ (
    .A(_4539_),
    .B(_4857_),
    .Y(_4858_)
);

AOI22X1 _15348_ (
    .A(breg_0_bF$buf5),
    .B(areg_24_bF$buf3),
    .C(breg_1_bF$buf5),
    .D(areg_23_bF$buf1),
    .Y(_4859_)
);

INVX2 _15349_ (
    .A(_4859_),
    .Y(_4860_)
);

NAND3X1 _15350_ (
    .A(_4856_),
    .B(_4860_),
    .C(_4858_),
    .Y(_4861_)
);

NAND2X1 _15351_ (
    .A(breg_1_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_4863_)
);

NOR2X1 _15352_ (
    .A(_4545_),
    .B(_4863_),
    .Y(_4864_)
);

OAI21X1 _15353_ (
    .A(_4864_),
    .B(_4859_),
    .C(_4855_),
    .Y(_4865_)
);

NAND3X1 _15354_ (
    .A(_4865_),
    .B(_4861_),
    .C(_4854_),
    .Y(_4866_)
);

AOI21X1 _15355_ (
    .A(_4538_),
    .B(_4542_),
    .C(_4546_),
    .Y(_4867_)
);

NOR3X1 _15356_ (
    .A(_4855_),
    .B(_4859_),
    .C(_4864_),
    .Y(_4868_)
);

AOI21X1 _15357_ (
    .A(_4860_),
    .B(_4858_),
    .C(_4856_),
    .Y(_4869_)
);

OAI21X1 _15358_ (
    .A(_4869_),
    .B(_4868_),
    .C(_4867_),
    .Y(_4870_)
);

NAND3X1 _15359_ (
    .A(_4853_),
    .B(_4870_),
    .C(_4866_),
    .Y(_4871_)
);

INVX2 _15360_ (
    .A(_4848_),
    .Y(_4872_)
);

XNOR2X1 _15361_ (
    .A(_4852_),
    .B(_4872_),
    .Y(_4874_)
);

OAI21X1 _15362_ (
    .A(_4869_),
    .B(_4868_),
    .C(_4854_),
    .Y(_4875_)
);

NAND3X1 _15363_ (
    .A(_4867_),
    .B(_4865_),
    .C(_4861_),
    .Y(_4876_)
);

NAND3X1 _15364_ (
    .A(_4874_),
    .B(_4876_),
    .C(_4875_),
    .Y(_4877_)
);

NAND3X1 _15365_ (
    .A(_4871_),
    .B(_4877_),
    .C(_4847_),
    .Y(_4878_)
);

NOR3X1 _15366_ (
    .A(_4556_),
    .B(_4550_),
    .C(_4554_),
    .Y(_4879_)
);

AOI21X1 _15367_ (
    .A(_4535_),
    .B(_4557_),
    .C(_4879_),
    .Y(_4880_)
);

AOI21X1 _15368_ (
    .A(_4876_),
    .B(_4875_),
    .C(_4874_),
    .Y(_4881_)
);

AOI21X1 _15369_ (
    .A(_4870_),
    .B(_4866_),
    .C(_4853_),
    .Y(_4882_)
);

OAI21X1 _15370_ (
    .A(_4882_),
    .B(_4881_),
    .C(_4880_),
    .Y(_4883_)
);

NAND3X1 _15371_ (
    .A(_4878_),
    .B(_4883_),
    .C(_4845_),
    .Y(_4885_)
);

NAND3X1 _15372_ (
    .A(_4816_),
    .B(_4839_),
    .C(_4834_),
    .Y(_4886_)
);

OAI21X1 _15373_ (
    .A(_4842_),
    .B(_4843_),
    .C(_4817_),
    .Y(_4887_)
);

NAND2X1 _15374_ (
    .A(_4886_),
    .B(_4887_),
    .Y(_4888_)
);

OAI21X1 _15375_ (
    .A(_4882_),
    .B(_4881_),
    .C(_4847_),
    .Y(_4889_)
);

NAND3X1 _15376_ (
    .A(_4871_),
    .B(_4877_),
    .C(_4880_),
    .Y(_4890_)
);

NAND3X1 _15377_ (
    .A(_4890_),
    .B(_4888_),
    .C(_4889_),
    .Y(_4891_)
);

NAND3X1 _15378_ (
    .A(_4885_),
    .B(_4814_),
    .C(_4891_),
    .Y(_4892_)
);

NOR3X1 _15379_ (
    .A(_4567_),
    .B(_4568_),
    .C(_4565_),
    .Y(_4893_)
);

AOI21X1 _15380_ (
    .A(_4526_),
    .B(_4569_),
    .C(_4893_),
    .Y(_4894_)
);

AOI21X1 _15381_ (
    .A(_4890_),
    .B(_4889_),
    .C(_4888_),
    .Y(_4896_)
);

AOI21X1 _15382_ (
    .A(_4878_),
    .B(_4883_),
    .C(_4845_),
    .Y(_4897_)
);

OAI21X1 _15383_ (
    .A(_4896_),
    .B(_4897_),
    .C(_4894_),
    .Y(_4898_)
);

NAND3X1 _15384_ (
    .A(_4892_),
    .B(_4898_),
    .C(_4812_),
    .Y(_4899_)
);

NAND3X1 _15385_ (
    .A(_4769_),
    .B(_4810_),
    .C(_4809_),
    .Y(_4900_)
);

OAI21X1 _15386_ (
    .A(_4805_),
    .B(_4801_),
    .C(_4808_),
    .Y(_4901_)
);

NAND2X1 _15387_ (
    .A(_4900_),
    .B(_4901_),
    .Y(_4902_)
);

NOR3X1 _15388_ (
    .A(_4896_),
    .B(_4897_),
    .C(_4894_),
    .Y(_4903_)
);

AOI21X1 _15389_ (
    .A(_4885_),
    .B(_4891_),
    .C(_4814_),
    .Y(_4904_)
);

OAI21X1 _15390_ (
    .A(_4903_),
    .B(_4904_),
    .C(_4902_),
    .Y(_4905_)
);

NAND3X1 _15391_ (
    .A(_4768_),
    .B(_4899_),
    .C(_4905_),
    .Y(_4907_)
);

NOR3X1 _15392_ (
    .A(_4581_),
    .B(_4582_),
    .C(_4580_),
    .Y(_4908_)
);

AOI21X1 _15393_ (
    .A(_4495_),
    .B(_4583_),
    .C(_4908_),
    .Y(_4909_)
);

OAI21X1 _15394_ (
    .A(_4896_),
    .B(_4897_),
    .C(_4814_),
    .Y(_4910_)
);

NAND3X1 _15395_ (
    .A(_4885_),
    .B(_4891_),
    .C(_4894_),
    .Y(_4911_)
);

AOI21X1 _15396_ (
    .A(_4910_),
    .B(_4911_),
    .C(_4902_),
    .Y(_4912_)
);

AOI21X1 _15397_ (
    .A(_4892_),
    .B(_4898_),
    .C(_4812_),
    .Y(_4913_)
);

OAI21X1 _15398_ (
    .A(_4912_),
    .B(_4913_),
    .C(_4909_),
    .Y(_4914_)
);

NAND3X1 _15399_ (
    .A(_4914_),
    .B(_4907_),
    .C(_4766_),
    .Y(_4915_)
);

NAND3X1 _15400_ (
    .A(_4677_),
    .B(_4764_),
    .C(_4762_),
    .Y(_4916_)
);

OAI21X1 _15401_ (
    .A(_4758_),
    .B(_4754_),
    .C(_4761_),
    .Y(_4918_)
);

NAND2X1 _15402_ (
    .A(_4916_),
    .B(_4918_),
    .Y(_4919_)
);

NOR3X1 _15403_ (
    .A(_4912_),
    .B(_4913_),
    .C(_4909_),
    .Y(_4920_)
);

AOI21X1 _15404_ (
    .A(_4899_),
    .B(_4905_),
    .C(_4768_),
    .Y(_4921_)
);

OAI21X1 _15405_ (
    .A(_4920_),
    .B(_4921_),
    .C(_4919_),
    .Y(_4922_)
);

NAND3X1 _15406_ (
    .A(_4676_),
    .B(_4915_),
    .C(_4922_),
    .Y(_4923_)
);

NOR3X1 _15407_ (
    .A(_4595_),
    .B(_4596_),
    .C(_4594_),
    .Y(_4924_)
);

AOI21X1 _15408_ (
    .A(_4444_),
    .B(_4597_),
    .C(_4924_),
    .Y(_4925_)
);

OAI21X1 _15409_ (
    .A(_4912_),
    .B(_4913_),
    .C(_4768_),
    .Y(_4926_)
);

NAND3X1 _15410_ (
    .A(_4909_),
    .B(_4899_),
    .C(_4905_),
    .Y(_4927_)
);

AOI21X1 _15411_ (
    .A(_4926_),
    .B(_4927_),
    .C(_4919_),
    .Y(_4929_)
);

AOI21X1 _15412_ (
    .A(_4914_),
    .B(_4907_),
    .C(_4766_),
    .Y(_4930_)
);

OAI21X1 _15413_ (
    .A(_4929_),
    .B(_4930_),
    .C(_4925_),
    .Y(_4931_)
);

NAND3X1 _15414_ (
    .A(_4673_),
    .B(_4931_),
    .C(_4923_),
    .Y(_4932_)
);

XOR2X1 _15415_ (
    .A(_4672_),
    .B(_4671_),
    .Y(_4933_)
);

OAI21X1 _15416_ (
    .A(_4929_),
    .B(_4930_),
    .C(_4676_),
    .Y(_4934_)
);

NAND3X1 _15417_ (
    .A(_4925_),
    .B(_4915_),
    .C(_4922_),
    .Y(_4935_)
);

NAND3X1 _15418_ (
    .A(_4933_),
    .B(_4934_),
    .C(_4935_),
    .Y(_4936_)
);

NAND3X1 _15419_ (
    .A(_4656_),
    .B(_4932_),
    .C(_4936_),
    .Y(_4937_)
);

NOR3X1 _15420_ (
    .A(_4609_),
    .B(_4611_),
    .C(_4608_),
    .Y(_4938_)
);

AOI21X1 _15421_ (
    .A(_4359_),
    .B(_4612_),
    .C(_4938_),
    .Y(_4940_)
);

AOI21X1 _15422_ (
    .A(_4934_),
    .B(_4935_),
    .C(_4933_),
    .Y(_4941_)
);

AOI21X1 _15423_ (
    .A(_4931_),
    .B(_4923_),
    .C(_4673_),
    .Y(_4942_)
);

OAI21X1 _15424_ (
    .A(_4941_),
    .B(_4942_),
    .C(_4940_),
    .Y(_4943_)
);

NAND3X1 _15425_ (
    .A(_4654_),
    .B(_4937_),
    .C(_4943_),
    .Y(_4944_)
);

NOR3X1 _15426_ (
    .A(_4941_),
    .B(_4942_),
    .C(_4940_),
    .Y(_4945_)
);

AOI21X1 _15427_ (
    .A(_4932_),
    .B(_4936_),
    .C(_4656_),
    .Y(_4946_)
);

OAI21X1 _15428_ (
    .A(_4945_),
    .B(_4946_),
    .C(_4652_),
    .Y(_4947_)
);

NAND3X1 _15429_ (
    .A(_4651_),
    .B(_4944_),
    .C(_4947_),
    .Y(_4948_)
);

NOR3X1 _15430_ (
    .A(_4622_),
    .B(_4623_),
    .C(_4620_),
    .Y(_4949_)
);

AOI21X1 _15431_ (
    .A(_4350_),
    .B(_4624_),
    .C(_4949_),
    .Y(_4951_)
);

OAI21X1 _15432_ (
    .A(_4941_),
    .B(_4942_),
    .C(_4656_),
    .Y(_4952_)
);

NAND3X1 _15433_ (
    .A(_4932_),
    .B(_4936_),
    .C(_4940_),
    .Y(_4953_)
);

AOI21X1 _15434_ (
    .A(_4953_),
    .B(_4952_),
    .C(_4652_),
    .Y(_4954_)
);

AOI21X1 _15435_ (
    .A(_4937_),
    .B(_4943_),
    .C(_4654_),
    .Y(_4955_)
);

OAI21X1 _15436_ (
    .A(_4955_),
    .B(_4954_),
    .C(_4951_),
    .Y(_4956_)
);

NAND3X1 _15437_ (
    .A(_4956_),
    .B(_4948_),
    .C(_4649_),
    .Y(_4957_)
);

OAI21X1 _15438_ (
    .A(_4955_),
    .B(_4954_),
    .C(_4651_),
    .Y(_4958_)
);

NAND3X1 _15439_ (
    .A(_4951_),
    .B(_4944_),
    .C(_4947_),
    .Y(_4959_)
);

NAND3X1 _15440_ (
    .A(_4629_),
    .B(_4958_),
    .C(_4959_),
    .Y(_4960_)
);

NAND2X1 _15441_ (
    .A(_4960_),
    .B(_4957_),
    .Y(_4961_)
);

XNOR2X1 _15442_ (
    .A(_4648_),
    .B(_4961_),
    .Y(_0_[24])
);

INVX1 _15443_ (
    .A(_4648_),
    .Y(_4962_)
);

OAI21X1 _15444_ (
    .A(_4962_),
    .B(_4961_),
    .C(_4957_),
    .Y(_4963_)
);

NOR3X1 _15445_ (
    .A(_4954_),
    .B(_4955_),
    .C(_4951_),
    .Y(_4964_)
);

OAI21X1 _15446_ (
    .A(_4946_),
    .B(_4652_),
    .C(_4937_),
    .Y(_4965_)
);

INVX1 _15447_ (
    .A(_4672_),
    .Y(_4966_)
);

NOR2X1 _15448_ (
    .A(_4671_),
    .B(_4966_),
    .Y(_4967_)
);

AOI21X1 _15449_ (
    .A(_4915_),
    .B(_4922_),
    .C(_4676_),
    .Y(_4968_)
);

OAI21X1 _15450_ (
    .A(_4968_),
    .B(_4933_),
    .C(_4923_),
    .Y(_4969_)
);

NAND2X1 _15451_ (
    .A(_4657_),
    .B(_4665_),
    .Y(_4971_)
);

INVX2 _15452_ (
    .A(_4662_),
    .Y(_4972_)
);

NAND2X1 _15453_ (
    .A(areg_1_bF$buf2),
    .B(breg_25_bF$buf5),
    .Y(_4973_)
);

NOR2X1 _15454_ (
    .A(_4658_),
    .B(_4973_),
    .Y(_4974_)
);

AOI22X1 _15455_ (
    .A(areg_1_bF$buf1),
    .B(breg_24_bF$buf4),
    .C(areg[0]),
    .D(breg_25_bF$buf4),
    .Y(_4975_)
);

NOR2X1 _15456_ (
    .A(_4975_),
    .B(_4974_),
    .Y(_4976_)
);

OAI22X1 _15457_ (
    .A(_4364_),
    .B(_4679_),
    .C(_4681_),
    .D(_4678_),
    .Y(_4977_)
);

NOR2X1 _15458_ (
    .A(_4977_),
    .B(_4976_),
    .Y(_4978_)
);

NAND2X1 _15459_ (
    .A(_4977_),
    .B(_4976_),
    .Y(_4979_)
);

INVX2 _15460_ (
    .A(_4979_),
    .Y(_4980_)
);

NOR2X1 _15461_ (
    .A(_4978_),
    .B(_4980_),
    .Y(_4982_)
);

AOI21X1 _15462_ (
    .A(_4693_),
    .B(_4696_),
    .C(_4685_),
    .Y(_4983_)
);

OAI21X1 _15463_ (
    .A(_4983_),
    .B(_4704_),
    .C(_4698_),
    .Y(_4984_)
);

AND2X2 _15464_ (
    .A(_4984_),
    .B(_4982_),
    .Y(_4985_)
);

NOR2X1 _15465_ (
    .A(_4982_),
    .B(_4984_),
    .Y(_4986_)
);

NOR3X1 _15466_ (
    .A(_4986_),
    .B(_4972_),
    .C(_4985_),
    .Y(_4987_)
);

NAND2X1 _15467_ (
    .A(_4982_),
    .B(_4984_),
    .Y(_4988_)
);

OR2X2 _15468_ (
    .A(_4984_),
    .B(_4982_),
    .Y(_4989_)
);

AOI21X1 _15469_ (
    .A(_4988_),
    .B(_4989_),
    .C(_4662_),
    .Y(_4990_)
);

OAI21X1 _15470_ (
    .A(_4987_),
    .B(_4990_),
    .C(_4971_),
    .Y(_4991_)
);

AND2X2 _15471_ (
    .A(_4665_),
    .B(_4657_),
    .Y(_4993_)
);

NAND3X1 _15472_ (
    .A(_4662_),
    .B(_4988_),
    .C(_4989_),
    .Y(_4994_)
);

OAI21X1 _15473_ (
    .A(_4985_),
    .B(_4986_),
    .C(_4972_),
    .Y(_4995_)
);

NAND3X1 _15474_ (
    .A(_4993_),
    .B(_4995_),
    .C(_4994_),
    .Y(_4996_)
);

AND2X2 _15475_ (
    .A(_4991_),
    .B(_4996_),
    .Y(_4997_)
);

OAI21X1 _15476_ (
    .A(_4754_),
    .B(_4761_),
    .C(_4764_),
    .Y(_4998_)
);

NAND2X1 _15477_ (
    .A(_4998_),
    .B(_4997_),
    .Y(_4999_)
);

NAND2X1 _15478_ (
    .A(_4996_),
    .B(_4991_),
    .Y(_5000_)
);

NAND3X1 _15479_ (
    .A(_4764_),
    .B(_5000_),
    .C(_4916_),
    .Y(_5001_)
);

NAND3X1 _15480_ (
    .A(_4670_),
    .B(_5001_),
    .C(_4999_),
    .Y(_5002_)
);

OR2X2 _15481_ (
    .A(_4998_),
    .B(_5000_),
    .Y(_5004_)
);

NAND2X1 _15482_ (
    .A(_5000_),
    .B(_4998_),
    .Y(_5005_)
);

NAND3X1 _15483_ (
    .A(_4669_),
    .B(_5005_),
    .C(_5004_),
    .Y(_5006_)
);

NAND2X1 _15484_ (
    .A(_5002_),
    .B(_5006_),
    .Y(_5007_)
);

OAI21X1 _15485_ (
    .A(_4921_),
    .B(_4919_),
    .C(_4907_),
    .Y(_5008_)
);

NAND2X1 _15486_ (
    .A(_4739_),
    .B(_4747_),
    .Y(_5009_)
);

NAND2X1 _15487_ (
    .A(areg_2_bF$buf1),
    .B(breg_23_bF$buf0),
    .Y(_5010_)
);

INVX2 _15488_ (
    .A(_5010_),
    .Y(_5011_)
);

NAND2X1 _15489_ (
    .A(areg_4_bF$buf3),
    .B(breg_21_bF$buf1),
    .Y(_5012_)
);

NOR2X1 _15490_ (
    .A(_4679_),
    .B(_5012_),
    .Y(_5013_)
);

AND2X2 _15491_ (
    .A(_4679_),
    .B(_5012_),
    .Y(_5015_)
);

NOR2X1 _15492_ (
    .A(_5013_),
    .B(_5015_),
    .Y(_5016_)
);

XNOR2X1 _15493_ (
    .A(_5016_),
    .B(_5011_),
    .Y(_5017_)
);

AOI21X1 _15494_ (
    .A(_4687_),
    .B(_4692_),
    .C(_4690_),
    .Y(_5018_)
);

INVX2 _15495_ (
    .A(_5018_),
    .Y(_5019_)
);

NAND2X1 _15496_ (
    .A(areg_5_bF$buf2),
    .B(breg_20_bF$buf0),
    .Y(_5020_)
);

NAND2X1 _15497_ (
    .A(areg_7_bF$buf4),
    .B(breg_18_bF$buf4),
    .Y(_5021_)
);

NOR2X1 _15498_ (
    .A(_4694_),
    .B(_5021_),
    .Y(_5022_)
);

AND2X2 _15499_ (
    .A(_4694_),
    .B(_5021_),
    .Y(_5023_)
);

NOR3X1 _15500_ (
    .A(_5020_),
    .B(_5022_),
    .C(_5023_),
    .Y(_5024_)
);

INVX2 _15501_ (
    .A(_5020_),
    .Y(_5026_)
);

INVX2 _15502_ (
    .A(_5022_),
    .Y(_5027_)
);

OAI21X1 _15503_ (
    .A(_4434__bF$buf0),
    .B(_3529__bF$buf0),
    .C(_4694_),
    .Y(_5028_)
);

AOI21X1 _15504_ (
    .A(_5028_),
    .B(_5027_),
    .C(_5026_),
    .Y(_5029_)
);

OAI21X1 _15505_ (
    .A(_5029_),
    .B(_5024_),
    .C(_5019_),
    .Y(_5030_)
);

NAND3X1 _15506_ (
    .A(_5026_),
    .B(_5028_),
    .C(_5027_),
    .Y(_5031_)
);

OAI21X1 _15507_ (
    .A(_5023_),
    .B(_5022_),
    .C(_5020_),
    .Y(_5032_)
);

NAND3X1 _15508_ (
    .A(_5018_),
    .B(_5032_),
    .C(_5031_),
    .Y(_5033_)
);

AOI21X1 _15509_ (
    .A(_5033_),
    .B(_5030_),
    .C(_5017_),
    .Y(_5034_)
);

XNOR2X1 _15510_ (
    .A(_5016_),
    .B(_5010_),
    .Y(_5035_)
);

NAND3X1 _15511_ (
    .A(_5032_),
    .B(_5031_),
    .C(_5019_),
    .Y(_5037_)
);

OAI21X1 _15512_ (
    .A(_5029_),
    .B(_5024_),
    .C(_5018_),
    .Y(_5038_)
);

AOI21X1 _15513_ (
    .A(_5037_),
    .B(_5038_),
    .C(_5035_),
    .Y(_5039_)
);

NOR2X1 _15514_ (
    .A(_5034_),
    .B(_5039_),
    .Y(_5040_)
);

OAI21X1 _15515_ (
    .A(_4737_),
    .B(_4735_),
    .C(_4726_),
    .Y(_5041_)
);

NAND2X1 _15516_ (
    .A(areg_9_bF$buf3),
    .B(breg_16_bF$buf5),
    .Y(_5042_)
);

OAI21X1 _15517_ (
    .A(_4400_),
    .B(_5042_),
    .C(_4718_),
    .Y(_5043_)
);

NAND2X1 _15518_ (
    .A(areg_8_bF$buf3),
    .B(breg_17_bF$buf0),
    .Y(_5044_)
);

INVX1 _15519_ (
    .A(_5044_),
    .Y(_5045_)
);

AND2X2 _15520_ (
    .A(areg_9_bF$buf2),
    .B(breg_16_bF$buf4),
    .Y(_5046_)
);

AND2X2 _15521_ (
    .A(areg_10_bF$buf3),
    .B(breg_15_bF$buf0),
    .Y(_5048_)
);

NAND2X1 _15522_ (
    .A(_5046_),
    .B(_5048_),
    .Y(_5049_)
);

OAI21X1 _15523_ (
    .A(_7711__bF$buf0),
    .B(_2362__bF$buf5),
    .C(_5042_),
    .Y(_5050_)
);

NAND3X1 _15524_ (
    .A(_5045_),
    .B(_5050_),
    .C(_5049_),
    .Y(_5051_)
);

OAI21X1 _15525_ (
    .A(_6582__bF$buf2),
    .B(_2560__bF$buf4),
    .C(_5048_),
    .Y(_5052_)
);

OAI21X1 _15526_ (
    .A(_7711__bF$buf3),
    .B(_2362__bF$buf4),
    .C(_5046_),
    .Y(_5053_)
);

NAND3X1 _15527_ (
    .A(_5044_),
    .B(_5052_),
    .C(_5053_),
    .Y(_5054_)
);

NAND2X1 _15528_ (
    .A(areg_12_bF$buf4),
    .B(breg_13_bF$buf2),
    .Y(_5055_)
);

AND2X2 _15529_ (
    .A(_4723_),
    .B(_4771_),
    .Y(_5056_)
);

OAI22X1 _15530_ (
    .A(_4451_),
    .B(_5055_),
    .C(_5056_),
    .D(_4770_),
    .Y(_5057_)
);

NAND3X1 _15531_ (
    .A(_5051_),
    .B(_5054_),
    .C(_5057_),
    .Y(_5059_)
);

AOI21X1 _15532_ (
    .A(_5052_),
    .B(_5053_),
    .C(_5044_),
    .Y(_5060_)
);

AOI21X1 _15533_ (
    .A(_5050_),
    .B(_5049_),
    .C(_5045_),
    .Y(_5061_)
);

NOR2X1 _15534_ (
    .A(_4723_),
    .B(_4771_),
    .Y(_5062_)
);

OAI21X1 _15535_ (
    .A(_10869__bF$buf2),
    .B(_2586__bF$buf1),
    .C(_4723_),
    .Y(_5063_)
);

AOI21X1 _15536_ (
    .A(_4794_),
    .B(_5063_),
    .C(_5062_),
    .Y(_5064_)
);

OAI21X1 _15537_ (
    .A(_5060_),
    .B(_5061_),
    .C(_5064_),
    .Y(_5065_)
);

NAND3X1 _15538_ (
    .A(_5043_),
    .B(_5059_),
    .C(_5065_),
    .Y(_5066_)
);

AOI21X1 _15539_ (
    .A(_4395_),
    .B(_5046_),
    .C(_4727_),
    .Y(_5067_)
);

NOR3X1 _15540_ (
    .A(_5061_),
    .B(_5064_),
    .C(_5060_),
    .Y(_5068_)
);

AOI21X1 _15541_ (
    .A(_5051_),
    .B(_5054_),
    .C(_5057_),
    .Y(_5070_)
);

OAI21X1 _15542_ (
    .A(_5068_),
    .B(_5070_),
    .C(_5067_),
    .Y(_5071_)
);

NAND3X1 _15543_ (
    .A(_5041_),
    .B(_5066_),
    .C(_5071_),
    .Y(_5072_)
);

AOI21X1 _15544_ (
    .A(_4711_),
    .B(_4733_),
    .C(_4736_),
    .Y(_5073_)
);

NAND3X1 _15545_ (
    .A(_5064_),
    .B(_5051_),
    .C(_5054_),
    .Y(_5074_)
);

OAI21X1 _15546_ (
    .A(_5060_),
    .B(_5061_),
    .C(_5057_),
    .Y(_5075_)
);

AOI21X1 _15547_ (
    .A(_5074_),
    .B(_5075_),
    .C(_5067_),
    .Y(_5076_)
);

AOI21X1 _15548_ (
    .A(_5059_),
    .B(_5065_),
    .C(_5043_),
    .Y(_5077_)
);

OAI21X1 _15549_ (
    .A(_5076_),
    .B(_5077_),
    .C(_5073_),
    .Y(_5078_)
);

NAND3X1 _15550_ (
    .A(_5072_),
    .B(_5078_),
    .C(_5040_),
    .Y(_5079_)
);

NAND3X1 _15551_ (
    .A(_5037_),
    .B(_5035_),
    .C(_5038_),
    .Y(_5081_)
);

NOR3X1 _15552_ (
    .A(_5018_),
    .B(_5024_),
    .C(_5029_),
    .Y(_5082_)
);

AOI21X1 _15553_ (
    .A(_5032_),
    .B(_5031_),
    .C(_5019_),
    .Y(_5083_)
);

OAI21X1 _15554_ (
    .A(_5082_),
    .B(_5083_),
    .C(_5017_),
    .Y(_5084_)
);

NAND2X1 _15555_ (
    .A(_5081_),
    .B(_5084_),
    .Y(_5085_)
);

OAI21X1 _15556_ (
    .A(_5076_),
    .B(_5077_),
    .C(_5041_),
    .Y(_5086_)
);

NAND3X1 _15557_ (
    .A(_5073_),
    .B(_5066_),
    .C(_5071_),
    .Y(_5087_)
);

NAND3X1 _15558_ (
    .A(_5086_),
    .B(_5087_),
    .C(_5085_),
    .Y(_5088_)
);

OAI21X1 _15559_ (
    .A(_4801_),
    .B(_4808_),
    .C(_4810_),
    .Y(_5089_)
);

AOI21X1 _15560_ (
    .A(_5088_),
    .B(_5079_),
    .C(_5089_),
    .Y(_5090_)
);

AOI21X1 _15561_ (
    .A(_5086_),
    .B(_5087_),
    .C(_5085_),
    .Y(_5092_)
);

AOI21X1 _15562_ (
    .A(_5072_),
    .B(_5078_),
    .C(_5040_),
    .Y(_5093_)
);

AOI21X1 _15563_ (
    .A(_4769_),
    .B(_4809_),
    .C(_4805_),
    .Y(_5094_)
);

NOR3X1 _15564_ (
    .A(_5093_),
    .B(_5092_),
    .C(_5094_),
    .Y(_5095_)
);

OAI21X1 _15565_ (
    .A(_5095_),
    .B(_5090_),
    .C(_5009_),
    .Y(_5096_)
);

AND2X2 _15566_ (
    .A(_4747_),
    .B(_4739_),
    .Y(_5097_)
);

OAI21X1 _15567_ (
    .A(_5093_),
    .B(_5092_),
    .C(_5094_),
    .Y(_5098_)
);

NAND3X1 _15568_ (
    .A(_5089_),
    .B(_5088_),
    .C(_5079_),
    .Y(_5099_)
);

NAND3X1 _15569_ (
    .A(_5098_),
    .B(_5099_),
    .C(_5097_),
    .Y(_5100_)
);

NAND2X1 _15570_ (
    .A(_5100_),
    .B(_5096_),
    .Y(_5101_)
);

OAI21X1 _15571_ (
    .A(_4902_),
    .B(_4904_),
    .C(_4892_),
    .Y(_5103_)
);

NAND2X1 _15572_ (
    .A(_4788_),
    .B(_4793_),
    .Y(_5104_)
);

NAND2X1 _15573_ (
    .A(areg_11_bF$buf4),
    .B(breg_14_bF$buf1),
    .Y(_5105_)
);

NAND2X1 _15574_ (
    .A(breg_12_bF$buf0),
    .B(areg_13_bF$buf2),
    .Y(_5106_)
);

XOR2X1 _15575_ (
    .A(_5055_),
    .B(_5106_),
    .Y(_5107_)
);

XNOR2X1 _15576_ (
    .A(_5107_),
    .B(_5105_),
    .Y(_5108_)
);

OAI21X1 _15577_ (
    .A(_4786_),
    .B(_4776_),
    .C(_4780_),
    .Y(_5109_)
);

NAND2X1 _15578_ (
    .A(breg_11_bF$buf2),
    .B(areg_14_bF$buf1),
    .Y(_5110_)
);

INVX2 _15579_ (
    .A(_5110_),
    .Y(_5111_)
);

AND2X2 _15580_ (
    .A(breg_10_bF$buf2),
    .B(areg_15_bF$buf4),
    .Y(_5112_)
);

AND2X2 _15581_ (
    .A(breg_9_bF$buf5),
    .B(areg_16_bF$buf0),
    .Y(_5114_)
);

NAND2X1 _15582_ (
    .A(_5112_),
    .B(_5114_),
    .Y(_5115_)
);

OAI21X1 _15583_ (
    .A(_6044__bF$buf5),
    .B(_2669__bF$buf1),
    .C(_4783_),
    .Y(_5116_)
);

NAND3X1 _15584_ (
    .A(_5111_),
    .B(_5116_),
    .C(_5115_),
    .Y(_5117_)
);

AND2X2 _15585_ (
    .A(_5112_),
    .B(_5114_),
    .Y(_5118_)
);

NOR2X1 _15586_ (
    .A(_5112_),
    .B(_5114_),
    .Y(_5119_)
);

OAI21X1 _15587_ (
    .A(_5118_),
    .B(_5119_),
    .C(_5110_),
    .Y(_5120_)
);

NAND3X1 _15588_ (
    .A(_5117_),
    .B(_5109_),
    .C(_5120_),
    .Y(_5121_)
);

AOI21X1 _15589_ (
    .A(_4777_),
    .B(_4781_),
    .C(_4784_),
    .Y(_5122_)
);

OAI21X1 _15590_ (
    .A(_7217__bF$buf0),
    .B(_2465__bF$buf0),
    .C(_5114_),
    .Y(_5123_)
);

OAI21X1 _15591_ (
    .A(_6044__bF$buf4),
    .B(_2669__bF$buf0),
    .C(_5112_),
    .Y(_5125_)
);

AOI21X1 _15592_ (
    .A(_5123_),
    .B(_5125_),
    .C(_5110_),
    .Y(_5126_)
);

AOI21X1 _15593_ (
    .A(_5116_),
    .B(_5115_),
    .C(_5111_),
    .Y(_5127_)
);

OAI21X1 _15594_ (
    .A(_5126_),
    .B(_5127_),
    .C(_5122_),
    .Y(_5128_)
);

NAND3X1 _15595_ (
    .A(_5121_),
    .B(_5128_),
    .C(_5108_),
    .Y(_5129_)
);

INVX2 _15596_ (
    .A(_5105_),
    .Y(_5130_)
);

XNOR2X1 _15597_ (
    .A(_5107_),
    .B(_5130_),
    .Y(_5131_)
);

OAI21X1 _15598_ (
    .A(_5126_),
    .B(_5127_),
    .C(_5109_),
    .Y(_5132_)
);

NAND3X1 _15599_ (
    .A(_5122_),
    .B(_5117_),
    .C(_5120_),
    .Y(_5133_)
);

NAND3X1 _15600_ (
    .A(_5132_),
    .B(_5133_),
    .C(_5131_),
    .Y(_5134_)
);

OAI21X1 _15601_ (
    .A(_4817_),
    .B(_4843_),
    .C(_4834_),
    .Y(_5136_)
);

AOI21X1 _15602_ (
    .A(_5129_),
    .B(_5134_),
    .C(_5136_),
    .Y(_5137_)
);

AOI21X1 _15603_ (
    .A(_5132_),
    .B(_5133_),
    .C(_5131_),
    .Y(_5138_)
);

AOI21X1 _15604_ (
    .A(_5128_),
    .B(_5121_),
    .C(_5108_),
    .Y(_5139_)
);

AOI21X1 _15605_ (
    .A(_4816_),
    .B(_4839_),
    .C(_4842_),
    .Y(_5140_)
);

NOR3X1 _15606_ (
    .A(_5138_),
    .B(_5139_),
    .C(_5140_),
    .Y(_5141_)
);

OAI21X1 _15607_ (
    .A(_5141_),
    .B(_5137_),
    .C(_5104_),
    .Y(_5142_)
);

AND2X2 _15608_ (
    .A(_4793_),
    .B(_4788_),
    .Y(_5143_)
);

OAI21X1 _15609_ (
    .A(_5138_),
    .B(_5139_),
    .C(_5140_),
    .Y(_5144_)
);

NAND3X1 _15610_ (
    .A(_5129_),
    .B(_5134_),
    .C(_5136_),
    .Y(_5145_)
);

NAND3X1 _15611_ (
    .A(_5143_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5147_)
);

NAND2X1 _15612_ (
    .A(_5147_),
    .B(_5142_),
    .Y(_5148_)
);

AOI21X1 _15613_ (
    .A(_4871_),
    .B(_4877_),
    .C(_4847_),
    .Y(_5149_)
);

OAI21X1 _15614_ (
    .A(_4888_),
    .B(_5149_),
    .C(_4878_),
    .Y(_5150_)
);

NAND2X1 _15615_ (
    .A(breg_7_bF$buf0),
    .B(areg_18_bF$buf0),
    .Y(_5151_)
);

OAI21X1 _15616_ (
    .A(_4815_),
    .B(_5151_),
    .C(_4824_),
    .Y(_5152_)
);

NAND2X1 _15617_ (
    .A(breg[8]),
    .B(areg_17_bF$buf5),
    .Y(_5153_)
);

INVX1 _15618_ (
    .A(_5153_),
    .Y(_5154_)
);

AND2X2 _15619_ (
    .A(breg_7_bF$buf5),
    .B(areg_18_bF$buf5),
    .Y(_5155_)
);

AND2X2 _15620_ (
    .A(breg_6_bF$buf2),
    .B(areg_19_bF$buf1),
    .Y(_5156_)
);

NAND2X1 _15621_ (
    .A(_5155_),
    .B(_5156_),
    .Y(_5158_)
);

OAI21X1 _15622_ (
    .A(_5453__bF$buf1),
    .B(_3402__bF$buf1),
    .C(_5151_),
    .Y(_5159_)
);

NAND3X1 _15623_ (
    .A(_5154_),
    .B(_5159_),
    .C(_5158_),
    .Y(_5160_)
);

OAI21X1 _15624_ (
    .A(_4116__bF$buf2),
    .B(_3146__bF$buf1),
    .C(_5156_),
    .Y(_5161_)
);

OAI21X1 _15625_ (
    .A(_5453__bF$buf0),
    .B(_3402__bF$buf0),
    .C(_5155_),
    .Y(_5162_)
);

NAND3X1 _15626_ (
    .A(_5153_),
    .B(_5161_),
    .C(_5162_),
    .Y(_5163_)
);

NAND2X1 _15627_ (
    .A(_4831_),
    .B(_4849_),
    .Y(_5164_)
);

OAI21X1 _15628_ (
    .A(_4848_),
    .B(_4850_),
    .C(_5164_),
    .Y(_5165_)
);

NAND3X1 _15629_ (
    .A(_5165_),
    .B(_5160_),
    .C(_5163_),
    .Y(_5166_)
);

AOI21X1 _15630_ (
    .A(_5161_),
    .B(_5162_),
    .C(_5153_),
    .Y(_5167_)
);

AOI21X1 _15631_ (
    .A(_5159_),
    .B(_5158_),
    .C(_5154_),
    .Y(_5169_)
);

INVX1 _15632_ (
    .A(_4850_),
    .Y(_5170_)
);

AOI22X1 _15633_ (
    .A(_4831_),
    .B(_4849_),
    .C(_5170_),
    .D(_4872_),
    .Y(_5171_)
);

OAI21X1 _15634_ (
    .A(_5167_),
    .B(_5169_),
    .C(_5171_),
    .Y(_5172_)
);

NAND3X1 _15635_ (
    .A(_5152_),
    .B(_5166_),
    .C(_5172_),
    .Y(_5173_)
);

AND2X2 _15636_ (
    .A(_4824_),
    .B(_4822_),
    .Y(_5174_)
);

NAND3X1 _15637_ (
    .A(_5171_),
    .B(_5160_),
    .C(_5163_),
    .Y(_5175_)
);

OAI21X1 _15638_ (
    .A(_5167_),
    .B(_5169_),
    .C(_5165_),
    .Y(_5176_)
);

NAND3X1 _15639_ (
    .A(_5174_),
    .B(_5175_),
    .C(_5176_),
    .Y(_5177_)
);

AND2X2 _15640_ (
    .A(_5173_),
    .B(_5177_),
    .Y(_5178_)
);

AOI21X1 _15641_ (
    .A(_4865_),
    .B(_4861_),
    .C(_4854_),
    .Y(_5180_)
);

OAI21X1 _15642_ (
    .A(_5180_),
    .B(_4874_),
    .C(_4866_),
    .Y(_5181_)
);

NOR2X1 _15643_ (
    .A(_4258__bF$buf0),
    .B(_3958__bF$buf2),
    .Y(_5182_)
);

NAND2X1 _15644_ (
    .A(breg_4_bF$buf1),
    .B(areg_21_bF$buf2),
    .Y(_5183_)
);

NAND2X1 _15645_ (
    .A(breg_3_bF$buf3),
    .B(areg_22_bF$buf4),
    .Y(_5184_)
);

OR2X2 _15646_ (
    .A(_5183_),
    .B(_5184_),
    .Y(_5185_)
);

OAI21X1 _15647_ (
    .A(_2365_),
    .B(_4551__bF$buf3),
    .C(_5183_),
    .Y(_5186_)
);

NAND3X1 _15648_ (
    .A(_5182_),
    .B(_5186_),
    .C(_5185_),
    .Y(_5187_)
);

INVX1 _15649_ (
    .A(_5182_),
    .Y(_5188_)
);

NOR2X1 _15650_ (
    .A(_5183_),
    .B(_5184_),
    .Y(_5189_)
);

AND2X2 _15651_ (
    .A(_5183_),
    .B(_5184_),
    .Y(_5191_)
);

OAI21X1 _15652_ (
    .A(_5191_),
    .B(_5189_),
    .C(_5188_),
    .Y(_5192_)
);

AND2X2 _15653_ (
    .A(_5192_),
    .B(_5187_),
    .Y(_5193_)
);

OAI21X1 _15654_ (
    .A(_4855_),
    .B(_4859_),
    .C(_4858_),
    .Y(_5194_)
);

NAND2X1 _15655_ (
    .A(breg_2_bF$buf3),
    .B(areg_23_bF$buf0),
    .Y(_5195_)
);

INVX2 _15656_ (
    .A(_5195_),
    .Y(_5196_)
);

AND2X2 _15657_ (
    .A(breg_0_bF$buf4),
    .B(areg_25_bF$buf4),
    .Y(_5197_)
);

NAND2X1 _15658_ (
    .A(_4857_),
    .B(_5197_),
    .Y(_5198_)
);

AOI22X1 _15659_ (
    .A(breg_0_bF$buf3),
    .B(areg_25_bF$buf3),
    .C(breg_1_bF$buf3),
    .D(areg_24_bF$buf1),
    .Y(_5199_)
);

INVX2 _15660_ (
    .A(_5199_),
    .Y(_5200_)
);

NAND3X1 _15661_ (
    .A(_5196_),
    .B(_5200_),
    .C(_5198_),
    .Y(_5202_)
);

NAND2X1 _15662_ (
    .A(breg_0_bF$buf2),
    .B(areg_25_bF$buf2),
    .Y(_5203_)
);

NOR2X1 _15663_ (
    .A(_4863_),
    .B(_5203_),
    .Y(_5204_)
);

OAI21X1 _15664_ (
    .A(_5204_),
    .B(_5199_),
    .C(_5195_),
    .Y(_5205_)
);

NAND3X1 _15665_ (
    .A(_5194_),
    .B(_5205_),
    .C(_5202_),
    .Y(_5206_)
);

AOI21X1 _15666_ (
    .A(_4856_),
    .B(_4860_),
    .C(_4864_),
    .Y(_5207_)
);

NOR3X1 _15667_ (
    .A(_5195_),
    .B(_5199_),
    .C(_5204_),
    .Y(_5208_)
);

AOI21X1 _15668_ (
    .A(_5200_),
    .B(_5198_),
    .C(_5196_),
    .Y(_5209_)
);

OAI21X1 _15669_ (
    .A(_5209_),
    .B(_5208_),
    .C(_5207_),
    .Y(_5210_)
);

NAND3X1 _15670_ (
    .A(_5206_),
    .B(_5210_),
    .C(_5193_),
    .Y(_5211_)
);

NAND2X1 _15671_ (
    .A(_5187_),
    .B(_5192_),
    .Y(_5213_)
);

OAI21X1 _15672_ (
    .A(_5209_),
    .B(_5208_),
    .C(_5194_),
    .Y(_5214_)
);

NAND3X1 _15673_ (
    .A(_5205_),
    .B(_5207_),
    .C(_5202_),
    .Y(_5215_)
);

NAND3X1 _15674_ (
    .A(_5213_),
    .B(_5215_),
    .C(_5214_),
    .Y(_5216_)
);

NAND3X1 _15675_ (
    .A(_5216_),
    .B(_5181_),
    .C(_5211_),
    .Y(_5217_)
);

NOR3X1 _15676_ (
    .A(_4868_),
    .B(_4867_),
    .C(_4869_),
    .Y(_5218_)
);

AOI21X1 _15677_ (
    .A(_4853_),
    .B(_4870_),
    .C(_5218_),
    .Y(_5219_)
);

AOI21X1 _15678_ (
    .A(_5215_),
    .B(_5214_),
    .C(_5213_),
    .Y(_5220_)
);

AOI21X1 _15679_ (
    .A(_5206_),
    .B(_5210_),
    .C(_5193_),
    .Y(_5221_)
);

OAI21X1 _15680_ (
    .A(_5220_),
    .B(_5221_),
    .C(_5219_),
    .Y(_5222_)
);

NAND3X1 _15681_ (
    .A(_5217_),
    .B(_5178_),
    .C(_5222_),
    .Y(_5223_)
);

NAND2X1 _15682_ (
    .A(_5177_),
    .B(_5173_),
    .Y(_5224_)
);

OAI21X1 _15683_ (
    .A(_5220_),
    .B(_5221_),
    .C(_5181_),
    .Y(_5225_)
);

NAND3X1 _15684_ (
    .A(_5211_),
    .B(_5216_),
    .C(_5219_),
    .Y(_5226_)
);

NAND3X1 _15685_ (
    .A(_5224_),
    .B(_5226_),
    .C(_5225_),
    .Y(_5227_)
);

NAND3X1 _15686_ (
    .A(_5223_),
    .B(_5227_),
    .C(_5150_),
    .Y(_5228_)
);

NOR3X1 _15687_ (
    .A(_4882_),
    .B(_4881_),
    .C(_4880_),
    .Y(_5229_)
);

AOI21X1 _15688_ (
    .A(_4845_),
    .B(_4883_),
    .C(_5229_),
    .Y(_5230_)
);

AOI21X1 _15689_ (
    .A(_5226_),
    .B(_5225_),
    .C(_5224_),
    .Y(_5231_)
);

AOI21X1 _15690_ (
    .A(_5217_),
    .B(_5222_),
    .C(_5178_),
    .Y(_5232_)
);

OAI21X1 _15691_ (
    .A(_5231_),
    .B(_5232_),
    .C(_5230_),
    .Y(_5234_)
);

NAND3X1 _15692_ (
    .A(_5228_),
    .B(_5234_),
    .C(_5148_),
    .Y(_5235_)
);

NAND3X1 _15693_ (
    .A(_5104_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5236_)
);

OAI21X1 _15694_ (
    .A(_5141_),
    .B(_5137_),
    .C(_5143_),
    .Y(_5237_)
);

NAND2X1 _15695_ (
    .A(_5236_),
    .B(_5237_),
    .Y(_5238_)
);

OAI21X1 _15696_ (
    .A(_5231_),
    .B(_5232_),
    .C(_5150_),
    .Y(_5239_)
);

NAND3X1 _15697_ (
    .A(_5223_),
    .B(_5227_),
    .C(_5230_),
    .Y(_5240_)
);

NAND3X1 _15698_ (
    .A(_5240_),
    .B(_5239_),
    .C(_5238_),
    .Y(_5241_)
);

NAND3X1 _15699_ (
    .A(_5235_),
    .B(_5241_),
    .C(_5103_),
    .Y(_5242_)
);

AOI21X1 _15700_ (
    .A(_4898_),
    .B(_4812_),
    .C(_4903_),
    .Y(_5243_)
);

AOI21X1 _15701_ (
    .A(_5240_),
    .B(_5239_),
    .C(_5238_),
    .Y(_5246_)
);

AOI21X1 _15702_ (
    .A(_5228_),
    .B(_5234_),
    .C(_5148_),
    .Y(_5247_)
);

OAI21X1 _15703_ (
    .A(_5246_),
    .B(_5247_),
    .C(_5243_),
    .Y(_5248_)
);

NAND3X1 _15704_ (
    .A(_5242_),
    .B(_5248_),
    .C(_5101_),
    .Y(_5249_)
);

NAND3X1 _15705_ (
    .A(_5009_),
    .B(_5099_),
    .C(_5098_),
    .Y(_5250_)
);

OAI21X1 _15706_ (
    .A(_5095_),
    .B(_5090_),
    .C(_5097_),
    .Y(_5251_)
);

NAND2X1 _15707_ (
    .A(_5250_),
    .B(_5251_),
    .Y(_5252_)
);

NOR3X1 _15708_ (
    .A(_5246_),
    .B(_5247_),
    .C(_5243_),
    .Y(_5253_)
);

AOI21X1 _15709_ (
    .A(_5235_),
    .B(_5241_),
    .C(_5103_),
    .Y(_5254_)
);

OAI21X1 _15710_ (
    .A(_5253_),
    .B(_5254_),
    .C(_5252_),
    .Y(_5255_)
);

NAND3X1 _15711_ (
    .A(_5249_),
    .B(_5008_),
    .C(_5255_),
    .Y(_5257_)
);

AOI21X1 _15712_ (
    .A(_4914_),
    .B(_4766_),
    .C(_4920_),
    .Y(_5258_)
);

OAI21X1 _15713_ (
    .A(_5246_),
    .B(_5247_),
    .C(_5103_),
    .Y(_5259_)
);

NAND3X1 _15714_ (
    .A(_5235_),
    .B(_5241_),
    .C(_5243_),
    .Y(_5260_)
);

AOI21X1 _15715_ (
    .A(_5259_),
    .B(_5260_),
    .C(_5252_),
    .Y(_5261_)
);

AOI21X1 _15716_ (
    .A(_5242_),
    .B(_5248_),
    .C(_5101_),
    .Y(_5262_)
);

OAI21X1 _15717_ (
    .A(_5261_),
    .B(_5262_),
    .C(_5258_),
    .Y(_5263_)
);

NAND3X1 _15718_ (
    .A(_5263_),
    .B(_5007_),
    .C(_5257_),
    .Y(_5264_)
);

AND2X2 _15719_ (
    .A(_5006_),
    .B(_5002_),
    .Y(_5265_)
);

NOR3X1 _15720_ (
    .A(_5261_),
    .B(_5262_),
    .C(_5258_),
    .Y(_5266_)
);

AOI21X1 _15721_ (
    .A(_5249_),
    .B(_5255_),
    .C(_5008_),
    .Y(_5268_)
);

OAI21X1 _15722_ (
    .A(_5266_),
    .B(_5268_),
    .C(_5265_),
    .Y(_5269_)
);

NAND3X1 _15723_ (
    .A(_5264_),
    .B(_4969_),
    .C(_5269_),
    .Y(_5270_)
);

NOR3X1 _15724_ (
    .A(_4929_),
    .B(_4930_),
    .C(_4925_),
    .Y(_5271_)
);

AOI21X1 _15725_ (
    .A(_4673_),
    .B(_4931_),
    .C(_5271_),
    .Y(_5272_)
);

OAI21X1 _15726_ (
    .A(_5261_),
    .B(_5262_),
    .C(_5008_),
    .Y(_5273_)
);

NAND3X1 _15727_ (
    .A(_5258_),
    .B(_5249_),
    .C(_5255_),
    .Y(_5274_)
);

AOI21X1 _15728_ (
    .A(_5273_),
    .B(_5274_),
    .C(_5265_),
    .Y(_5275_)
);

AOI21X1 _15729_ (
    .A(_5263_),
    .B(_5257_),
    .C(_5007_),
    .Y(_5276_)
);

OAI21X1 _15730_ (
    .A(_5275_),
    .B(_5276_),
    .C(_5272_),
    .Y(_5277_)
);

NAND3X1 _15731_ (
    .A(_4967_),
    .B(_5277_),
    .C(_5270_),
    .Y(_5279_)
);

INVX2 _15732_ (
    .A(_4967_),
    .Y(_5280_)
);

NOR3X1 _15733_ (
    .A(_5275_),
    .B(_5276_),
    .C(_5272_),
    .Y(_5281_)
);

AOI21X1 _15734_ (
    .A(_5264_),
    .B(_5269_),
    .C(_4969_),
    .Y(_5282_)
);

OAI21X1 _15735_ (
    .A(_5281_),
    .B(_5282_),
    .C(_5280_),
    .Y(_5283_)
);

NAND3X1 _15736_ (
    .A(_4965_),
    .B(_5279_),
    .C(_5283_),
    .Y(_5284_)
);

AOI21X1 _15737_ (
    .A(_4943_),
    .B(_4654_),
    .C(_4945_),
    .Y(_5285_)
);

OAI21X1 _15738_ (
    .A(_5275_),
    .B(_5276_),
    .C(_4969_),
    .Y(_5286_)
);

NAND3X1 _15739_ (
    .A(_5264_),
    .B(_5272_),
    .C(_5269_),
    .Y(_5287_)
);

AOI21X1 _15740_ (
    .A(_5286_),
    .B(_5287_),
    .C(_5280_),
    .Y(_5288_)
);

AOI21X1 _15741_ (
    .A(_5277_),
    .B(_5270_),
    .C(_4967_),
    .Y(_5290_)
);

OAI21X1 _15742_ (
    .A(_5288_),
    .B(_5290_),
    .C(_5285_),
    .Y(_5291_)
);

NAND3X1 _15743_ (
    .A(_5284_),
    .B(_5291_),
    .C(_4964_),
    .Y(_5292_)
);

OAI21X1 _15744_ (
    .A(_5288_),
    .B(_5290_),
    .C(_4965_),
    .Y(_5293_)
);

NAND3X1 _15745_ (
    .A(_5279_),
    .B(_5285_),
    .C(_5283_),
    .Y(_5294_)
);

NAND3X1 _15746_ (
    .A(_5293_),
    .B(_4948_),
    .C(_5294_),
    .Y(_5295_)
);

NAND2X1 _15747_ (
    .A(_5295_),
    .B(_5292_),
    .Y(_5296_)
);

XNOR2X1 _15748_ (
    .A(_4963_),
    .B(_5296_),
    .Y(_0_[25])
);

NAND2X1 _15749_ (
    .A(_4957_),
    .B(_5292_),
    .Y(_5297_)
);

NAND2X1 _15750_ (
    .A(_5295_),
    .B(_5297_),
    .Y(_5298_)
);

INVX1 _15751_ (
    .A(_5298_),
    .Y(_5300_)
);

NOR2X1 _15752_ (
    .A(_4961_),
    .B(_5296_),
    .Y(_5301_)
);

AOI21X1 _15753_ (
    .A(_5301_),
    .B(_4648_),
    .C(_5300_),
    .Y(_5302_)
);

OAI21X1 _15754_ (
    .A(_5282_),
    .B(_5280_),
    .C(_5270_),
    .Y(_5303_)
);

INVX1 _15755_ (
    .A(_4999_),
    .Y(_5304_)
);

AOI21X1 _15756_ (
    .A(_4669_),
    .B(_5001_),
    .C(_5304_),
    .Y(_5305_)
);

INVX2 _15757_ (
    .A(_5305_),
    .Y(_5306_)
);

OAI21X1 _15758_ (
    .A(_5265_),
    .B(_5268_),
    .C(_5257_),
    .Y(_5307_)
);

AOI21X1 _15759_ (
    .A(_4662_),
    .B(_4989_),
    .C(_4985_),
    .Y(_5308_)
);

NAND2X1 _15760_ (
    .A(areg[0]),
    .B(breg_26_bF$buf4),
    .Y(_5309_)
);

INVX1 _15761_ (
    .A(_5309_),
    .Y(_5311_)
);

AND2X2 _15762_ (
    .A(areg_1_bF$buf0),
    .B(breg_25_bF$buf3),
    .Y(_5312_)
);

AND2X2 _15763_ (
    .A(areg_2_bF$buf0),
    .B(breg_24_bF$buf3),
    .Y(_5313_)
);

NAND2X1 _15764_ (
    .A(_5312_),
    .B(_5313_),
    .Y(_5314_)
);

INVX8 _15765_ (
    .A(breg_24_bF$buf2),
    .Y(_5315_)
);

OAI21X1 _15766_ (
    .A(_2519__bF$buf1),
    .B(_5315__bF$buf4),
    .C(_4973_),
    .Y(_5316_)
);

NAND3X1 _15767_ (
    .A(_5311_),
    .B(_5316_),
    .C(_5314_),
    .Y(_5317_)
);

INVX4 _15768_ (
    .A(breg_25_bF$buf2),
    .Y(_5318_)
);

OAI21X1 _15769_ (
    .A(_2661_),
    .B(_5318_),
    .C(_5313_),
    .Y(_5319_)
);

OAI21X1 _15770_ (
    .A(_2519__bF$buf0),
    .B(_5315__bF$buf3),
    .C(_5312_),
    .Y(_5320_)
);

NAND3X1 _15771_ (
    .A(_5309_),
    .B(_5319_),
    .C(_5320_),
    .Y(_5322_)
);

OR2X2 _15772_ (
    .A(_4679_),
    .B(_5012_),
    .Y(_5323_)
);

OAI21X1 _15773_ (
    .A(_5015_),
    .B(_5010_),
    .C(_5323_),
    .Y(_5324_)
);

NAND3X1 _15774_ (
    .A(_5317_),
    .B(_5322_),
    .C(_5324_),
    .Y(_5325_)
);

AOI21X1 _15775_ (
    .A(_5319_),
    .B(_5320_),
    .C(_5309_),
    .Y(_5326_)
);

AOI21X1 _15776_ (
    .A(_5316_),
    .B(_5314_),
    .C(_5311_),
    .Y(_5327_)
);

OAI21X1 _15777_ (
    .A(_2562__bF$buf3),
    .B(_3781__bF$buf1),
    .C(_4679_),
    .Y(_5328_)
);

AOI21X1 _15778_ (
    .A(_5011_),
    .B(_5328_),
    .C(_5013_),
    .Y(_5329_)
);

OAI21X1 _15779_ (
    .A(_5326_),
    .B(_5327_),
    .C(_5329_),
    .Y(_5330_)
);

NAND3X1 _15780_ (
    .A(_4974_),
    .B(_5325_),
    .C(_5330_),
    .Y(_5331_)
);

INVX1 _15781_ (
    .A(_4974_),
    .Y(_5333_)
);

NAND3X1 _15782_ (
    .A(_5329_),
    .B(_5317_),
    .C(_5322_),
    .Y(_5334_)
);

OAI21X1 _15783_ (
    .A(_5326_),
    .B(_5327_),
    .C(_5324_),
    .Y(_5335_)
);

NAND3X1 _15784_ (
    .A(_5333_),
    .B(_5334_),
    .C(_5335_),
    .Y(_5336_)
);

AOI21X1 _15785_ (
    .A(_5035_),
    .B(_5038_),
    .C(_5082_),
    .Y(_5337_)
);

NAND3X1 _15786_ (
    .A(_5331_),
    .B(_5336_),
    .C(_5337_),
    .Y(_5338_)
);

AOI21X1 _15787_ (
    .A(_5334_),
    .B(_5335_),
    .C(_5333_),
    .Y(_5339_)
);

AOI21X1 _15788_ (
    .A(_5325_),
    .B(_5330_),
    .C(_4974_),
    .Y(_5340_)
);

OAI21X1 _15789_ (
    .A(_5083_),
    .B(_5017_),
    .C(_5037_),
    .Y(_5341_)
);

OAI21X1 _15790_ (
    .A(_5339_),
    .B(_5340_),
    .C(_5341_),
    .Y(_5342_)
);

AOI21X1 _15791_ (
    .A(_5342_),
    .B(_5338_),
    .C(_4979_),
    .Y(_5344_)
);

NAND3X1 _15792_ (
    .A(_5331_),
    .B(_5336_),
    .C(_5341_),
    .Y(_5345_)
);

OAI21X1 _15793_ (
    .A(_5339_),
    .B(_5340_),
    .C(_5337_),
    .Y(_5346_)
);

AOI21X1 _15794_ (
    .A(_5346_),
    .B(_5345_),
    .C(_4980_),
    .Y(_5347_)
);

OAI21X1 _15795_ (
    .A(_5344_),
    .B(_5347_),
    .C(_5308_),
    .Y(_5348_)
);

OAI21X1 _15796_ (
    .A(_4986_),
    .B(_4972_),
    .C(_4988_),
    .Y(_5349_)
);

NAND3X1 _15797_ (
    .A(_4980_),
    .B(_5346_),
    .C(_5345_),
    .Y(_5350_)
);

NAND3X1 _15798_ (
    .A(_4979_),
    .B(_5342_),
    .C(_5338_),
    .Y(_5351_)
);

NAND3X1 _15799_ (
    .A(_5350_),
    .B(_5349_),
    .C(_5351_),
    .Y(_5352_)
);

AND2X2 _15800_ (
    .A(_5348_),
    .B(_5352_),
    .Y(_5353_)
);

OAI21X1 _15801_ (
    .A(_5097_),
    .B(_5090_),
    .C(_5099_),
    .Y(_5355_)
);

NAND2X1 _15802_ (
    .A(_5355_),
    .B(_5353_),
    .Y(_5356_)
);

NAND2X1 _15803_ (
    .A(_5352_),
    .B(_5348_),
    .Y(_5357_)
);

AOI21X1 _15804_ (
    .A(_5009_),
    .B(_5098_),
    .C(_5095_),
    .Y(_5358_)
);

NAND2X1 _15805_ (
    .A(_5357_),
    .B(_5358_),
    .Y(_5359_)
);

NAND3X1 _15806_ (
    .A(_4996_),
    .B(_5359_),
    .C(_5356_),
    .Y(_5360_)
);

INVX1 _15807_ (
    .A(_4996_),
    .Y(_5361_)
);

NOR2X1 _15808_ (
    .A(_5357_),
    .B(_5358_),
    .Y(_5362_)
);

NOR2X1 _15809_ (
    .A(_5355_),
    .B(_5353_),
    .Y(_5363_)
);

OAI21X1 _15810_ (
    .A(_5363_),
    .B(_5362_),
    .C(_5361_),
    .Y(_5364_)
);

NAND2X1 _15811_ (
    .A(_5360_),
    .B(_5364_),
    .Y(_5366_)
);

OAI21X1 _15812_ (
    .A(_5252_),
    .B(_5254_),
    .C(_5242_),
    .Y(_5367_)
);

NAND2X1 _15813_ (
    .A(_5072_),
    .B(_5079_),
    .Y(_5368_)
);

INVX4 _15814_ (
    .A(breg_23_bF$buf3),
    .Y(_5369_)
);

NOR2X1 _15815_ (
    .A(_2792_),
    .B(_5369_),
    .Y(_5370_)
);

INVX2 _15816_ (
    .A(_5370_),
    .Y(_5371_)
);

NAND2X1 _15817_ (
    .A(areg_4_bF$buf2),
    .B(breg_22_bF$buf0),
    .Y(_5372_)
);

NAND2X1 _15818_ (
    .A(areg_5_bF$buf1),
    .B(breg_21_bF$buf0),
    .Y(_5373_)
);

NOR2X1 _15819_ (
    .A(_5372_),
    .B(_5373_),
    .Y(_5374_)
);

AND2X2 _15820_ (
    .A(_5372_),
    .B(_5373_),
    .Y(_5375_)
);

NOR2X1 _15821_ (
    .A(_5374_),
    .B(_5375_),
    .Y(_5377_)
);

XNOR2X1 _15822_ (
    .A(_5377_),
    .B(_5371_),
    .Y(_5378_)
);

OAI21X1 _15823_ (
    .A(_5020_),
    .B(_5023_),
    .C(_5027_),
    .Y(_5379_)
);

NAND2X1 _15824_ (
    .A(areg_6_bF$buf1),
    .B(breg_20_bF$buf4),
    .Y(_5380_)
);

INVX2 _15825_ (
    .A(_5380_),
    .Y(_5381_)
);

AND2X2 _15826_ (
    .A(areg_7_bF$buf3),
    .B(breg_19_bF$buf4),
    .Y(_5382_)
);

AND2X2 _15827_ (
    .A(areg_8_bF$buf2),
    .B(breg_18_bF$buf3),
    .Y(_5383_)
);

NAND2X1 _15828_ (
    .A(_5382_),
    .B(_5383_),
    .Y(_5384_)
);

NAND2X1 _15829_ (
    .A(areg_7_bF$buf2),
    .B(breg_19_bF$buf3),
    .Y(_5385_)
);

OAI21X1 _15830_ (
    .A(_5190__bF$buf1),
    .B(_3529__bF$buf4),
    .C(_5385_),
    .Y(_5386_)
);

NAND3X1 _15831_ (
    .A(_5381_),
    .B(_5386_),
    .C(_5384_),
    .Y(_5388_)
);

NAND2X1 _15832_ (
    .A(areg_8_bF$buf1),
    .B(breg_18_bF$buf2),
    .Y(_5389_)
);

NOR2X1 _15833_ (
    .A(_5385_),
    .B(_5389_),
    .Y(_5390_)
);

NOR2X1 _15834_ (
    .A(_5382_),
    .B(_5383_),
    .Y(_5391_)
);

OAI21X1 _15835_ (
    .A(_5391_),
    .B(_5390_),
    .C(_5380_),
    .Y(_5392_)
);

NAND3X1 _15836_ (
    .A(_5388_),
    .B(_5392_),
    .C(_5379_),
    .Y(_5393_)
);

AOI21X1 _15837_ (
    .A(_5026_),
    .B(_5028_),
    .C(_5022_),
    .Y(_5394_)
);

NOR3X1 _15838_ (
    .A(_5380_),
    .B(_5390_),
    .C(_5391_),
    .Y(_5395_)
);

AOI21X1 _15839_ (
    .A(_5386_),
    .B(_5384_),
    .C(_5381_),
    .Y(_5396_)
);

OAI21X1 _15840_ (
    .A(_5395_),
    .B(_5396_),
    .C(_5394_),
    .Y(_5397_)
);

NAND3X1 _15841_ (
    .A(_5393_),
    .B(_5397_),
    .C(_5378_),
    .Y(_5399_)
);

XNOR2X1 _15842_ (
    .A(_5377_),
    .B(_5370_),
    .Y(_5400_)
);

NOR3X1 _15843_ (
    .A(_5394_),
    .B(_5396_),
    .C(_5395_),
    .Y(_5401_)
);

AOI21X1 _15844_ (
    .A(_5388_),
    .B(_5392_),
    .C(_5379_),
    .Y(_5402_)
);

OAI21X1 _15845_ (
    .A(_5401_),
    .B(_5402_),
    .C(_5400_),
    .Y(_5403_)
);

AND2X2 _15846_ (
    .A(_5403_),
    .B(_5399_),
    .Y(_5404_)
);

OAI21X1 _15847_ (
    .A(_5070_),
    .B(_5067_),
    .C(_5059_),
    .Y(_5405_)
);

INVX1 _15848_ (
    .A(_5048_),
    .Y(_5406_)
);

OAI21X1 _15849_ (
    .A(_5042_),
    .B(_5406_),
    .C(_5051_),
    .Y(_5407_)
);

NAND2X1 _15850_ (
    .A(areg_9_bF$buf1),
    .B(breg_17_bF$buf4),
    .Y(_5408_)
);

INVX1 _15851_ (
    .A(_5408_),
    .Y(_5410_)
);

AND2X2 _15852_ (
    .A(areg_10_bF$buf2),
    .B(breg_16_bF$buf3),
    .Y(_5411_)
);

AND2X2 _15853_ (
    .A(areg_11_bF$buf3),
    .B(breg_15_bF$buf5),
    .Y(_5412_)
);

NAND2X1 _15854_ (
    .A(_5411_),
    .B(_5412_),
    .Y(_5413_)
);

OAI22X1 _15855_ (
    .A(_7711__bF$buf2),
    .B(_2560__bF$buf3),
    .C(_9104__bF$buf0),
    .D(_2362__bF$buf3),
    .Y(_5414_)
);

NAND3X1 _15856_ (
    .A(_5410_),
    .B(_5414_),
    .C(_5413_),
    .Y(_5415_)
);

OAI21X1 _15857_ (
    .A(_7711__bF$buf1),
    .B(_2560__bF$buf2),
    .C(_5412_),
    .Y(_5416_)
);

OAI21X1 _15858_ (
    .A(_9104__bF$buf3),
    .B(_2362__bF$buf2),
    .C(_5411_),
    .Y(_5417_)
);

NAND3X1 _15859_ (
    .A(_5408_),
    .B(_5416_),
    .C(_5417_),
    .Y(_5418_)
);

NAND2X1 _15860_ (
    .A(areg_13_bF$buf1),
    .B(breg_13_bF$buf1),
    .Y(_5419_)
);

AND2X2 _15861_ (
    .A(_5055_),
    .B(_5106_),
    .Y(_5421_)
);

OAI22X1 _15862_ (
    .A(_4771_),
    .B(_5419_),
    .C(_5421_),
    .D(_5105_),
    .Y(_5422_)
);

NAND3X1 _15863_ (
    .A(_5415_),
    .B(_5418_),
    .C(_5422_),
    .Y(_5423_)
);

AOI21X1 _15864_ (
    .A(_5416_),
    .B(_5417_),
    .C(_5408_),
    .Y(_5424_)
);

AOI21X1 _15865_ (
    .A(_5414_),
    .B(_5413_),
    .C(_5410_),
    .Y(_5425_)
);

NOR2X1 _15866_ (
    .A(_5055_),
    .B(_5106_),
    .Y(_5426_)
);

OAI21X1 _15867_ (
    .A(_2586__bF$buf0),
    .B(_549__bF$buf3),
    .C(_5055_),
    .Y(_5427_)
);

AOI21X1 _15868_ (
    .A(_5130_),
    .B(_5427_),
    .C(_5426_),
    .Y(_5428_)
);

OAI21X1 _15869_ (
    .A(_5424_),
    .B(_5425_),
    .C(_5428_),
    .Y(_5429_)
);

NAND3X1 _15870_ (
    .A(_5407_),
    .B(_5423_),
    .C(_5429_),
    .Y(_5430_)
);

AOI21X1 _15871_ (
    .A(_4715_),
    .B(_5411_),
    .C(_5060_),
    .Y(_5432_)
);

NOR3X1 _15872_ (
    .A(_5425_),
    .B(_5428_),
    .C(_5424_),
    .Y(_5433_)
);

AOI21X1 _15873_ (
    .A(_5415_),
    .B(_5418_),
    .C(_5422_),
    .Y(_5434_)
);

OAI21X1 _15874_ (
    .A(_5433_),
    .B(_5434_),
    .C(_5432_),
    .Y(_5435_)
);

NAND3X1 _15875_ (
    .A(_5405_),
    .B(_5430_),
    .C(_5435_),
    .Y(_5436_)
);

AOI21X1 _15876_ (
    .A(_5043_),
    .B(_5065_),
    .C(_5068_),
    .Y(_5437_)
);

NAND3X1 _15877_ (
    .A(_5428_),
    .B(_5415_),
    .C(_5418_),
    .Y(_5438_)
);

OAI21X1 _15878_ (
    .A(_5424_),
    .B(_5425_),
    .C(_5422_),
    .Y(_5439_)
);

AOI21X1 _15879_ (
    .A(_5438_),
    .B(_5439_),
    .C(_5432_),
    .Y(_5440_)
);

AOI21X1 _15880_ (
    .A(_5423_),
    .B(_5429_),
    .C(_5407_),
    .Y(_5441_)
);

OAI21X1 _15881_ (
    .A(_5440_),
    .B(_5441_),
    .C(_5437_),
    .Y(_5443_)
);

NAND3X1 _15882_ (
    .A(_5436_),
    .B(_5443_),
    .C(_5404_),
    .Y(_5444_)
);

NAND2X1 _15883_ (
    .A(_5399_),
    .B(_5403_),
    .Y(_5445_)
);

OAI21X1 _15884_ (
    .A(_5440_),
    .B(_5441_),
    .C(_5405_),
    .Y(_5446_)
);

NAND3X1 _15885_ (
    .A(_5437_),
    .B(_5430_),
    .C(_5435_),
    .Y(_5447_)
);

NAND3X1 _15886_ (
    .A(_5446_),
    .B(_5445_),
    .C(_5447_),
    .Y(_5448_)
);

OAI21X1 _15887_ (
    .A(_5137_),
    .B(_5143_),
    .C(_5145_),
    .Y(_5449_)
);

AOI21X1 _15888_ (
    .A(_5448_),
    .B(_5444_),
    .C(_5449_),
    .Y(_5450_)
);

AOI21X1 _15889_ (
    .A(_5446_),
    .B(_5447_),
    .C(_5445_),
    .Y(_5451_)
);

AOI21X1 _15890_ (
    .A(_5436_),
    .B(_5443_),
    .C(_5404_),
    .Y(_5452_)
);

AOI21X1 _15891_ (
    .A(_5104_),
    .B(_5144_),
    .C(_5141_),
    .Y(_5454_)
);

NOR3X1 _15892_ (
    .A(_5452_),
    .B(_5451_),
    .C(_5454_),
    .Y(_5455_)
);

OAI21X1 _15893_ (
    .A(_5455_),
    .B(_5450_),
    .C(_5368_),
    .Y(_5456_)
);

AND2X2 _15894_ (
    .A(_5079_),
    .B(_5072_),
    .Y(_5457_)
);

OAI21X1 _15895_ (
    .A(_5452_),
    .B(_5451_),
    .C(_5454_),
    .Y(_5458_)
);

NAND3X1 _15896_ (
    .A(_5448_),
    .B(_5449_),
    .C(_5444_),
    .Y(_5459_)
);

NAND3X1 _15897_ (
    .A(_5459_),
    .B(_5458_),
    .C(_5457_),
    .Y(_5460_)
);

NAND2X1 _15898_ (
    .A(_5460_),
    .B(_5456_),
    .Y(_5461_)
);

AOI21X1 _15899_ (
    .A(_5223_),
    .B(_5227_),
    .C(_5150_),
    .Y(_5462_)
);

OAI21X1 _15900_ (
    .A(_5238_),
    .B(_5462_),
    .C(_5228_),
    .Y(_5463_)
);

NAND2X1 _15901_ (
    .A(_5121_),
    .B(_5129_),
    .Y(_5465_)
);

NAND2X1 _15902_ (
    .A(areg_12_bF$buf3),
    .B(breg_14_bF$buf0),
    .Y(_5466_)
);

INVX2 _15903_ (
    .A(_5466_),
    .Y(_5467_)
);

NAND2X1 _15904_ (
    .A(breg_13_bF$buf0),
    .B(areg_14_bF$buf0),
    .Y(_5468_)
);

OAI21X1 _15905_ (
    .A(_2586__bF$buf4),
    .B(_2287__bF$buf2),
    .C(_5419_),
    .Y(_5469_)
);

OAI21X1 _15906_ (
    .A(_5106_),
    .B(_5468_),
    .C(_5469_),
    .Y(_5470_)
);

XNOR2X1 _15907_ (
    .A(_5470_),
    .B(_5467_),
    .Y(_5471_)
);

OAI21X1 _15908_ (
    .A(_5119_),
    .B(_5110_),
    .C(_5115_),
    .Y(_5472_)
);

NAND2X1 _15909_ (
    .A(breg_11_bF$buf1),
    .B(areg_15_bF$buf3),
    .Y(_5473_)
);

INVX2 _15910_ (
    .A(_5473_),
    .Y(_5474_)
);

AND2X2 _15911_ (
    .A(breg_10_bF$buf1),
    .B(areg_17_bF$buf4),
    .Y(_5476_)
);

NAND2X1 _15912_ (
    .A(_5114_),
    .B(_5476_),
    .Y(_5477_)
);

NAND2X1 _15913_ (
    .A(breg_10_bF$buf0),
    .B(areg_16_bF$buf5),
    .Y(_5478_)
);

OAI21X1 _15914_ (
    .A(_6044__bF$buf3),
    .B(_2884__bF$buf1),
    .C(_5478_),
    .Y(_5479_)
);

NAND3X1 _15915_ (
    .A(_5474_),
    .B(_5479_),
    .C(_5477_),
    .Y(_5480_)
);

NAND2X1 _15916_ (
    .A(breg_9_bF$buf4),
    .B(areg_17_bF$buf3),
    .Y(_5481_)
);

NOR2X1 _15917_ (
    .A(_5478_),
    .B(_5481_),
    .Y(_5482_)
);

AND2X2 _15918_ (
    .A(_5478_),
    .B(_5481_),
    .Y(_5483_)
);

OAI21X1 _15919_ (
    .A(_5483_),
    .B(_5482_),
    .C(_5473_),
    .Y(_5484_)
);

NAND3X1 _15920_ (
    .A(_5480_),
    .B(_5484_),
    .C(_5472_),
    .Y(_5485_)
);

AOI21X1 _15921_ (
    .A(_5111_),
    .B(_5116_),
    .C(_5118_),
    .Y(_5487_)
);

NOR3X1 _15922_ (
    .A(_5473_),
    .B(_5482_),
    .C(_5483_),
    .Y(_5488_)
);

AOI21X1 _15923_ (
    .A(_5479_),
    .B(_5477_),
    .C(_5474_),
    .Y(_5489_)
);

OAI21X1 _15924_ (
    .A(_5488_),
    .B(_5489_),
    .C(_5487_),
    .Y(_5490_)
);

NAND3X1 _15925_ (
    .A(_5485_),
    .B(_5490_),
    .C(_5471_),
    .Y(_5491_)
);

XNOR2X1 _15926_ (
    .A(_5470_),
    .B(_5466_),
    .Y(_5492_)
);

OAI21X1 _15927_ (
    .A(_5488_),
    .B(_5489_),
    .C(_5472_),
    .Y(_5493_)
);

NAND3X1 _15928_ (
    .A(_5480_),
    .B(_5484_),
    .C(_5487_),
    .Y(_5494_)
);

NAND3X1 _15929_ (
    .A(_5494_),
    .B(_5493_),
    .C(_5492_),
    .Y(_5495_)
);

AOI21X1 _15930_ (
    .A(_5160_),
    .B(_5163_),
    .C(_5165_),
    .Y(_5496_)
);

OAI21X1 _15931_ (
    .A(_5496_),
    .B(_5174_),
    .C(_5166_),
    .Y(_5498_)
);

AOI21X1 _15932_ (
    .A(_5495_),
    .B(_5491_),
    .C(_5498_),
    .Y(_5499_)
);

AOI21X1 _15933_ (
    .A(_5494_),
    .B(_5493_),
    .C(_5492_),
    .Y(_5500_)
);

AOI21X1 _15934_ (
    .A(_5485_),
    .B(_5490_),
    .C(_5471_),
    .Y(_5501_)
);

NOR3X1 _15935_ (
    .A(_5169_),
    .B(_5171_),
    .C(_5167_),
    .Y(_5502_)
);

AOI21X1 _15936_ (
    .A(_5152_),
    .B(_5172_),
    .C(_5502_),
    .Y(_5503_)
);

NOR3X1 _15937_ (
    .A(_5500_),
    .B(_5501_),
    .C(_5503_),
    .Y(_5504_)
);

OAI21X1 _15938_ (
    .A(_5504_),
    .B(_5499_),
    .C(_5465_),
    .Y(_5505_)
);

AND2X2 _15939_ (
    .A(_5129_),
    .B(_5121_),
    .Y(_5506_)
);

OAI21X1 _15940_ (
    .A(_5500_),
    .B(_5501_),
    .C(_5503_),
    .Y(_5507_)
);

NAND3X1 _15941_ (
    .A(_5498_),
    .B(_5491_),
    .C(_5495_),
    .Y(_5509_)
);

NAND3X1 _15942_ (
    .A(_5509_),
    .B(_5507_),
    .C(_5506_),
    .Y(_5510_)
);

NAND2X1 _15943_ (
    .A(_5510_),
    .B(_5505_),
    .Y(_5511_)
);

AOI21X1 _15944_ (
    .A(_5216_),
    .B(_5211_),
    .C(_5181_),
    .Y(_5512_)
);

OAI21X1 _15945_ (
    .A(_5512_),
    .B(_5224_),
    .C(_5217_),
    .Y(_5513_)
);

INVX1 _15946_ (
    .A(_5156_),
    .Y(_5514_)
);

OAI21X1 _15947_ (
    .A(_5151_),
    .B(_5514_),
    .C(_5160_),
    .Y(_5515_)
);

NOR2X1 _15948_ (
    .A(_5420__bF$buf2),
    .B(_3146__bF$buf0),
    .Y(_5516_)
);

AND2X2 _15949_ (
    .A(breg_7_bF$buf4),
    .B(areg_19_bF$buf0),
    .Y(_5517_)
);

AND2X2 _15950_ (
    .A(breg_6_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_5518_)
);

NAND2X1 _15951_ (
    .A(_5517_),
    .B(_5518_),
    .Y(_5520_)
);

OAI22X1 _15952_ (
    .A(_5453__bF$buf5),
    .B(_3958__bF$buf1),
    .C(_4116__bF$buf1),
    .D(_3402__bF$buf3),
    .Y(_5521_)
);

NAND3X1 _15953_ (
    .A(_5516_),
    .B(_5521_),
    .C(_5520_),
    .Y(_5522_)
);

INVX1 _15954_ (
    .A(_5516_),
    .Y(_5523_)
);

OAI21X1 _15955_ (
    .A(_4116__bF$buf0),
    .B(_3402__bF$buf2),
    .C(_5518_),
    .Y(_5524_)
);

OAI21X1 _15956_ (
    .A(_5453__bF$buf4),
    .B(_3958__bF$buf0),
    .C(_5517_),
    .Y(_5525_)
);

NAND3X1 _15957_ (
    .A(_5524_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5526_)
);

AOI21X1 _15958_ (
    .A(_5182_),
    .B(_5186_),
    .C(_5189_),
    .Y(_5527_)
);

INVX1 _15959_ (
    .A(_5527_),
    .Y(_5528_)
);

AOI21X1 _15960_ (
    .A(_5522_),
    .B(_5526_),
    .C(_5528_),
    .Y(_5529_)
);

AOI21X1 _15961_ (
    .A(_5524_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5531_)
);

AOI21X1 _15962_ (
    .A(_5521_),
    .B(_5520_),
    .C(_5516_),
    .Y(_5532_)
);

NOR3X1 _15963_ (
    .A(_5532_),
    .B(_5527_),
    .C(_5531_),
    .Y(_5533_)
);

OAI21X1 _15964_ (
    .A(_5529_),
    .B(_5533_),
    .C(_5515_),
    .Y(_5534_)
);

INVX2 _15965_ (
    .A(_5515_),
    .Y(_5535_)
);

OAI21X1 _15966_ (
    .A(_5531_),
    .B(_5532_),
    .C(_5527_),
    .Y(_5536_)
);

NAND3X1 _15967_ (
    .A(_5522_),
    .B(_5526_),
    .C(_5528_),
    .Y(_5537_)
);

NAND3X1 _15968_ (
    .A(_5536_),
    .B(_5535_),
    .C(_5537_),
    .Y(_5538_)
);

NAND2X1 _15969_ (
    .A(_5538_),
    .B(_5534_),
    .Y(_5539_)
);

AOI21X1 _15970_ (
    .A(_5205_),
    .B(_5202_),
    .C(_5194_),
    .Y(_5540_)
);

OAI21X1 _15971_ (
    .A(_5540_),
    .B(_5213_),
    .C(_5206_),
    .Y(_5542_)
);

NAND2X1 _15972_ (
    .A(breg_5_bF$buf3),
    .B(areg_21_bF$buf1),
    .Y(_5543_)
);

INVX1 _15973_ (
    .A(_5543_),
    .Y(_5544_)
);

NAND2X1 _15974_ (
    .A(breg_4_bF$buf0),
    .B(areg_22_bF$buf3),
    .Y(_5545_)
);

NAND2X1 _15975_ (
    .A(breg_3_bF$buf2),
    .B(areg_23_bF$buf4),
    .Y(_5546_)
);

OR2X2 _15976_ (
    .A(_5545_),
    .B(_5546_),
    .Y(_5547_)
);

OAI21X1 _15977_ (
    .A(_2365_),
    .B(_4541__bF$buf2),
    .C(_5545_),
    .Y(_5548_)
);

NAND3X1 _15978_ (
    .A(_5544_),
    .B(_5548_),
    .C(_5547_),
    .Y(_5549_)
);

NOR2X1 _15979_ (
    .A(_5545_),
    .B(_5546_),
    .Y(_5550_)
);

AND2X2 _15980_ (
    .A(_5545_),
    .B(_5546_),
    .Y(_5551_)
);

OAI21X1 _15981_ (
    .A(_5551_),
    .B(_5550_),
    .C(_5543_),
    .Y(_5553_)
);

AND2X2 _15982_ (
    .A(_5549_),
    .B(_5553_),
    .Y(_5554_)
);

OAI21X1 _15983_ (
    .A(_5195_),
    .B(_5199_),
    .C(_5198_),
    .Y(_5555_)
);

NAND2X1 _15984_ (
    .A(breg_2_bF$buf2),
    .B(areg_24_bF$buf0),
    .Y(_5556_)
);

INVX2 _15985_ (
    .A(_5556_),
    .Y(_5557_)
);

AND2X2 _15986_ (
    .A(breg_1_bF$buf2),
    .B(areg_26_bF$buf4),
    .Y(_5558_)
);

NAND2X1 _15987_ (
    .A(_5197_),
    .B(_5558_),
    .Y(_5559_)
);

AOI22X1 _15988_ (
    .A(breg_0_bF$buf1),
    .B(areg_26_bF$buf3),
    .C(breg_1_bF$buf1),
    .D(areg_25_bF$buf1),
    .Y(_5560_)
);

INVX2 _15989_ (
    .A(_5560_),
    .Y(_5561_)
);

NAND3X1 _15990_ (
    .A(_5557_),
    .B(_5561_),
    .C(_5559_),
    .Y(_5562_)
);

NAND2X1 _15991_ (
    .A(breg_1_bF$buf0),
    .B(areg_26_bF$buf2),
    .Y(_5564_)
);

NOR2X1 _15992_ (
    .A(_5203_),
    .B(_5564_),
    .Y(_5565_)
);

OAI21X1 _15993_ (
    .A(_5565_),
    .B(_5560_),
    .C(_5556_),
    .Y(_5566_)
);

NAND3X1 _15994_ (
    .A(_5555_),
    .B(_5566_),
    .C(_5562_),
    .Y(_5567_)
);

AOI21X1 _15995_ (
    .A(_5196_),
    .B(_5200_),
    .C(_5204_),
    .Y(_5568_)
);

NOR3X1 _15996_ (
    .A(_5556_),
    .B(_5560_),
    .C(_5565_),
    .Y(_5569_)
);

AOI21X1 _15997_ (
    .A(_5561_),
    .B(_5559_),
    .C(_5557_),
    .Y(_5570_)
);

OAI21X1 _15998_ (
    .A(_5570_),
    .B(_5569_),
    .C(_5568_),
    .Y(_5571_)
);

NAND3X1 _15999_ (
    .A(_5567_),
    .B(_5571_),
    .C(_5554_),
    .Y(_5572_)
);

NAND2X1 _16000_ (
    .A(_5553_),
    .B(_5549_),
    .Y(_5573_)
);

OAI21X1 _16001_ (
    .A(_5570_),
    .B(_5569_),
    .C(_5555_),
    .Y(_5575_)
);

NAND3X1 _16002_ (
    .A(_5566_),
    .B(_5568_),
    .C(_5562_),
    .Y(_5576_)
);

NAND3X1 _16003_ (
    .A(_5573_),
    .B(_5576_),
    .C(_5575_),
    .Y(_5577_)
);

NAND3X1 _16004_ (
    .A(_5542_),
    .B(_5577_),
    .C(_5572_),
    .Y(_5578_)
);

NOR3X1 _16005_ (
    .A(_5208_),
    .B(_5207_),
    .C(_5209_),
    .Y(_5579_)
);

AOI21X1 _16006_ (
    .A(_5210_),
    .B(_5193_),
    .C(_5579_),
    .Y(_5580_)
);

AOI21X1 _16007_ (
    .A(_5576_),
    .B(_5575_),
    .C(_5573_),
    .Y(_5581_)
);

AOI21X1 _16008_ (
    .A(_5567_),
    .B(_5571_),
    .C(_5554_),
    .Y(_5582_)
);

OAI21X1 _16009_ (
    .A(_5581_),
    .B(_5582_),
    .C(_5580_),
    .Y(_5583_)
);

NAND3X1 _16010_ (
    .A(_5578_),
    .B(_5583_),
    .C(_5539_),
    .Y(_5584_)
);

NAND3X1 _16011_ (
    .A(_5515_),
    .B(_5536_),
    .C(_5537_),
    .Y(_5586_)
);

OAI21X1 _16012_ (
    .A(_5529_),
    .B(_5533_),
    .C(_5535_),
    .Y(_5587_)
);

NAND2X1 _16013_ (
    .A(_5586_),
    .B(_5587_),
    .Y(_5588_)
);

OAI21X1 _16014_ (
    .A(_5581_),
    .B(_5582_),
    .C(_5542_),
    .Y(_5589_)
);

NAND3X1 _16015_ (
    .A(_5572_),
    .B(_5577_),
    .C(_5580_),
    .Y(_5590_)
);

NAND3X1 _16016_ (
    .A(_5590_),
    .B(_5589_),
    .C(_5588_),
    .Y(_5591_)
);

NAND3X1 _16017_ (
    .A(_5513_),
    .B(_5584_),
    .C(_5591_),
    .Y(_5592_)
);

NOR3X1 _16018_ (
    .A(_5220_),
    .B(_5221_),
    .C(_5219_),
    .Y(_5593_)
);

AOI21X1 _16019_ (
    .A(_5178_),
    .B(_5222_),
    .C(_5593_),
    .Y(_5594_)
);

AOI21X1 _16020_ (
    .A(_5590_),
    .B(_5589_),
    .C(_5588_),
    .Y(_5595_)
);

AOI21X1 _16021_ (
    .A(_5578_),
    .B(_5583_),
    .C(_5539_),
    .Y(_5597_)
);

OAI21X1 _16022_ (
    .A(_5595_),
    .B(_5597_),
    .C(_5594_),
    .Y(_5598_)
);

NAND3X1 _16023_ (
    .A(_5592_),
    .B(_5511_),
    .C(_5598_),
    .Y(_5599_)
);

NAND3X1 _16024_ (
    .A(_5465_),
    .B(_5509_),
    .C(_5507_),
    .Y(_5600_)
);

OAI21X1 _16025_ (
    .A(_5504_),
    .B(_5499_),
    .C(_5506_),
    .Y(_5601_)
);

NAND2X1 _16026_ (
    .A(_5600_),
    .B(_5601_),
    .Y(_5602_)
);

OAI21X1 _16027_ (
    .A(_5595_),
    .B(_5597_),
    .C(_5513_),
    .Y(_5603_)
);

NAND3X1 _16028_ (
    .A(_5584_),
    .B(_5591_),
    .C(_5594_),
    .Y(_5604_)
);

NAND3X1 _16029_ (
    .A(_5604_),
    .B(_5602_),
    .C(_5603_),
    .Y(_5605_)
);

NAND3X1 _16030_ (
    .A(_5599_),
    .B(_5605_),
    .C(_5463_),
    .Y(_5606_)
);

NOR3X1 _16031_ (
    .A(_5231_),
    .B(_5232_),
    .C(_5230_),
    .Y(_5608_)
);

AOI21X1 _16032_ (
    .A(_5148_),
    .B(_5234_),
    .C(_5608_),
    .Y(_5609_)
);

AOI21X1 _16033_ (
    .A(_5604_),
    .B(_5603_),
    .C(_5602_),
    .Y(_5610_)
);

AOI21X1 _16034_ (
    .A(_5592_),
    .B(_5598_),
    .C(_5511_),
    .Y(_5611_)
);

OAI21X1 _16035_ (
    .A(_5610_),
    .B(_5611_),
    .C(_5609_),
    .Y(_5612_)
);

NAND3X1 _16036_ (
    .A(_5606_),
    .B(_5612_),
    .C(_5461_),
    .Y(_5613_)
);

NAND3X1 _16037_ (
    .A(_5368_),
    .B(_5459_),
    .C(_5458_),
    .Y(_5614_)
);

OAI21X1 _16038_ (
    .A(_5455_),
    .B(_5450_),
    .C(_5457_),
    .Y(_5615_)
);

NAND2X1 _16039_ (
    .A(_5614_),
    .B(_5615_),
    .Y(_5616_)
);

OAI21X1 _16040_ (
    .A(_5610_),
    .B(_5611_),
    .C(_5463_),
    .Y(_5617_)
);

NAND3X1 _16041_ (
    .A(_5599_),
    .B(_5605_),
    .C(_5609_),
    .Y(_5619_)
);

NAND3X1 _16042_ (
    .A(_5617_),
    .B(_5619_),
    .C(_5616_),
    .Y(_5620_)
);

NAND3X1 _16043_ (
    .A(_5613_),
    .B(_5620_),
    .C(_5367_),
    .Y(_5621_)
);

AOI21X1 _16044_ (
    .A(_5248_),
    .B(_5101_),
    .C(_5253_),
    .Y(_5622_)
);

AOI21X1 _16045_ (
    .A(_5619_),
    .B(_5617_),
    .C(_5616_),
    .Y(_5623_)
);

AOI21X1 _16046_ (
    .A(_5606_),
    .B(_5612_),
    .C(_5461_),
    .Y(_5624_)
);

OAI21X1 _16047_ (
    .A(_5623_),
    .B(_5624_),
    .C(_5622_),
    .Y(_5625_)
);

NAND3X1 _16048_ (
    .A(_5366_),
    .B(_5621_),
    .C(_5625_),
    .Y(_5626_)
);

NAND3X1 _16049_ (
    .A(_5361_),
    .B(_5359_),
    .C(_5356_),
    .Y(_5627_)
);

OAI21X1 _16050_ (
    .A(_5363_),
    .B(_5362_),
    .C(_4996_),
    .Y(_5628_)
);

NAND2X1 _16051_ (
    .A(_5627_),
    .B(_5628_),
    .Y(_5630_)
);

NOR3X1 _16052_ (
    .A(_5623_),
    .B(_5624_),
    .C(_5622_),
    .Y(_5631_)
);

AOI21X1 _16053_ (
    .A(_5613_),
    .B(_5620_),
    .C(_5367_),
    .Y(_5632_)
);

OAI21X1 _16054_ (
    .A(_5631_),
    .B(_5632_),
    .C(_5630_),
    .Y(_5633_)
);

NAND3X1 _16055_ (
    .A(_5626_),
    .B(_5633_),
    .C(_5307_),
    .Y(_5634_)
);

AOI21X1 _16056_ (
    .A(_5007_),
    .B(_5263_),
    .C(_5266_),
    .Y(_5635_)
);

OAI21X1 _16057_ (
    .A(_5623_),
    .B(_5624_),
    .C(_5367_),
    .Y(_5636_)
);

NAND3X1 _16058_ (
    .A(_5613_),
    .B(_5620_),
    .C(_5622_),
    .Y(_5637_)
);

AOI21X1 _16059_ (
    .A(_5637_),
    .B(_5636_),
    .C(_5630_),
    .Y(_5638_)
);

AOI21X1 _16060_ (
    .A(_5621_),
    .B(_5625_),
    .C(_5366_),
    .Y(_5639_)
);

OAI21X1 _16061_ (
    .A(_5638_),
    .B(_5639_),
    .C(_5635_),
    .Y(_5641_)
);

NAND3X1 _16062_ (
    .A(_5306_),
    .B(_5641_),
    .C(_5634_),
    .Y(_5642_)
);

NOR3X1 _16063_ (
    .A(_5638_),
    .B(_5639_),
    .C(_5635_),
    .Y(_5643_)
);

AOI21X1 _16064_ (
    .A(_5626_),
    .B(_5633_),
    .C(_5307_),
    .Y(_5644_)
);

OAI21X1 _16065_ (
    .A(_5643_),
    .B(_5644_),
    .C(_5305_),
    .Y(_5645_)
);

NAND3X1 _16066_ (
    .A(_5642_),
    .B(_5303_),
    .C(_5645_),
    .Y(_5646_)
);

AOI21X1 _16067_ (
    .A(_5277_),
    .B(_4967_),
    .C(_5281_),
    .Y(_5647_)
);

OAI21X1 _16068_ (
    .A(_5638_),
    .B(_5639_),
    .C(_5307_),
    .Y(_5648_)
);

NAND3X1 _16069_ (
    .A(_5635_),
    .B(_5626_),
    .C(_5633_),
    .Y(_5649_)
);

AOI21X1 _16070_ (
    .A(_5648_),
    .B(_5649_),
    .C(_5305_),
    .Y(_5650_)
);

AOI21X1 _16071_ (
    .A(_5641_),
    .B(_5634_),
    .C(_5306_),
    .Y(_5652_)
);

OAI21X1 _16072_ (
    .A(_5652_),
    .B(_5650_),
    .C(_5647_),
    .Y(_5653_)
);

NAND3X1 _16073_ (
    .A(_5653_),
    .B(_5646_),
    .C(_5284_),
    .Y(_5654_)
);

INVX1 _16074_ (
    .A(_5284_),
    .Y(_5655_)
);

NAND2X1 _16075_ (
    .A(_5653_),
    .B(_5646_),
    .Y(_5656_)
);

NAND2X1 _16076_ (
    .A(_5655_),
    .B(_5656_),
    .Y(_5657_)
);

NAND2X1 _16077_ (
    .A(_5654_),
    .B(_5657_),
    .Y(_5658_)
);

XNOR2X1 _16078_ (
    .A(_5302_),
    .B(_5658_),
    .Y(_0_[26])
);

NOR2X1 _16079_ (
    .A(_5284_),
    .B(_5656_),
    .Y(_5659_)
);

INVX1 _16080_ (
    .A(_5659_),
    .Y(_5660_)
);

INVX1 _16081_ (
    .A(_5658_),
    .Y(_5662_)
);

OAI21X1 _16082_ (
    .A(_5302_),
    .B(_5662_),
    .C(_5660_),
    .Y(_5663_)
);

NOR3X1 _16083_ (
    .A(_5652_),
    .B(_5650_),
    .C(_5647_),
    .Y(_5664_)
);

OAI21X1 _16084_ (
    .A(_5644_),
    .B(_5305_),
    .C(_5634_),
    .Y(_5665_)
);

OAI21X1 _16085_ (
    .A(_5363_),
    .B(_4996_),
    .C(_5356_),
    .Y(_5666_)
);

OAI21X1 _16086_ (
    .A(_5632_),
    .B(_5630_),
    .C(_5621_),
    .Y(_5667_)
);

INVX8 _16087_ (
    .A(breg_27_bF$buf5),
    .Y(_5668_)
);

NOR2X1 _16088_ (
    .A(_2376__bF$buf1),
    .B(_5668__bF$buf5),
    .Y(_5669_)
);

AOI21X1 _16089_ (
    .A(_5331_),
    .B(_5336_),
    .C(_5341_),
    .Y(_5670_)
);

OAI21X1 _16090_ (
    .A(_5670_),
    .B(_4979_),
    .C(_5345_),
    .Y(_5671_)
);

NAND2X1 _16091_ (
    .A(_5325_),
    .B(_5331_),
    .Y(_5673_)
);

NAND2X1 _16092_ (
    .A(areg_2_bF$buf4),
    .B(breg_24_bF$buf1),
    .Y(_5674_)
);

OAI21X1 _16093_ (
    .A(_4973_),
    .B(_5674_),
    .C(_5317_),
    .Y(_5675_)
);

INVX8 _16094_ (
    .A(breg_26_bF$buf3),
    .Y(_5676_)
);

NOR2X1 _16095_ (
    .A(_2661_),
    .B(_5676_),
    .Y(_5677_)
);

AND2X2 _16096_ (
    .A(areg_2_bF$buf3),
    .B(breg_25_bF$buf1),
    .Y(_5678_)
);

AND2X2 _16097_ (
    .A(areg_3_bF$buf3),
    .B(breg_24_bF$buf0),
    .Y(_5679_)
);

NAND2X1 _16098_ (
    .A(_5678_),
    .B(_5679_),
    .Y(_5680_)
);

NAND2X1 _16099_ (
    .A(areg_2_bF$buf2),
    .B(breg_25_bF$buf0),
    .Y(_5681_)
);

OAI21X1 _16100_ (
    .A(_2792_),
    .B(_5315__bF$buf2),
    .C(_5681_),
    .Y(_5682_)
);

NAND3X1 _16101_ (
    .A(_5677_),
    .B(_5682_),
    .C(_5680_),
    .Y(_5684_)
);

NAND2X1 _16102_ (
    .A(areg_3_bF$buf2),
    .B(breg_25_bF$buf5),
    .Y(_5685_)
);

OAI21X1 _16103_ (
    .A(_5674_),
    .B(_5685_),
    .C(_5682_),
    .Y(_5686_)
);

OAI21X1 _16104_ (
    .A(_2661_),
    .B(_5676_),
    .C(_5686_),
    .Y(_5687_)
);

NAND2X1 _16105_ (
    .A(areg_5_bF$buf0),
    .B(breg_22_bF$buf4),
    .Y(_5688_)
);

OAI22X1 _16106_ (
    .A(_5012_),
    .B(_5688_),
    .C(_5371_),
    .D(_5375_),
    .Y(_5689_)
);

NAND3X1 _16107_ (
    .A(_5684_),
    .B(_5689_),
    .C(_5687_),
    .Y(_5690_)
);

INVX1 _16108_ (
    .A(_5677_),
    .Y(_5691_)
);

OAI21X1 _16109_ (
    .A(_2519__bF$buf3),
    .B(_5318_),
    .C(_5679_),
    .Y(_5692_)
);

OAI21X1 _16110_ (
    .A(_2792_),
    .B(_5315__bF$buf1),
    .C(_5678_),
    .Y(_5693_)
);

AOI21X1 _16111_ (
    .A(_5692_),
    .B(_5693_),
    .C(_5691_),
    .Y(_5695_)
);

AOI21X1 _16112_ (
    .A(_5682_),
    .B(_5680_),
    .C(_5677_),
    .Y(_5696_)
);

OAI21X1 _16113_ (
    .A(_2825__bF$buf4),
    .B(_3781__bF$buf0),
    .C(_5372_),
    .Y(_5697_)
);

AOI21X1 _16114_ (
    .A(_5370_),
    .B(_5697_),
    .C(_5374_),
    .Y(_5698_)
);

OAI21X1 _16115_ (
    .A(_5695_),
    .B(_5696_),
    .C(_5698_),
    .Y(_5699_)
);

NAND3X1 _16116_ (
    .A(_5675_),
    .B(_5699_),
    .C(_5690_),
    .Y(_5700_)
);

INVX1 _16117_ (
    .A(_5675_),
    .Y(_5701_)
);

NAND3X1 _16118_ (
    .A(_5684_),
    .B(_5698_),
    .C(_5687_),
    .Y(_5702_)
);

OAI21X1 _16119_ (
    .A(_5695_),
    .B(_5696_),
    .C(_5689_),
    .Y(_5703_)
);

NAND3X1 _16120_ (
    .A(_5703_),
    .B(_5701_),
    .C(_5702_),
    .Y(_5704_)
);

OAI21X1 _16121_ (
    .A(_5400_),
    .B(_5402_),
    .C(_5393_),
    .Y(_5706_)
);

NAND3X1 _16122_ (
    .A(_5700_),
    .B(_5704_),
    .C(_5706_),
    .Y(_5707_)
);

AOI21X1 _16123_ (
    .A(_5703_),
    .B(_5702_),
    .C(_5701_),
    .Y(_5708_)
);

AOI21X1 _16124_ (
    .A(_5699_),
    .B(_5690_),
    .C(_5675_),
    .Y(_5709_)
);

AOI21X1 _16125_ (
    .A(_5397_),
    .B(_5378_),
    .C(_5401_),
    .Y(_5710_)
);

OAI21X1 _16126_ (
    .A(_5708_),
    .B(_5709_),
    .C(_5710_),
    .Y(_5711_)
);

NAND3X1 _16127_ (
    .A(_5673_),
    .B(_5707_),
    .C(_5711_),
    .Y(_5712_)
);

INVX2 _16128_ (
    .A(_5673_),
    .Y(_5713_)
);

NAND3X1 _16129_ (
    .A(_5700_),
    .B(_5704_),
    .C(_5710_),
    .Y(_5714_)
);

OAI21X1 _16130_ (
    .A(_5708_),
    .B(_5709_),
    .C(_5706_),
    .Y(_5715_)
);

NAND3X1 _16131_ (
    .A(_5714_),
    .B(_5713_),
    .C(_5715_),
    .Y(_5717_)
);

NAND3X1 _16132_ (
    .A(_5712_),
    .B(_5671_),
    .C(_5717_),
    .Y(_5718_)
);

NAND2X1 _16133_ (
    .A(_5331_),
    .B(_5336_),
    .Y(_5719_)
);

NOR2X1 _16134_ (
    .A(_5337_),
    .B(_5719_),
    .Y(_5720_)
);

AOI21X1 _16135_ (
    .A(_4980_),
    .B(_5346_),
    .C(_5720_),
    .Y(_5721_)
);

AOI21X1 _16136_ (
    .A(_5714_),
    .B(_5715_),
    .C(_5713_),
    .Y(_5722_)
);

AOI21X1 _16137_ (
    .A(_5707_),
    .B(_5711_),
    .C(_5673_),
    .Y(_5723_)
);

OAI21X1 _16138_ (
    .A(_5722_),
    .B(_5723_),
    .C(_5721_),
    .Y(_5724_)
);

NAND3X1 _16139_ (
    .A(_5669_),
    .B(_5718_),
    .C(_5724_),
    .Y(_5725_)
);

INVX2 _16140_ (
    .A(_5669_),
    .Y(_5726_)
);

OAI21X1 _16141_ (
    .A(_5722_),
    .B(_5723_),
    .C(_5671_),
    .Y(_5728_)
);

NAND3X1 _16142_ (
    .A(_5712_),
    .B(_5717_),
    .C(_5721_),
    .Y(_5729_)
);

NAND3X1 _16143_ (
    .A(_5726_),
    .B(_5728_),
    .C(_5729_),
    .Y(_5730_)
);

OAI21X1 _16144_ (
    .A(_5457_),
    .B(_5450_),
    .C(_5459_),
    .Y(_5731_)
);

NAND3X1 _16145_ (
    .A(_5731_),
    .B(_5725_),
    .C(_5730_),
    .Y(_5732_)
);

AOI21X1 _16146_ (
    .A(_5728_),
    .B(_5729_),
    .C(_5726_),
    .Y(_5733_)
);

AOI21X1 _16147_ (
    .A(_5718_),
    .B(_5724_),
    .C(_5669_),
    .Y(_5734_)
);

AOI21X1 _16148_ (
    .A(_5368_),
    .B(_5458_),
    .C(_5455_),
    .Y(_5735_)
);

OAI21X1 _16149_ (
    .A(_5733_),
    .B(_5734_),
    .C(_5735_),
    .Y(_5736_)
);

NAND3X1 _16150_ (
    .A(_5352_),
    .B(_5732_),
    .C(_5736_),
    .Y(_5737_)
);

INVX1 _16151_ (
    .A(_5352_),
    .Y(_5739_)
);

NAND3X1 _16152_ (
    .A(_5725_),
    .B(_5730_),
    .C(_5735_),
    .Y(_5740_)
);

OAI21X1 _16153_ (
    .A(_5733_),
    .B(_5734_),
    .C(_5731_),
    .Y(_5741_)
);

NAND3X1 _16154_ (
    .A(_5739_),
    .B(_5740_),
    .C(_5741_),
    .Y(_5742_)
);

NAND2X1 _16155_ (
    .A(_5737_),
    .B(_5742_),
    .Y(_5743_)
);

AOI21X1 _16156_ (
    .A(_5599_),
    .B(_5605_),
    .C(_5463_),
    .Y(_5744_)
);

OAI21X1 _16157_ (
    .A(_5616_),
    .B(_5744_),
    .C(_5606_),
    .Y(_5745_)
);

NAND2X1 _16158_ (
    .A(_5436_),
    .B(_5444_),
    .Y(_5746_)
);

NAND2X1 _16159_ (
    .A(areg_4_bF$buf1),
    .B(breg_23_bF$buf2),
    .Y(_5747_)
);

INVX2 _16160_ (
    .A(_5747_),
    .Y(_5748_)
);

NAND2X1 _16161_ (
    .A(areg_6_bF$buf0),
    .B(breg_21_bF$buf4),
    .Y(_5750_)
);

XOR2X1 _16162_ (
    .A(_5688_),
    .B(_5750_),
    .Y(_5751_)
);

XNOR2X1 _16163_ (
    .A(_5751_),
    .B(_5748_),
    .Y(_5752_)
);

OAI21X1 _16164_ (
    .A(_5391_),
    .B(_5380_),
    .C(_5384_),
    .Y(_5753_)
);

NAND2X1 _16165_ (
    .A(areg_7_bF$buf1),
    .B(breg_20_bF$buf3),
    .Y(_5754_)
);

AND2X2 _16166_ (
    .A(areg_9_bF$buf0),
    .B(breg_18_bF$buf1),
    .Y(_5755_)
);

OAI21X1 _16167_ (
    .A(_5190__bF$buf0),
    .B(_3253__bF$buf1),
    .C(_5755_),
    .Y(_5756_)
);

AND2X2 _16168_ (
    .A(areg_8_bF$buf0),
    .B(breg_19_bF$buf2),
    .Y(_5757_)
);

OAI21X1 _16169_ (
    .A(_6582__bF$buf1),
    .B(_3529__bF$buf3),
    .C(_5757_),
    .Y(_5758_)
);

AOI21X1 _16170_ (
    .A(_5756_),
    .B(_5758_),
    .C(_5754_),
    .Y(_5759_)
);

INVX2 _16171_ (
    .A(_5754_),
    .Y(_5761_)
);

NAND2X1 _16172_ (
    .A(_5757_),
    .B(_5755_),
    .Y(_5762_)
);

OAI22X1 _16173_ (
    .A(_5190__bF$buf3),
    .B(_3253__bF$buf0),
    .C(_6582__bF$buf0),
    .D(_3529__bF$buf2),
    .Y(_5763_)
);

AOI21X1 _16174_ (
    .A(_5763_),
    .B(_5762_),
    .C(_5761_),
    .Y(_5764_)
);

OAI21X1 _16175_ (
    .A(_5759_),
    .B(_5764_),
    .C(_5753_),
    .Y(_5765_)
);

AOI21X1 _16176_ (
    .A(_5381_),
    .B(_5386_),
    .C(_5390_),
    .Y(_5766_)
);

NAND3X1 _16177_ (
    .A(_5761_),
    .B(_5763_),
    .C(_5762_),
    .Y(_5767_)
);

NAND2X1 _16178_ (
    .A(areg_9_bF$buf4),
    .B(breg_19_bF$buf1),
    .Y(_5768_)
);

NOR2X1 _16179_ (
    .A(_5389_),
    .B(_5768_),
    .Y(_5769_)
);

NOR2X1 _16180_ (
    .A(_5757_),
    .B(_5755_),
    .Y(_5770_)
);

OAI21X1 _16181_ (
    .A(_5770_),
    .B(_5769_),
    .C(_5754_),
    .Y(_5772_)
);

NAND3X1 _16182_ (
    .A(_5766_),
    .B(_5767_),
    .C(_5772_),
    .Y(_5773_)
);

AOI21X1 _16183_ (
    .A(_5765_),
    .B(_5773_),
    .C(_5752_),
    .Y(_5774_)
);

XNOR2X1 _16184_ (
    .A(_5751_),
    .B(_5747_),
    .Y(_5775_)
);

NAND3X1 _16185_ (
    .A(_5767_),
    .B(_5753_),
    .C(_5772_),
    .Y(_5776_)
);

OAI21X1 _16186_ (
    .A(_5759_),
    .B(_5764_),
    .C(_5766_),
    .Y(_5777_)
);

AOI21X1 _16187_ (
    .A(_5777_),
    .B(_5776_),
    .C(_5775_),
    .Y(_5778_)
);

NOR2X1 _16188_ (
    .A(_5774_),
    .B(_5778_),
    .Y(_5779_)
);

OAI21X1 _16189_ (
    .A(_5434_),
    .B(_5432_),
    .C(_5423_),
    .Y(_5780_)
);

NAND2X1 _16190_ (
    .A(areg_11_bF$buf2),
    .B(breg_16_bF$buf2),
    .Y(_5781_)
);

OAI21X1 _16191_ (
    .A(_5406_),
    .B(_5781_),
    .C(_5415_),
    .Y(_5782_)
);

NAND2X1 _16192_ (
    .A(areg_10_bF$buf1),
    .B(breg_17_bF$buf3),
    .Y(_5783_)
);

INVX1 _16193_ (
    .A(_5783_),
    .Y(_5784_)
);

AND2X2 _16194_ (
    .A(areg_11_bF$buf1),
    .B(breg_16_bF$buf1),
    .Y(_5785_)
);

AND2X2 _16195_ (
    .A(areg_12_bF$buf2),
    .B(breg_15_bF$buf4),
    .Y(_5786_)
);

NAND2X1 _16196_ (
    .A(_5785_),
    .B(_5786_),
    .Y(_5787_)
);

OAI21X1 _16197_ (
    .A(_10869__bF$buf1),
    .B(_2362__bF$buf1),
    .C(_5781_),
    .Y(_5788_)
);

NAND3X1 _16198_ (
    .A(_5784_),
    .B(_5788_),
    .C(_5787_),
    .Y(_5789_)
);

OAI21X1 _16199_ (
    .A(_9104__bF$buf2),
    .B(_2560__bF$buf1),
    .C(_5786_),
    .Y(_5790_)
);

OAI21X1 _16200_ (
    .A(_10869__bF$buf0),
    .B(_2362__bF$buf0),
    .C(_5785_),
    .Y(_5791_)
);

NAND3X1 _16201_ (
    .A(_5783_),
    .B(_5790_),
    .C(_5791_),
    .Y(_5794_)
);

NAND2X1 _16202_ (
    .A(breg_12_bF$buf4),
    .B(areg_14_bF$buf4),
    .Y(_5795_)
);

AND2X2 _16203_ (
    .A(_5419_),
    .B(_5795_),
    .Y(_5796_)
);

OAI22X1 _16204_ (
    .A(_5106_),
    .B(_5468_),
    .C(_5796_),
    .D(_5466_),
    .Y(_5797_)
);

NAND3X1 _16205_ (
    .A(_5789_),
    .B(_5794_),
    .C(_5797_),
    .Y(_5798_)
);

AOI21X1 _16206_ (
    .A(_5790_),
    .B(_5791_),
    .C(_5783_),
    .Y(_5799_)
);

AOI21X1 _16207_ (
    .A(_5788_),
    .B(_5787_),
    .C(_5784_),
    .Y(_5800_)
);

NOR2X1 _16208_ (
    .A(_5419_),
    .B(_5795_),
    .Y(_5801_)
);

AOI21X1 _16209_ (
    .A(_5467_),
    .B(_5469_),
    .C(_5801_),
    .Y(_5802_)
);

OAI21X1 _16210_ (
    .A(_5799_),
    .B(_5800_),
    .C(_5802_),
    .Y(_5803_)
);

NAND3X1 _16211_ (
    .A(_5782_),
    .B(_5798_),
    .C(_5803_),
    .Y(_5805_)
);

AOI21X1 _16212_ (
    .A(_5048_),
    .B(_5785_),
    .C(_5424_),
    .Y(_5806_)
);

NOR3X1 _16213_ (
    .A(_5800_),
    .B(_5802_),
    .C(_5799_),
    .Y(_5807_)
);

AOI21X1 _16214_ (
    .A(_5789_),
    .B(_5794_),
    .C(_5797_),
    .Y(_5808_)
);

OAI21X1 _16215_ (
    .A(_5807_),
    .B(_5808_),
    .C(_5806_),
    .Y(_5809_)
);

NAND3X1 _16216_ (
    .A(_5805_),
    .B(_5780_),
    .C(_5809_),
    .Y(_5810_)
);

AOI21X1 _16217_ (
    .A(_5407_),
    .B(_5429_),
    .C(_5433_),
    .Y(_5811_)
);

NAND3X1 _16218_ (
    .A(_5802_),
    .B(_5789_),
    .C(_5794_),
    .Y(_5812_)
);

OAI21X1 _16219_ (
    .A(_5799_),
    .B(_5800_),
    .C(_5797_),
    .Y(_5813_)
);

AOI21X1 _16220_ (
    .A(_5812_),
    .B(_5813_),
    .C(_5806_),
    .Y(_5814_)
);

AOI21X1 _16221_ (
    .A(_5798_),
    .B(_5803_),
    .C(_5782_),
    .Y(_5816_)
);

OAI21X1 _16222_ (
    .A(_5814_),
    .B(_5816_),
    .C(_5811_),
    .Y(_5817_)
);

NAND3X1 _16223_ (
    .A(_5779_),
    .B(_5817_),
    .C(_5810_),
    .Y(_5818_)
);

OR2X2 _16224_ (
    .A(_5774_),
    .B(_5778_),
    .Y(_5819_)
);

OAI21X1 _16225_ (
    .A(_5814_),
    .B(_5816_),
    .C(_5780_),
    .Y(_5820_)
);

NAND3X1 _16226_ (
    .A(_5811_),
    .B(_5805_),
    .C(_5809_),
    .Y(_5821_)
);

NAND3X1 _16227_ (
    .A(_5820_),
    .B(_5821_),
    .C(_5819_),
    .Y(_5822_)
);

OAI21X1 _16228_ (
    .A(_5506_),
    .B(_5499_),
    .C(_5509_),
    .Y(_5823_)
);

AOI21X1 _16229_ (
    .A(_5818_),
    .B(_5822_),
    .C(_5823_),
    .Y(_5824_)
);

AOI21X1 _16230_ (
    .A(_5821_),
    .B(_5820_),
    .C(_5819_),
    .Y(_5825_)
);

AOI21X1 _16231_ (
    .A(_5817_),
    .B(_5810_),
    .C(_5779_),
    .Y(_5827_)
);

AOI21X1 _16232_ (
    .A(_5465_),
    .B(_5507_),
    .C(_5504_),
    .Y(_5828_)
);

NOR3X1 _16233_ (
    .A(_5825_),
    .B(_5827_),
    .C(_5828_),
    .Y(_5829_)
);

OAI21X1 _16234_ (
    .A(_5829_),
    .B(_5824_),
    .C(_5746_),
    .Y(_5830_)
);

AND2X2 _16235_ (
    .A(_5444_),
    .B(_5436_),
    .Y(_5831_)
);

OAI21X1 _16236_ (
    .A(_5825_),
    .B(_5827_),
    .C(_5828_),
    .Y(_5832_)
);

NAND3X1 _16237_ (
    .A(_5818_),
    .B(_5823_),
    .C(_5822_),
    .Y(_5833_)
);

NAND3X1 _16238_ (
    .A(_5832_),
    .B(_5833_),
    .C(_5831_),
    .Y(_5834_)
);

NAND2X1 _16239_ (
    .A(_5834_),
    .B(_5830_),
    .Y(_5835_)
);

AOI21X1 _16240_ (
    .A(_5584_),
    .B(_5591_),
    .C(_5513_),
    .Y(_5836_)
);

OAI21X1 _16241_ (
    .A(_5602_),
    .B(_5836_),
    .C(_5592_),
    .Y(_5838_)
);

NAND2X1 _16242_ (
    .A(_5485_),
    .B(_5491_),
    .Y(_5839_)
);

NAND2X1 _16243_ (
    .A(areg_13_bF$buf0),
    .B(breg_14_bF$buf3),
    .Y(_5840_)
);

INVX2 _16244_ (
    .A(_5840_),
    .Y(_5841_)
);

NAND2X1 _16245_ (
    .A(breg_13_bF$buf4),
    .B(areg_15_bF$buf2),
    .Y(_5842_)
);

OAI21X1 _16246_ (
    .A(_2586__bF$buf3),
    .B(_2465__bF$buf4),
    .C(_5468_),
    .Y(_5843_)
);

OAI21X1 _16247_ (
    .A(_5795_),
    .B(_5842_),
    .C(_5843_),
    .Y(_5844_)
);

XNOR2X1 _16248_ (
    .A(_5844_),
    .B(_5841_),
    .Y(_5845_)
);

OAI21X1 _16249_ (
    .A(_5483_),
    .B(_5473_),
    .C(_5477_),
    .Y(_5846_)
);

NAND2X1 _16250_ (
    .A(breg_11_bF$buf0),
    .B(areg_16_bF$buf4),
    .Y(_5847_)
);

INVX2 _16251_ (
    .A(_5847_),
    .Y(_5849_)
);

AND2X2 _16252_ (
    .A(breg_9_bF$buf3),
    .B(areg_18_bF$buf4),
    .Y(_5850_)
);

NAND2X1 _16253_ (
    .A(_5476_),
    .B(_5850_),
    .Y(_5851_)
);

OAI22X1 _16254_ (
    .A(_6044__bF$buf2),
    .B(_3146__bF$buf3),
    .C(_7217__bF$buf4),
    .D(_2884__bF$buf0),
    .Y(_5852_)
);

NAND3X1 _16255_ (
    .A(_5849_),
    .B(_5852_),
    .C(_5851_),
    .Y(_5853_)
);

NAND2X1 _16256_ (
    .A(breg_10_bF$buf5),
    .B(areg_18_bF$buf3),
    .Y(_5854_)
);

NOR2X1 _16257_ (
    .A(_5481_),
    .B(_5854_),
    .Y(_5855_)
);

NOR2X1 _16258_ (
    .A(_5476_),
    .B(_5850_),
    .Y(_5856_)
);

OAI21X1 _16259_ (
    .A(_5856_),
    .B(_5855_),
    .C(_5847_),
    .Y(_5857_)
);

NAND3X1 _16260_ (
    .A(_5846_),
    .B(_5853_),
    .C(_5857_),
    .Y(_5858_)
);

AOI21X1 _16261_ (
    .A(_5474_),
    .B(_5479_),
    .C(_5482_),
    .Y(_5860_)
);

OAI21X1 _16262_ (
    .A(_7217__bF$buf3),
    .B(_2884__bF$buf3),
    .C(_5850_),
    .Y(_5861_)
);

OAI21X1 _16263_ (
    .A(_6044__bF$buf1),
    .B(_3146__bF$buf2),
    .C(_5476_),
    .Y(_5862_)
);

AOI21X1 _16264_ (
    .A(_5861_),
    .B(_5862_),
    .C(_5847_),
    .Y(_5863_)
);

AOI21X1 _16265_ (
    .A(_5852_),
    .B(_5851_),
    .C(_5849_),
    .Y(_5864_)
);

OAI21X1 _16266_ (
    .A(_5863_),
    .B(_5864_),
    .C(_5860_),
    .Y(_5865_)
);

NAND3X1 _16267_ (
    .A(_5858_),
    .B(_5865_),
    .C(_5845_),
    .Y(_5866_)
);

XNOR2X1 _16268_ (
    .A(_5844_),
    .B(_5840_),
    .Y(_5867_)
);

OAI21X1 _16269_ (
    .A(_5863_),
    .B(_5864_),
    .C(_5846_),
    .Y(_5868_)
);

NAND3X1 _16270_ (
    .A(_5860_),
    .B(_5853_),
    .C(_5857_),
    .Y(_5869_)
);

NAND3X1 _16271_ (
    .A(_5868_),
    .B(_5869_),
    .C(_5867_),
    .Y(_5871_)
);

OAI21X1 _16272_ (
    .A(_5529_),
    .B(_5535_),
    .C(_5537_),
    .Y(_5872_)
);

AOI21X1 _16273_ (
    .A(_5871_),
    .B(_5866_),
    .C(_5872_),
    .Y(_5873_)
);

AOI21X1 _16274_ (
    .A(_5868_),
    .B(_5869_),
    .C(_5867_),
    .Y(_5874_)
);

AOI21X1 _16275_ (
    .A(_5865_),
    .B(_5858_),
    .C(_5845_),
    .Y(_5875_)
);

AOI21X1 _16276_ (
    .A(_5515_),
    .B(_5536_),
    .C(_5533_),
    .Y(_5876_)
);

NOR3X1 _16277_ (
    .A(_5874_),
    .B(_5875_),
    .C(_5876_),
    .Y(_5877_)
);

OAI21X1 _16278_ (
    .A(_5877_),
    .B(_5873_),
    .C(_5839_),
    .Y(_5878_)
);

AND2X2 _16279_ (
    .A(_5491_),
    .B(_5485_),
    .Y(_5879_)
);

OAI21X1 _16280_ (
    .A(_5874_),
    .B(_5875_),
    .C(_5876_),
    .Y(_5880_)
);

NAND3X1 _16281_ (
    .A(_5866_),
    .B(_5871_),
    .C(_5872_),
    .Y(_5882_)
);

NAND3X1 _16282_ (
    .A(_5879_),
    .B(_5880_),
    .C(_5882_),
    .Y(_5883_)
);

NAND2X1 _16283_ (
    .A(_5883_),
    .B(_5878_),
    .Y(_5884_)
);

AOI21X1 _16284_ (
    .A(_5577_),
    .B(_5572_),
    .C(_5542_),
    .Y(_5885_)
);

OAI21X1 _16285_ (
    .A(_5588_),
    .B(_5885_),
    .C(_5578_),
    .Y(_5886_)
);

NAND2X1 _16286_ (
    .A(breg_7_bF$buf3),
    .B(areg_20_bF$buf4),
    .Y(_5887_)
);

OAI21X1 _16287_ (
    .A(_5514_),
    .B(_5887_),
    .C(_5522_),
    .Y(_5888_)
);

NAND2X1 _16288_ (
    .A(breg[8]),
    .B(areg_19_bF$buf5),
    .Y(_5889_)
);

INVX1 _16289_ (
    .A(_5889_),
    .Y(_5890_)
);

AND2X2 _16290_ (
    .A(breg_7_bF$buf2),
    .B(areg_20_bF$buf3),
    .Y(_5891_)
);

AND2X2 _16291_ (
    .A(breg_6_bF$buf0),
    .B(areg_21_bF$buf0),
    .Y(_5893_)
);

NAND2X1 _16292_ (
    .A(_5891_),
    .B(_5893_),
    .Y(_5894_)
);

OAI21X1 _16293_ (
    .A(_5453__bF$buf3),
    .B(_3961__bF$buf2),
    .C(_5887_),
    .Y(_5895_)
);

NAND3X1 _16294_ (
    .A(_5890_),
    .B(_5895_),
    .C(_5894_),
    .Y(_5896_)
);

OAI21X1 _16295_ (
    .A(_4116__bF$buf4),
    .B(_3958__bF$buf3),
    .C(_5893_),
    .Y(_5897_)
);

OAI21X1 _16296_ (
    .A(_5453__bF$buf2),
    .B(_3961__bF$buf1),
    .C(_5891_),
    .Y(_5898_)
);

NAND3X1 _16297_ (
    .A(_5889_),
    .B(_5897_),
    .C(_5898_),
    .Y(_5899_)
);

OAI21X1 _16298_ (
    .A(_5551_),
    .B(_5543_),
    .C(_5547_),
    .Y(_5900_)
);

AOI21X1 _16299_ (
    .A(_5896_),
    .B(_5899_),
    .C(_5900_),
    .Y(_5901_)
);

AOI21X1 _16300_ (
    .A(_5897_),
    .B(_5898_),
    .C(_5889_),
    .Y(_5902_)
);

AOI21X1 _16301_ (
    .A(_5895_),
    .B(_5894_),
    .C(_5890_),
    .Y(_5904_)
);

AOI21X1 _16302_ (
    .A(_5544_),
    .B(_5548_),
    .C(_5550_),
    .Y(_5905_)
);

NOR3X1 _16303_ (
    .A(_5904_),
    .B(_5905_),
    .C(_5902_),
    .Y(_5906_)
);

OAI21X1 _16304_ (
    .A(_5906_),
    .B(_5901_),
    .C(_5888_),
    .Y(_5907_)
);

INVX2 _16305_ (
    .A(_5888_),
    .Y(_5908_)
);

OAI21X1 _16306_ (
    .A(_5902_),
    .B(_5904_),
    .C(_5905_),
    .Y(_5909_)
);

NAND3X1 _16307_ (
    .A(_5896_),
    .B(_5899_),
    .C(_5900_),
    .Y(_5910_)
);

NAND3X1 _16308_ (
    .A(_5909_),
    .B(_5910_),
    .C(_5908_),
    .Y(_5911_)
);

NAND2X1 _16309_ (
    .A(_5907_),
    .B(_5911_),
    .Y(_5912_)
);

AOI21X1 _16310_ (
    .A(_5566_),
    .B(_5562_),
    .C(_5555_),
    .Y(_5913_)
);

OAI21X1 _16311_ (
    .A(_5913_),
    .B(_5573_),
    .C(_5567_),
    .Y(_5915_)
);

NAND2X1 _16312_ (
    .A(breg_5_bF$buf2),
    .B(areg_22_bF$buf2),
    .Y(_5916_)
);

INVX1 _16313_ (
    .A(_5916_),
    .Y(_5917_)
);

NAND2X1 _16314_ (
    .A(breg_4_bF$buf5),
    .B(areg_23_bF$buf3),
    .Y(_5918_)
);

NAND2X1 _16315_ (
    .A(breg_3_bF$buf1),
    .B(areg_24_bF$buf4),
    .Y(_5919_)
);

OR2X2 _16316_ (
    .A(_5918_),
    .B(_5919_),
    .Y(_5920_)
);

INVX8 _16317_ (
    .A(areg_24_bF$buf3),
    .Y(_5921_)
);

OAI21X1 _16318_ (
    .A(_2365_),
    .B(_5921__bF$buf3),
    .C(_5918_),
    .Y(_5922_)
);

NAND3X1 _16319_ (
    .A(_5917_),
    .B(_5922_),
    .C(_5920_),
    .Y(_5923_)
);

NOR2X1 _16320_ (
    .A(_5918_),
    .B(_5919_),
    .Y(_5924_)
);

AND2X2 _16321_ (
    .A(_5918_),
    .B(_5919_),
    .Y(_5926_)
);

OAI21X1 _16322_ (
    .A(_5926_),
    .B(_5924_),
    .C(_5916_),
    .Y(_5927_)
);

AND2X2 _16323_ (
    .A(_5923_),
    .B(_5927_),
    .Y(_5928_)
);

OAI21X1 _16324_ (
    .A(_5556_),
    .B(_5560_),
    .C(_5559_),
    .Y(_5929_)
);

NAND2X1 _16325_ (
    .A(breg_2_bF$buf1),
    .B(areg_25_bF$buf0),
    .Y(_5930_)
);

INVX2 _16326_ (
    .A(_5930_),
    .Y(_5931_)
);

AND2X2 _16327_ (
    .A(breg_0_bF$buf0),
    .B(areg_27_bF$buf5),
    .Y(_5932_)
);

NAND2X1 _16328_ (
    .A(_5558_),
    .B(_5932_),
    .Y(_5933_)
);

AOI22X1 _16329_ (
    .A(breg_0_bF$buf6),
    .B(areg_27_bF$buf4),
    .C(breg_1_bF$buf6),
    .D(areg_26_bF$buf1),
    .Y(_5934_)
);

INVX2 _16330_ (
    .A(_5934_),
    .Y(_5935_)
);

NAND3X1 _16331_ (
    .A(_5931_),
    .B(_5935_),
    .C(_5933_),
    .Y(_5937_)
);

NAND2X1 _16332_ (
    .A(breg_0_bF$buf5),
    .B(areg_27_bF$buf3),
    .Y(_5938_)
);

NOR2X1 _16333_ (
    .A(_5564_),
    .B(_5938_),
    .Y(_5939_)
);

OAI21X1 _16334_ (
    .A(_5939_),
    .B(_5934_),
    .C(_5930_),
    .Y(_5940_)
);

NAND3X1 _16335_ (
    .A(_5929_),
    .B(_5940_),
    .C(_5937_),
    .Y(_5941_)
);

AOI21X1 _16336_ (
    .A(_5557_),
    .B(_5561_),
    .C(_5565_),
    .Y(_5942_)
);

NAND2X1 _16337_ (
    .A(_5564_),
    .B(_5932_),
    .Y(_5943_)
);

NAND2X1 _16338_ (
    .A(_5938_),
    .B(_5558_),
    .Y(_5944_)
);

AOI21X1 _16339_ (
    .A(_5943_),
    .B(_5944_),
    .C(_5930_),
    .Y(_5945_)
);

AOI21X1 _16340_ (
    .A(_5935_),
    .B(_5933_),
    .C(_5931_),
    .Y(_5946_)
);

OAI21X1 _16341_ (
    .A(_5946_),
    .B(_5945_),
    .C(_5942_),
    .Y(_5948_)
);

NAND3X1 _16342_ (
    .A(_5941_),
    .B(_5948_),
    .C(_5928_),
    .Y(_5949_)
);

NAND2X1 _16343_ (
    .A(_5927_),
    .B(_5923_),
    .Y(_5950_)
);

OAI21X1 _16344_ (
    .A(_5946_),
    .B(_5945_),
    .C(_5929_),
    .Y(_5951_)
);

NAND3X1 _16345_ (
    .A(_5940_),
    .B(_5942_),
    .C(_5937_),
    .Y(_5952_)
);

NAND3X1 _16346_ (
    .A(_5950_),
    .B(_5952_),
    .C(_5951_),
    .Y(_5953_)
);

NAND3X1 _16347_ (
    .A(_5915_),
    .B(_5953_),
    .C(_5949_),
    .Y(_5954_)
);

NOR3X1 _16348_ (
    .A(_5569_),
    .B(_5568_),
    .C(_5570_),
    .Y(_5955_)
);

AOI21X1 _16349_ (
    .A(_5554_),
    .B(_5571_),
    .C(_5955_),
    .Y(_5956_)
);

AOI21X1 _16350_ (
    .A(_5952_),
    .B(_5951_),
    .C(_5950_),
    .Y(_5957_)
);

AOI21X1 _16351_ (
    .A(_5941_),
    .B(_5948_),
    .C(_5928_),
    .Y(_5959_)
);

OAI21X1 _16352_ (
    .A(_5957_),
    .B(_5959_),
    .C(_5956_),
    .Y(_5960_)
);

NAND3X1 _16353_ (
    .A(_5954_),
    .B(_5912_),
    .C(_5960_),
    .Y(_5961_)
);

NAND3X1 _16354_ (
    .A(_5888_),
    .B(_5910_),
    .C(_5909_),
    .Y(_5962_)
);

OAI21X1 _16355_ (
    .A(_5906_),
    .B(_5901_),
    .C(_5908_),
    .Y(_5963_)
);

NAND2X1 _16356_ (
    .A(_5962_),
    .B(_5963_),
    .Y(_5964_)
);

OAI21X1 _16357_ (
    .A(_5957_),
    .B(_5959_),
    .C(_5915_),
    .Y(_5965_)
);

NAND3X1 _16358_ (
    .A(_5949_),
    .B(_5953_),
    .C(_5956_),
    .Y(_5966_)
);

NAND3X1 _16359_ (
    .A(_5964_),
    .B(_5966_),
    .C(_5965_),
    .Y(_5967_)
);

NAND3X1 _16360_ (
    .A(_5961_),
    .B(_5967_),
    .C(_5886_),
    .Y(_5968_)
);

NOR3X1 _16361_ (
    .A(_5581_),
    .B(_5582_),
    .C(_5580_),
    .Y(_5970_)
);

AOI21X1 _16362_ (
    .A(_5539_),
    .B(_5583_),
    .C(_5970_),
    .Y(_5971_)
);

AOI21X1 _16363_ (
    .A(_5966_),
    .B(_5965_),
    .C(_5964_),
    .Y(_5972_)
);

AOI21X1 _16364_ (
    .A(_5954_),
    .B(_5960_),
    .C(_5912_),
    .Y(_5973_)
);

OAI21X1 _16365_ (
    .A(_5972_),
    .B(_5973_),
    .C(_5971_),
    .Y(_5974_)
);

NAND3X1 _16366_ (
    .A(_5968_),
    .B(_5884_),
    .C(_5974_),
    .Y(_5975_)
);

NAND3X1 _16367_ (
    .A(_5839_),
    .B(_5880_),
    .C(_5882_),
    .Y(_5976_)
);

OAI21X1 _16368_ (
    .A(_5877_),
    .B(_5873_),
    .C(_5879_),
    .Y(_5977_)
);

NAND2X1 _16369_ (
    .A(_5976_),
    .B(_5977_),
    .Y(_5978_)
);

OAI21X1 _16370_ (
    .A(_5972_),
    .B(_5973_),
    .C(_5886_),
    .Y(_5979_)
);

NAND3X1 _16371_ (
    .A(_5961_),
    .B(_5967_),
    .C(_5971_),
    .Y(_5980_)
);

NAND3X1 _16372_ (
    .A(_5978_),
    .B(_5979_),
    .C(_5980_),
    .Y(_5981_)
);

NAND3X1 _16373_ (
    .A(_5975_),
    .B(_5981_),
    .C(_5838_),
    .Y(_5982_)
);

NOR3X1 _16374_ (
    .A(_5595_),
    .B(_5597_),
    .C(_5594_),
    .Y(_5983_)
);

AOI21X1 _16375_ (
    .A(_5511_),
    .B(_5598_),
    .C(_5983_),
    .Y(_5984_)
);

AOI21X1 _16376_ (
    .A(_5979_),
    .B(_5980_),
    .C(_5978_),
    .Y(_5985_)
);

AOI21X1 _16377_ (
    .A(_5968_),
    .B(_5974_),
    .C(_5884_),
    .Y(_5986_)
);

OAI21X1 _16378_ (
    .A(_5985_),
    .B(_5986_),
    .C(_5984_),
    .Y(_5987_)
);

NAND3X1 _16379_ (
    .A(_5982_),
    .B(_5987_),
    .C(_5835_),
    .Y(_5988_)
);

NAND3X1 _16380_ (
    .A(_5746_),
    .B(_5833_),
    .C(_5832_),
    .Y(_5989_)
);

OAI21X1 _16381_ (
    .A(_5829_),
    .B(_5824_),
    .C(_5831_),
    .Y(_5991_)
);

NAND2X1 _16382_ (
    .A(_5989_),
    .B(_5991_),
    .Y(_5992_)
);

OAI21X1 _16383_ (
    .A(_5985_),
    .B(_5986_),
    .C(_5838_),
    .Y(_5993_)
);

NAND3X1 _16384_ (
    .A(_5975_),
    .B(_5981_),
    .C(_5984_),
    .Y(_5994_)
);

NAND3X1 _16385_ (
    .A(_5993_),
    .B(_5992_),
    .C(_5994_),
    .Y(_5995_)
);

NAND3X1 _16386_ (
    .A(_5988_),
    .B(_5995_),
    .C(_5745_),
    .Y(_5996_)
);

NOR3X1 _16387_ (
    .A(_5610_),
    .B(_5611_),
    .C(_5609_),
    .Y(_5997_)
);

AOI21X1 _16388_ (
    .A(_5612_),
    .B(_5461_),
    .C(_5997_),
    .Y(_5998_)
);

AOI21X1 _16389_ (
    .A(_5993_),
    .B(_5994_),
    .C(_5992_),
    .Y(_5999_)
);

AOI21X1 _16390_ (
    .A(_5982_),
    .B(_5987_),
    .C(_5835_),
    .Y(_6000_)
);

OAI21X1 _16391_ (
    .A(_5999_),
    .B(_6000_),
    .C(_5998_),
    .Y(_6002_)
);

NAND3X1 _16392_ (
    .A(_5996_),
    .B(_5743_),
    .C(_6002_),
    .Y(_6003_)
);

NAND3X1 _16393_ (
    .A(_5739_),
    .B(_5732_),
    .C(_5736_),
    .Y(_6004_)
);

NAND3X1 _16394_ (
    .A(_5352_),
    .B(_5740_),
    .C(_5741_),
    .Y(_6005_)
);

NAND2X1 _16395_ (
    .A(_6004_),
    .B(_6005_),
    .Y(_6006_)
);

OAI21X1 _16396_ (
    .A(_5999_),
    .B(_6000_),
    .C(_5745_),
    .Y(_6007_)
);

NAND3X1 _16397_ (
    .A(_5988_),
    .B(_5995_),
    .C(_5998_),
    .Y(_6008_)
);

NAND3X1 _16398_ (
    .A(_6007_),
    .B(_6006_),
    .C(_6008_),
    .Y(_6009_)
);

NAND3X1 _16399_ (
    .A(_6003_),
    .B(_5667_),
    .C(_6009_),
    .Y(_6010_)
);

AOI21X1 _16400_ (
    .A(_5366_),
    .B(_5625_),
    .C(_5631_),
    .Y(_6011_)
);

AOI21X1 _16401_ (
    .A(_6007_),
    .B(_6008_),
    .C(_6006_),
    .Y(_6013_)
);

AOI21X1 _16402_ (
    .A(_5996_),
    .B(_6002_),
    .C(_5743_),
    .Y(_6014_)
);

OAI21X1 _16403_ (
    .A(_6013_),
    .B(_6014_),
    .C(_6011_),
    .Y(_6015_)
);

NAND3X1 _16404_ (
    .A(_5666_),
    .B(_6010_),
    .C(_6015_),
    .Y(_6016_)
);

INVX2 _16405_ (
    .A(_5666_),
    .Y(_6017_)
);

NOR3X1 _16406_ (
    .A(_6013_),
    .B(_6014_),
    .C(_6011_),
    .Y(_6018_)
);

AOI21X1 _16407_ (
    .A(_6003_),
    .B(_6009_),
    .C(_5667_),
    .Y(_6019_)
);

OAI21X1 _16408_ (
    .A(_6018_),
    .B(_6019_),
    .C(_6017_),
    .Y(_6020_)
);

NAND3X1 _16409_ (
    .A(_6016_),
    .B(_5665_),
    .C(_6020_),
    .Y(_6021_)
);

AOI21X1 _16410_ (
    .A(_5306_),
    .B(_5641_),
    .C(_5643_),
    .Y(_6022_)
);

OAI21X1 _16411_ (
    .A(_6013_),
    .B(_6014_),
    .C(_5667_),
    .Y(_6024_)
);

NAND3X1 _16412_ (
    .A(_6003_),
    .B(_6009_),
    .C(_6011_),
    .Y(_6025_)
);

AOI21X1 _16413_ (
    .A(_6024_),
    .B(_6025_),
    .C(_6017_),
    .Y(_6026_)
);

AOI21X1 _16414_ (
    .A(_6010_),
    .B(_6015_),
    .C(_5666_),
    .Y(_6027_)
);

OAI21X1 _16415_ (
    .A(_6026_),
    .B(_6027_),
    .C(_6022_),
    .Y(_6028_)
);

NAND3X1 _16416_ (
    .A(_6021_),
    .B(_6028_),
    .C(_5664_),
    .Y(_6029_)
);

NOR3X1 _16417_ (
    .A(_6026_),
    .B(_6027_),
    .C(_6022_),
    .Y(_6030_)
);

AOI21X1 _16418_ (
    .A(_6016_),
    .B(_6020_),
    .C(_5665_),
    .Y(_6031_)
);

OAI21X1 _16419_ (
    .A(_6030_),
    .B(_6031_),
    .C(_5646_),
    .Y(_6032_)
);

NAND2X1 _16420_ (
    .A(_6032_),
    .B(_6029_),
    .Y(_6033_)
);

XNOR2X1 _16421_ (
    .A(_5663_),
    .B(_6033_),
    .Y(_0_[27])
);

NAND3X1 _16422_ (
    .A(_6029_),
    .B(_6032_),
    .C(_5658_),
    .Y(_6035_)
);

NAND2X1 _16423_ (
    .A(_6032_),
    .B(_5659_),
    .Y(_6036_)
);

AND2X2 _16424_ (
    .A(_6036_),
    .B(_6029_),
    .Y(_6037_)
);

OAI21X1 _16425_ (
    .A(_6035_),
    .B(_5298_),
    .C(_6037_),
    .Y(_6038_)
);

AOI21X1 _16426_ (
    .A(_5654_),
    .B(_5657_),
    .C(_6033_),
    .Y(_6039_)
);

NAND2X1 _16427_ (
    .A(_5301_),
    .B(_6039_),
    .Y(_6040_)
);

NOR2X1 _16428_ (
    .A(_6040_),
    .B(_4962_),
    .Y(_6041_)
);

NOR2X1 _16429_ (
    .A(_6038_),
    .B(_6041_),
    .Y(_6042_)
);

OAI21X1 _16430_ (
    .A(_6019_),
    .B(_6017_),
    .C(_6010_),
    .Y(_6043_)
);

NAND2X1 _16431_ (
    .A(_5732_),
    .B(_6004_),
    .Y(_6045_)
);

AOI21X1 _16432_ (
    .A(_5988_),
    .B(_5995_),
    .C(_5745_),
    .Y(_6046_)
);

OAI21X1 _16433_ (
    .A(_6006_),
    .B(_6046_),
    .C(_5996_),
    .Y(_6047_)
);

AND2X2 _16434_ (
    .A(_5725_),
    .B(_5718_),
    .Y(_6048_)
);

NAND2X1 _16435_ (
    .A(areg_1_bF$buf4),
    .B(breg_28_bF$buf5),
    .Y(_6049_)
);

INVX8 _16436_ (
    .A(breg_28_bF$buf4),
    .Y(_6050_)
);

NAND2X1 _16437_ (
    .A(areg_1_bF$buf3),
    .B(breg_27_bF$buf4),
    .Y(_6051_)
);

OAI21X1 _16438_ (
    .A(_2376__bF$buf0),
    .B(_6050__bF$buf3),
    .C(_6051_),
    .Y(_6052_)
);

OAI21X1 _16439_ (
    .A(_5726_),
    .B(_6049_),
    .C(_6052_),
    .Y(_6053_)
);

INVX1 _16440_ (
    .A(_6053_),
    .Y(_6054_)
);

AOI21X1 _16441_ (
    .A(_5700_),
    .B(_5704_),
    .C(_5706_),
    .Y(_6056_)
);

OAI21X1 _16442_ (
    .A(_5713_),
    .B(_6056_),
    .C(_5707_),
    .Y(_6057_)
);

NAND2X1 _16443_ (
    .A(_5690_),
    .B(_5700_),
    .Y(_6058_)
);

OAI21X1 _16444_ (
    .A(_5686_),
    .B(_5691_),
    .C(_5680_),
    .Y(_6059_)
);

NAND2X1 _16445_ (
    .A(areg_2_bF$buf1),
    .B(breg_26_bF$buf2),
    .Y(_6060_)
);

INVX1 _16446_ (
    .A(_6060_),
    .Y(_6061_)
);

AND2X2 _16447_ (
    .A(areg_3_bF$buf1),
    .B(breg_25_bF$buf4),
    .Y(_6062_)
);

AND2X2 _16448_ (
    .A(areg_4_bF$buf0),
    .B(breg_24_bF$buf5),
    .Y(_6063_)
);

NAND2X1 _16449_ (
    .A(_6062_),
    .B(_6063_),
    .Y(_6064_)
);

OAI21X1 _16450_ (
    .A(_2562__bF$buf2),
    .B(_5315__bF$buf0),
    .C(_5685_),
    .Y(_6065_)
);

NAND3X1 _16451_ (
    .A(_6061_),
    .B(_6065_),
    .C(_6064_),
    .Y(_6066_)
);

OAI21X1 _16452_ (
    .A(_2792_),
    .B(_5318_),
    .C(_6063_),
    .Y(_6067_)
);

OAI21X1 _16453_ (
    .A(_2562__bF$buf1),
    .B(_5315__bF$buf4),
    .C(_6062_),
    .Y(_6068_)
);

NAND3X1 _16454_ (
    .A(_6060_),
    .B(_6067_),
    .C(_6068_),
    .Y(_6069_)
);

NAND2X1 _16455_ (
    .A(areg_6_bF$buf4),
    .B(breg_22_bF$buf3),
    .Y(_6070_)
);

AND2X2 _16456_ (
    .A(_5688_),
    .B(_5750_),
    .Y(_6071_)
);

OAI22X1 _16457_ (
    .A(_5373_),
    .B(_6070_),
    .C(_6071_),
    .D(_5747_),
    .Y(_6072_)
);

NAND3X1 _16458_ (
    .A(_6066_),
    .B(_6069_),
    .C(_6072_),
    .Y(_6073_)
);

AOI21X1 _16459_ (
    .A(_6067_),
    .B(_6068_),
    .C(_6060_),
    .Y(_6074_)
);

AOI21X1 _16460_ (
    .A(_6065_),
    .B(_6064_),
    .C(_6061_),
    .Y(_6075_)
);

NOR2X1 _16461_ (
    .A(_5688_),
    .B(_5750_),
    .Y(_6077_)
);

OAI21X1 _16462_ (
    .A(_3646__bF$buf2),
    .B(_3781__bF$buf3),
    .C(_5688_),
    .Y(_6078_)
);

AOI21X1 _16463_ (
    .A(_5748_),
    .B(_6078_),
    .C(_6077_),
    .Y(_6079_)
);

OAI21X1 _16464_ (
    .A(_6074_),
    .B(_6075_),
    .C(_6079_),
    .Y(_6080_)
);

NAND3X1 _16465_ (
    .A(_6059_),
    .B(_6073_),
    .C(_6080_),
    .Y(_6081_)
);

INVX1 _16466_ (
    .A(_6059_),
    .Y(_6082_)
);

NAND3X1 _16467_ (
    .A(_6079_),
    .B(_6066_),
    .C(_6069_),
    .Y(_6083_)
);

OAI21X1 _16468_ (
    .A(_6074_),
    .B(_6075_),
    .C(_6072_),
    .Y(_6084_)
);

NAND3X1 _16469_ (
    .A(_6083_),
    .B(_6084_),
    .C(_6082_),
    .Y(_6085_)
);

AOI21X1 _16470_ (
    .A(_5767_),
    .B(_5772_),
    .C(_5753_),
    .Y(_6086_)
);

OAI21X1 _16471_ (
    .A(_5752_),
    .B(_6086_),
    .C(_5776_),
    .Y(_6089_)
);

NAND3X1 _16472_ (
    .A(_6081_),
    .B(_6085_),
    .C(_6089_),
    .Y(_6090_)
);

AOI21X1 _16473_ (
    .A(_6083_),
    .B(_6084_),
    .C(_6082_),
    .Y(_6091_)
);

AOI21X1 _16474_ (
    .A(_6073_),
    .B(_6080_),
    .C(_6059_),
    .Y(_6092_)
);

NOR3X1 _16475_ (
    .A(_5764_),
    .B(_5766_),
    .C(_5759_),
    .Y(_6093_)
);

AOI21X1 _16476_ (
    .A(_5777_),
    .B(_5775_),
    .C(_6093_),
    .Y(_6094_)
);

OAI21X1 _16477_ (
    .A(_6091_),
    .B(_6092_),
    .C(_6094_),
    .Y(_6095_)
);

NAND3X1 _16478_ (
    .A(_6058_),
    .B(_6095_),
    .C(_6090_),
    .Y(_6096_)
);

AND2X2 _16479_ (
    .A(_5700_),
    .B(_5690_),
    .Y(_6097_)
);

NOR3X1 _16480_ (
    .A(_6091_),
    .B(_6092_),
    .C(_6094_),
    .Y(_6098_)
);

AOI21X1 _16481_ (
    .A(_6081_),
    .B(_6085_),
    .C(_6089_),
    .Y(_6100_)
);

OAI21X1 _16482_ (
    .A(_6098_),
    .B(_6100_),
    .C(_6097_),
    .Y(_6101_)
);

NAND3X1 _16483_ (
    .A(_6096_),
    .B(_6057_),
    .C(_6101_),
    .Y(_6102_)
);

NOR3X1 _16484_ (
    .A(_5708_),
    .B(_5709_),
    .C(_5710_),
    .Y(_6103_)
);

AOI21X1 _16485_ (
    .A(_5673_),
    .B(_5711_),
    .C(_6103_),
    .Y(_6104_)
);

NAND3X1 _16486_ (
    .A(_6081_),
    .B(_6085_),
    .C(_6094_),
    .Y(_6105_)
);

OAI21X1 _16487_ (
    .A(_6091_),
    .B(_6092_),
    .C(_6089_),
    .Y(_6106_)
);

AOI21X1 _16488_ (
    .A(_6106_),
    .B(_6105_),
    .C(_6097_),
    .Y(_6107_)
);

AOI21X1 _16489_ (
    .A(_6095_),
    .B(_6090_),
    .C(_6058_),
    .Y(_6108_)
);

OAI21X1 _16490_ (
    .A(_6108_),
    .B(_6107_),
    .C(_6104_),
    .Y(_6109_)
);

NAND3X1 _16491_ (
    .A(_6054_),
    .B(_6109_),
    .C(_6102_),
    .Y(_6111_)
);

OAI21X1 _16492_ (
    .A(_6107_),
    .B(_6108_),
    .C(_6057_),
    .Y(_6112_)
);

NAND3X1 _16493_ (
    .A(_6096_),
    .B(_6101_),
    .C(_6104_),
    .Y(_6113_)
);

NAND3X1 _16494_ (
    .A(_6053_),
    .B(_6112_),
    .C(_6113_),
    .Y(_6114_)
);

AOI21X1 _16495_ (
    .A(_5746_),
    .B(_5832_),
    .C(_5829_),
    .Y(_6115_)
);

NAND3X1 _16496_ (
    .A(_6111_),
    .B(_6115_),
    .C(_6114_),
    .Y(_6116_)
);

AOI21X1 _16497_ (
    .A(_6112_),
    .B(_6113_),
    .C(_6053_),
    .Y(_6117_)
);

AOI21X1 _16498_ (
    .A(_6109_),
    .B(_6102_),
    .C(_6054_),
    .Y(_6118_)
);

OAI21X1 _16499_ (
    .A(_5831_),
    .B(_5824_),
    .C(_5833_),
    .Y(_6119_)
);

OAI21X1 _16500_ (
    .A(_6117_),
    .B(_6118_),
    .C(_6119_),
    .Y(_6120_)
);

AOI21X1 _16501_ (
    .A(_6116_),
    .B(_6120_),
    .C(_6048_),
    .Y(_6122_)
);

NAND2X1 _16502_ (
    .A(_5718_),
    .B(_5725_),
    .Y(_6123_)
);

NAND3X1 _16503_ (
    .A(_6111_),
    .B(_6119_),
    .C(_6114_),
    .Y(_6124_)
);

OAI21X1 _16504_ (
    .A(_6117_),
    .B(_6118_),
    .C(_6115_),
    .Y(_6125_)
);

AOI21X1 _16505_ (
    .A(_6124_),
    .B(_6125_),
    .C(_6123_),
    .Y(_6126_)
);

NOR2X1 _16506_ (
    .A(_6122_),
    .B(_6126_),
    .Y(_6127_)
);

AOI21X1 _16507_ (
    .A(_5975_),
    .B(_5981_),
    .C(_5838_),
    .Y(_6128_)
);

OAI21X1 _16508_ (
    .A(_5992_),
    .B(_6128_),
    .C(_5982_),
    .Y(_6129_)
);

NAND2X1 _16509_ (
    .A(_5810_),
    .B(_5818_),
    .Y(_6130_)
);

NAND2X1 _16510_ (
    .A(areg_5_bF$buf4),
    .B(breg_23_bF$buf1),
    .Y(_6131_)
);

INVX2 _16511_ (
    .A(_6131_),
    .Y(_6133_)
);

NAND2X1 _16512_ (
    .A(areg_7_bF$buf0),
    .B(breg_21_bF$buf3),
    .Y(_6134_)
);

XOR2X1 _16513_ (
    .A(_6070_),
    .B(_6134_),
    .Y(_6135_)
);

XNOR2X1 _16514_ (
    .A(_6135_),
    .B(_6133_),
    .Y(_6136_)
);

OAI21X1 _16515_ (
    .A(_5770_),
    .B(_5754_),
    .C(_5762_),
    .Y(_6137_)
);

NAND2X1 _16516_ (
    .A(areg_8_bF$buf4),
    .B(breg_20_bF$buf2),
    .Y(_6138_)
);

NAND2X1 _16517_ (
    .A(areg_10_bF$buf0),
    .B(breg_18_bF$buf0),
    .Y(_6139_)
);

NOR2X1 _16518_ (
    .A(_5768_),
    .B(_6139_),
    .Y(_6140_)
);

AND2X2 _16519_ (
    .A(areg_9_bF$buf3),
    .B(breg_19_bF$buf0),
    .Y(_6141_)
);

AND2X2 _16520_ (
    .A(areg_10_bF$buf4),
    .B(breg_18_bF$buf5),
    .Y(_6142_)
);

NOR2X1 _16521_ (
    .A(_6141_),
    .B(_6142_),
    .Y(_6144_)
);

NOR3X1 _16522_ (
    .A(_6138_),
    .B(_6140_),
    .C(_6144_),
    .Y(_6145_)
);

INVX2 _16523_ (
    .A(_6138_),
    .Y(_6146_)
);

NAND2X1 _16524_ (
    .A(_6141_),
    .B(_6142_),
    .Y(_6147_)
);

OAI21X1 _16525_ (
    .A(_7711__bF$buf0),
    .B(_3529__bF$buf1),
    .C(_5768_),
    .Y(_6148_)
);

AOI21X1 _16526_ (
    .A(_6148_),
    .B(_6147_),
    .C(_6146_),
    .Y(_6149_)
);

OAI21X1 _16527_ (
    .A(_6145_),
    .B(_6149_),
    .C(_6137_),
    .Y(_6150_)
);

AOI21X1 _16528_ (
    .A(_5761_),
    .B(_5763_),
    .C(_5769_),
    .Y(_6151_)
);

NAND3X1 _16529_ (
    .A(_6146_),
    .B(_6148_),
    .C(_6147_),
    .Y(_6152_)
);

OAI21X1 _16530_ (
    .A(_6144_),
    .B(_6140_),
    .C(_6138_),
    .Y(_6153_)
);

NAND3X1 _16531_ (
    .A(_6151_),
    .B(_6152_),
    .C(_6153_),
    .Y(_6155_)
);

AOI21X1 _16532_ (
    .A(_6155_),
    .B(_6150_),
    .C(_6136_),
    .Y(_6156_)
);

XNOR2X1 _16533_ (
    .A(_6135_),
    .B(_6131_),
    .Y(_6157_)
);

NAND3X1 _16534_ (
    .A(_6152_),
    .B(_6137_),
    .C(_6153_),
    .Y(_6158_)
);

OAI21X1 _16535_ (
    .A(_6145_),
    .B(_6149_),
    .C(_6151_),
    .Y(_6159_)
);

AOI21X1 _16536_ (
    .A(_6158_),
    .B(_6159_),
    .C(_6157_),
    .Y(_6160_)
);

NOR2X1 _16537_ (
    .A(_6156_),
    .B(_6160_),
    .Y(_6161_)
);

OAI21X1 _16538_ (
    .A(_5808_),
    .B(_5806_),
    .C(_5798_),
    .Y(_6162_)
);

INVX1 _16539_ (
    .A(_5786_),
    .Y(_6163_)
);

OAI21X1 _16540_ (
    .A(_5781_),
    .B(_6163_),
    .C(_5789_),
    .Y(_6164_)
);

NAND2X1 _16541_ (
    .A(areg_11_bF$buf0),
    .B(breg_17_bF$buf2),
    .Y(_6166_)
);

INVX1 _16542_ (
    .A(_6166_),
    .Y(_6167_)
);

AND2X2 _16543_ (
    .A(areg_12_bF$buf1),
    .B(breg_16_bF$buf0),
    .Y(_6168_)
);

AND2X2 _16544_ (
    .A(areg_13_bF$buf4),
    .B(breg_15_bF$buf3),
    .Y(_6169_)
);

NAND2X1 _16545_ (
    .A(_6168_),
    .B(_6169_),
    .Y(_6170_)
);

OAI22X1 _16546_ (
    .A(_10869__bF$buf3),
    .B(_2560__bF$buf0),
    .C(_549__bF$buf2),
    .D(_2362__bF$buf5),
    .Y(_6171_)
);

NAND3X1 _16547_ (
    .A(_6167_),
    .B(_6171_),
    .C(_6170_),
    .Y(_6172_)
);

OAI21X1 _16548_ (
    .A(_10869__bF$buf2),
    .B(_2560__bF$buf4),
    .C(_6169_),
    .Y(_6173_)
);

OAI21X1 _16549_ (
    .A(_549__bF$buf1),
    .B(_2362__bF$buf4),
    .C(_6168_),
    .Y(_6174_)
);

NAND3X1 _16550_ (
    .A(_6166_),
    .B(_6173_),
    .C(_6174_),
    .Y(_6175_)
);

NAND2X1 _16551_ (
    .A(breg_12_bF$buf3),
    .B(areg_15_bF$buf1),
    .Y(_6177_)
);

AND2X2 _16552_ (
    .A(_5468_),
    .B(_6177_),
    .Y(_6178_)
);

OAI22X1 _16553_ (
    .A(_5795_),
    .B(_5842_),
    .C(_6178_),
    .D(_5840_),
    .Y(_6179_)
);

NAND3X1 _16554_ (
    .A(_6172_),
    .B(_6175_),
    .C(_6179_),
    .Y(_6180_)
);

AOI21X1 _16555_ (
    .A(_6173_),
    .B(_6174_),
    .C(_6166_),
    .Y(_6181_)
);

AOI21X1 _16556_ (
    .A(_6171_),
    .B(_6170_),
    .C(_6167_),
    .Y(_6182_)
);

NOR2X1 _16557_ (
    .A(_5468_),
    .B(_6177_),
    .Y(_6183_)
);

AOI21X1 _16558_ (
    .A(_5841_),
    .B(_5843_),
    .C(_6183_),
    .Y(_6184_)
);

OAI21X1 _16559_ (
    .A(_6181_),
    .B(_6182_),
    .C(_6184_),
    .Y(_6185_)
);

NAND3X1 _16560_ (
    .A(_6164_),
    .B(_6180_),
    .C(_6185_),
    .Y(_6186_)
);

AOI21X1 _16561_ (
    .A(_5412_),
    .B(_6168_),
    .C(_5799_),
    .Y(_6188_)
);

NOR3X1 _16562_ (
    .A(_6182_),
    .B(_6184_),
    .C(_6181_),
    .Y(_6189_)
);

AOI21X1 _16563_ (
    .A(_6172_),
    .B(_6175_),
    .C(_6179_),
    .Y(_6190_)
);

OAI21X1 _16564_ (
    .A(_6189_),
    .B(_6190_),
    .C(_6188_),
    .Y(_6191_)
);

NAND3X1 _16565_ (
    .A(_6162_),
    .B(_6186_),
    .C(_6191_),
    .Y(_6192_)
);

AOI21X1 _16566_ (
    .A(_5782_),
    .B(_5803_),
    .C(_5807_),
    .Y(_6193_)
);

NAND3X1 _16567_ (
    .A(_6184_),
    .B(_6172_),
    .C(_6175_),
    .Y(_6194_)
);

OAI21X1 _16568_ (
    .A(_6181_),
    .B(_6182_),
    .C(_6179_),
    .Y(_6195_)
);

AOI21X1 _16569_ (
    .A(_6194_),
    .B(_6195_),
    .C(_6188_),
    .Y(_6196_)
);

AOI21X1 _16570_ (
    .A(_6180_),
    .B(_6185_),
    .C(_6164_),
    .Y(_6197_)
);

OAI21X1 _16571_ (
    .A(_6196_),
    .B(_6197_),
    .C(_6193_),
    .Y(_6199_)
);

NAND3X1 _16572_ (
    .A(_6199_),
    .B(_6161_),
    .C(_6192_),
    .Y(_6200_)
);

OR2X2 _16573_ (
    .A(_6160_),
    .B(_6156_),
    .Y(_6201_)
);

OAI21X1 _16574_ (
    .A(_6196_),
    .B(_6197_),
    .C(_6162_),
    .Y(_6202_)
);

NAND3X1 _16575_ (
    .A(_6193_),
    .B(_6186_),
    .C(_6191_),
    .Y(_6203_)
);

NAND3X1 _16576_ (
    .A(_6202_),
    .B(_6203_),
    .C(_6201_),
    .Y(_6204_)
);

OAI21X1 _16577_ (
    .A(_5873_),
    .B(_5879_),
    .C(_5882_),
    .Y(_6205_)
);

AOI21X1 _16578_ (
    .A(_6200_),
    .B(_6204_),
    .C(_6205_),
    .Y(_6206_)
);

AOI21X1 _16579_ (
    .A(_6202_),
    .B(_6203_),
    .C(_6201_),
    .Y(_6207_)
);

AOI21X1 _16580_ (
    .A(_6199_),
    .B(_6192_),
    .C(_6161_),
    .Y(_6208_)
);

AOI21X1 _16581_ (
    .A(_5839_),
    .B(_5880_),
    .C(_5877_),
    .Y(_6210_)
);

NOR3X1 _16582_ (
    .A(_6210_),
    .B(_6208_),
    .C(_6207_),
    .Y(_6211_)
);

OAI21X1 _16583_ (
    .A(_6211_),
    .B(_6206_),
    .C(_6130_),
    .Y(_6212_)
);

INVX2 _16584_ (
    .A(_6130_),
    .Y(_6213_)
);

OAI21X1 _16585_ (
    .A(_6207_),
    .B(_6208_),
    .C(_6210_),
    .Y(_6214_)
);

NAND3X1 _16586_ (
    .A(_6200_),
    .B(_6205_),
    .C(_6204_),
    .Y(_6215_)
);

NAND3X1 _16587_ (
    .A(_6214_),
    .B(_6215_),
    .C(_6213_),
    .Y(_6216_)
);

NAND2X1 _16588_ (
    .A(_6216_),
    .B(_6212_),
    .Y(_6217_)
);

AOI21X1 _16589_ (
    .A(_5961_),
    .B(_5967_),
    .C(_5886_),
    .Y(_6218_)
);

OAI21X1 _16590_ (
    .A(_5978_),
    .B(_6218_),
    .C(_5968_),
    .Y(_6219_)
);

NAND2X1 _16591_ (
    .A(_5858_),
    .B(_5866_),
    .Y(_6221_)
);

NAND2X1 _16592_ (
    .A(areg_14_bF$buf3),
    .B(breg_14_bF$buf2),
    .Y(_6222_)
);

NAND2X1 _16593_ (
    .A(breg_12_bF$buf2),
    .B(areg_16_bF$buf3),
    .Y(_6223_)
);

XOR2X1 _16594_ (
    .A(_5842_),
    .B(_6223_),
    .Y(_6224_)
);

XNOR2X1 _16595_ (
    .A(_6224_),
    .B(_6222_),
    .Y(_6225_)
);

OAI21X1 _16596_ (
    .A(_5856_),
    .B(_5847_),
    .C(_5851_),
    .Y(_6226_)
);

NAND2X1 _16597_ (
    .A(breg_11_bF$buf4),
    .B(areg_17_bF$buf2),
    .Y(_6227_)
);

INVX2 _16598_ (
    .A(_6227_),
    .Y(_6228_)
);

AND2X2 _16599_ (
    .A(breg_10_bF$buf4),
    .B(areg_19_bF$buf4),
    .Y(_6229_)
);

NAND2X1 _16600_ (
    .A(_5850_),
    .B(_6229_),
    .Y(_6230_)
);

OAI21X1 _16601_ (
    .A(_6044__bF$buf0),
    .B(_3402__bF$buf1),
    .C(_5854_),
    .Y(_6232_)
);

NAND3X1 _16602_ (
    .A(_6228_),
    .B(_6232_),
    .C(_6230_),
    .Y(_6233_)
);

NAND2X1 _16603_ (
    .A(breg_9_bF$buf2),
    .B(areg_19_bF$buf3),
    .Y(_6234_)
);

NOR2X1 _16604_ (
    .A(_5854_),
    .B(_6234_),
    .Y(_6235_)
);

AND2X2 _16605_ (
    .A(_5854_),
    .B(_6234_),
    .Y(_6236_)
);

OAI21X1 _16606_ (
    .A(_6236_),
    .B(_6235_),
    .C(_6227_),
    .Y(_6237_)
);

NAND3X1 _16607_ (
    .A(_6233_),
    .B(_6237_),
    .C(_6226_),
    .Y(_6238_)
);

AOI21X1 _16608_ (
    .A(_5849_),
    .B(_5852_),
    .C(_5855_),
    .Y(_6239_)
);

NOR3X1 _16609_ (
    .A(_6227_),
    .B(_6235_),
    .C(_6236_),
    .Y(_6240_)
);

AOI21X1 _16610_ (
    .A(_6232_),
    .B(_6230_),
    .C(_6228_),
    .Y(_6241_)
);

OAI21X1 _16611_ (
    .A(_6240_),
    .B(_6241_),
    .C(_6239_),
    .Y(_6243_)
);

NAND3X1 _16612_ (
    .A(_6238_),
    .B(_6243_),
    .C(_6225_),
    .Y(_6244_)
);

INVX2 _16613_ (
    .A(_6222_),
    .Y(_6245_)
);

XNOR2X1 _16614_ (
    .A(_6224_),
    .B(_6245_),
    .Y(_6246_)
);

OAI21X1 _16615_ (
    .A(_6240_),
    .B(_6241_),
    .C(_6226_),
    .Y(_6247_)
);

NAND3X1 _16616_ (
    .A(_6239_),
    .B(_6233_),
    .C(_6237_),
    .Y(_6248_)
);

NAND3X1 _16617_ (
    .A(_6247_),
    .B(_6248_),
    .C(_6246_),
    .Y(_6249_)
);

OAI21X1 _16618_ (
    .A(_5908_),
    .B(_5901_),
    .C(_5910_),
    .Y(_6250_)
);

AOI21X1 _16619_ (
    .A(_6244_),
    .B(_6249_),
    .C(_6250_),
    .Y(_6251_)
);

AOI21X1 _16620_ (
    .A(_6247_),
    .B(_6248_),
    .C(_6246_),
    .Y(_6252_)
);

AOI21X1 _16621_ (
    .A(_6238_),
    .B(_6243_),
    .C(_6225_),
    .Y(_6254_)
);

AOI21X1 _16622_ (
    .A(_5888_),
    .B(_5909_),
    .C(_5906_),
    .Y(_6255_)
);

NOR3X1 _16623_ (
    .A(_6254_),
    .B(_6255_),
    .C(_6252_),
    .Y(_6256_)
);

OAI21X1 _16624_ (
    .A(_6256_),
    .B(_6251_),
    .C(_6221_),
    .Y(_6257_)
);

AND2X2 _16625_ (
    .A(_5866_),
    .B(_5858_),
    .Y(_6258_)
);

OAI21X1 _16626_ (
    .A(_6252_),
    .B(_6254_),
    .C(_6255_),
    .Y(_6259_)
);

NAND3X1 _16627_ (
    .A(_6244_),
    .B(_6249_),
    .C(_6250_),
    .Y(_6260_)
);

NAND3X1 _16628_ (
    .A(_6258_),
    .B(_6259_),
    .C(_6260_),
    .Y(_6261_)
);

NAND2X1 _16629_ (
    .A(_6261_),
    .B(_6257_),
    .Y(_6262_)
);

AOI21X1 _16630_ (
    .A(_5953_),
    .B(_5949_),
    .C(_5915_),
    .Y(_6263_)
);

OAI21X1 _16631_ (
    .A(_5964_),
    .B(_6263_),
    .C(_5954_),
    .Y(_6265_)
);

INVX1 _16632_ (
    .A(_5893_),
    .Y(_6266_)
);

OAI21X1 _16633_ (
    .A(_5887_),
    .B(_6266_),
    .C(_5896_),
    .Y(_6267_)
);

NOR2X1 _16634_ (
    .A(_5420__bF$buf1),
    .B(_3958__bF$buf2),
    .Y(_6268_)
);

AND2X2 _16635_ (
    .A(breg_7_bF$buf1),
    .B(areg_21_bF$buf4),
    .Y(_6269_)
);

AND2X2 _16636_ (
    .A(breg_6_bF$buf5),
    .B(areg_22_bF$buf1),
    .Y(_6270_)
);

NAND2X1 _16637_ (
    .A(_6269_),
    .B(_6270_),
    .Y(_6271_)
);

OAI22X1 _16638_ (
    .A(_5453__bF$buf1),
    .B(_4551__bF$buf2),
    .C(_4116__bF$buf3),
    .D(_3961__bF$buf0),
    .Y(_6272_)
);

NAND3X1 _16639_ (
    .A(_6268_),
    .B(_6272_),
    .C(_6271_),
    .Y(_6273_)
);

INVX1 _16640_ (
    .A(_6268_),
    .Y(_6274_)
);

OAI21X1 _16641_ (
    .A(_4116__bF$buf2),
    .B(_3961__bF$buf4),
    .C(_6270_),
    .Y(_6276_)
);

OAI21X1 _16642_ (
    .A(_5453__bF$buf0),
    .B(_4551__bF$buf1),
    .C(_6269_),
    .Y(_6277_)
);

NAND3X1 _16643_ (
    .A(_6276_),
    .B(_6277_),
    .C(_6274_),
    .Y(_6278_)
);

AOI21X1 _16644_ (
    .A(_5917_),
    .B(_5922_),
    .C(_5924_),
    .Y(_6279_)
);

INVX1 _16645_ (
    .A(_6279_),
    .Y(_6280_)
);

AOI21X1 _16646_ (
    .A(_6273_),
    .B(_6278_),
    .C(_6280_),
    .Y(_6281_)
);

AOI21X1 _16647_ (
    .A(_6276_),
    .B(_6277_),
    .C(_6274_),
    .Y(_6282_)
);

AOI21X1 _16648_ (
    .A(_6272_),
    .B(_6271_),
    .C(_6268_),
    .Y(_6283_)
);

NOR3X1 _16649_ (
    .A(_6283_),
    .B(_6279_),
    .C(_6282_),
    .Y(_6284_)
);

OAI21X1 _16650_ (
    .A(_6281_),
    .B(_6284_),
    .C(_6267_),
    .Y(_6285_)
);

INVX2 _16651_ (
    .A(_6267_),
    .Y(_6287_)
);

OAI21X1 _16652_ (
    .A(_6282_),
    .B(_6283_),
    .C(_6279_),
    .Y(_6288_)
);

NAND3X1 _16653_ (
    .A(_6273_),
    .B(_6278_),
    .C(_6280_),
    .Y(_6289_)
);

NAND3X1 _16654_ (
    .A(_6288_),
    .B(_6287_),
    .C(_6289_),
    .Y(_6290_)
);

NAND2X1 _16655_ (
    .A(_6290_),
    .B(_6285_),
    .Y(_6291_)
);

AOI21X1 _16656_ (
    .A(_5940_),
    .B(_5937_),
    .C(_5929_),
    .Y(_6292_)
);

OAI21X1 _16657_ (
    .A(_6292_),
    .B(_5950_),
    .C(_5941_),
    .Y(_6293_)
);

NAND2X1 _16658_ (
    .A(breg_5_bF$buf1),
    .B(areg_23_bF$buf2),
    .Y(_6294_)
);

INVX1 _16659_ (
    .A(_6294_),
    .Y(_6295_)
);

NAND2X1 _16660_ (
    .A(breg_4_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_6296_)
);

NAND2X1 _16661_ (
    .A(breg_3_bF$buf0),
    .B(areg_25_bF$buf4),
    .Y(_6298_)
);

OR2X2 _16662_ (
    .A(_6296_),
    .B(_6298_),
    .Y(_6299_)
);

INVX8 _16663_ (
    .A(areg_25_bF$buf3),
    .Y(_6300_)
);

OAI21X1 _16664_ (
    .A(_2365_),
    .B(_6300__bF$buf3),
    .C(_6296_),
    .Y(_6301_)
);

NAND3X1 _16665_ (
    .A(_6295_),
    .B(_6301_),
    .C(_6299_),
    .Y(_6302_)
);

NOR2X1 _16666_ (
    .A(_6296_),
    .B(_6298_),
    .Y(_6303_)
);

AND2X2 _16667_ (
    .A(_6296_),
    .B(_6298_),
    .Y(_6304_)
);

OAI21X1 _16668_ (
    .A(_6304_),
    .B(_6303_),
    .C(_6294_),
    .Y(_6305_)
);

AND2X2 _16669_ (
    .A(_6302_),
    .B(_6305_),
    .Y(_6306_)
);

OAI21X1 _16670_ (
    .A(_5930_),
    .B(_5934_),
    .C(_5933_),
    .Y(_6307_)
);

NAND2X1 _16671_ (
    .A(breg_2_bF$buf0),
    .B(areg_26_bF$buf0),
    .Y(_6309_)
);

INVX2 _16672_ (
    .A(_6309_),
    .Y(_6310_)
);

AND2X2 _16673_ (
    .A(breg_1_bF$buf5),
    .B(areg_27_bF$buf2),
    .Y(_6311_)
);

AND2X2 _16674_ (
    .A(breg_0_bF$buf4),
    .B(areg_28_bF$buf5),
    .Y(_6312_)
);

NAND2X1 _16675_ (
    .A(_6311_),
    .B(_6312_),
    .Y(_6313_)
);

AOI22X1 _16676_ (
    .A(breg_0_bF$buf3),
    .B(areg_28_bF$buf4),
    .C(breg_1_bF$buf4),
    .D(areg_27_bF$buf1),
    .Y(_6314_)
);

INVX2 _16677_ (
    .A(_6314_),
    .Y(_6315_)
);

NAND3X1 _16678_ (
    .A(_6310_),
    .B(_6315_),
    .C(_6313_),
    .Y(_6316_)
);

NAND2X1 _16679_ (
    .A(breg_1_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_6317_)
);

NAND2X1 _16680_ (
    .A(breg_0_bF$buf2),
    .B(areg_28_bF$buf3),
    .Y(_6318_)
);

NOR2X1 _16681_ (
    .A(_6317_),
    .B(_6318_),
    .Y(_6320_)
);

OAI21X1 _16682_ (
    .A(_6320_),
    .B(_6314_),
    .C(_6309_),
    .Y(_6321_)
);

NAND3X1 _16683_ (
    .A(_6307_),
    .B(_6321_),
    .C(_6316_),
    .Y(_6322_)
);

AOI21X1 _16684_ (
    .A(_5931_),
    .B(_5935_),
    .C(_5939_),
    .Y(_6323_)
);

NAND2X1 _16685_ (
    .A(_6317_),
    .B(_6312_),
    .Y(_6324_)
);

NAND2X1 _16686_ (
    .A(_6318_),
    .B(_6311_),
    .Y(_6325_)
);

AOI21X1 _16687_ (
    .A(_6324_),
    .B(_6325_),
    .C(_6309_),
    .Y(_6326_)
);

AOI21X1 _16688_ (
    .A(_6315_),
    .B(_6313_),
    .C(_6310_),
    .Y(_6327_)
);

OAI21X1 _16689_ (
    .A(_6327_),
    .B(_6326_),
    .C(_6323_),
    .Y(_6328_)
);

NAND3X1 _16690_ (
    .A(_6322_),
    .B(_6328_),
    .C(_6306_),
    .Y(_6329_)
);

NAND2X1 _16691_ (
    .A(_6305_),
    .B(_6302_),
    .Y(_6331_)
);

OAI21X1 _16692_ (
    .A(_6327_),
    .B(_6326_),
    .C(_6307_),
    .Y(_6332_)
);

NAND3X1 _16693_ (
    .A(_6321_),
    .B(_6323_),
    .C(_6316_),
    .Y(_6333_)
);

NAND3X1 _16694_ (
    .A(_6331_),
    .B(_6333_),
    .C(_6332_),
    .Y(_6334_)
);

NAND3X1 _16695_ (
    .A(_6293_),
    .B(_6334_),
    .C(_6329_),
    .Y(_6335_)
);

NOR3X1 _16696_ (
    .A(_5945_),
    .B(_5942_),
    .C(_5946_),
    .Y(_6336_)
);

AOI21X1 _16697_ (
    .A(_5928_),
    .B(_5948_),
    .C(_6336_),
    .Y(_6337_)
);

AOI21X1 _16698_ (
    .A(_6333_),
    .B(_6332_),
    .C(_6331_),
    .Y(_6338_)
);

AOI21X1 _16699_ (
    .A(_6322_),
    .B(_6328_),
    .C(_6306_),
    .Y(_6339_)
);

OAI21X1 _16700_ (
    .A(_6338_),
    .B(_6339_),
    .C(_6337_),
    .Y(_6340_)
);

NAND3X1 _16701_ (
    .A(_6335_),
    .B(_6340_),
    .C(_6291_),
    .Y(_6342_)
);

NAND3X1 _16702_ (
    .A(_6267_),
    .B(_6288_),
    .C(_6289_),
    .Y(_6343_)
);

OAI21X1 _16703_ (
    .A(_6281_),
    .B(_6284_),
    .C(_6287_),
    .Y(_6344_)
);

NAND2X1 _16704_ (
    .A(_6343_),
    .B(_6344_),
    .Y(_6345_)
);

OAI21X1 _16705_ (
    .A(_6338_),
    .B(_6339_),
    .C(_6293_),
    .Y(_6346_)
);

NAND3X1 _16706_ (
    .A(_6329_),
    .B(_6334_),
    .C(_6337_),
    .Y(_6347_)
);

NAND3X1 _16707_ (
    .A(_6347_),
    .B(_6346_),
    .C(_6345_),
    .Y(_6348_)
);

NAND3X1 _16708_ (
    .A(_6265_),
    .B(_6342_),
    .C(_6348_),
    .Y(_6349_)
);

NOR3X1 _16709_ (
    .A(_5957_),
    .B(_5959_),
    .C(_5956_),
    .Y(_6350_)
);

AOI21X1 _16710_ (
    .A(_5912_),
    .B(_5960_),
    .C(_6350_),
    .Y(_6351_)
);

AOI21X1 _16711_ (
    .A(_6347_),
    .B(_6346_),
    .C(_6345_),
    .Y(_6353_)
);

AOI21X1 _16712_ (
    .A(_6335_),
    .B(_6340_),
    .C(_6291_),
    .Y(_6354_)
);

OAI21X1 _16713_ (
    .A(_6353_),
    .B(_6354_),
    .C(_6351_),
    .Y(_6355_)
);

NAND3X1 _16714_ (
    .A(_6349_),
    .B(_6355_),
    .C(_6262_),
    .Y(_6356_)
);

NAND3X1 _16715_ (
    .A(_6221_),
    .B(_6259_),
    .C(_6260_),
    .Y(_6357_)
);

OAI21X1 _16716_ (
    .A(_6256_),
    .B(_6251_),
    .C(_6258_),
    .Y(_6358_)
);

NAND2X1 _16717_ (
    .A(_6357_),
    .B(_6358_),
    .Y(_6359_)
);

OAI21X1 _16718_ (
    .A(_6353_),
    .B(_6354_),
    .C(_6265_),
    .Y(_6360_)
);

NAND3X1 _16719_ (
    .A(_6342_),
    .B(_6348_),
    .C(_6351_),
    .Y(_6361_)
);

NAND3X1 _16720_ (
    .A(_6361_),
    .B(_6360_),
    .C(_6359_),
    .Y(_6362_)
);

NAND3X1 _16721_ (
    .A(_6356_),
    .B(_6219_),
    .C(_6362_),
    .Y(_6364_)
);

NOR3X1 _16722_ (
    .A(_5972_),
    .B(_5973_),
    .C(_5971_),
    .Y(_6365_)
);

AOI21X1 _16723_ (
    .A(_5884_),
    .B(_5974_),
    .C(_6365_),
    .Y(_6366_)
);

AOI21X1 _16724_ (
    .A(_6361_),
    .B(_6360_),
    .C(_6359_),
    .Y(_6367_)
);

AOI21X1 _16725_ (
    .A(_6349_),
    .B(_6355_),
    .C(_6262_),
    .Y(_6368_)
);

OAI21X1 _16726_ (
    .A(_6367_),
    .B(_6368_),
    .C(_6366_),
    .Y(_6369_)
);

NAND3X1 _16727_ (
    .A(_6364_),
    .B(_6369_),
    .C(_6217_),
    .Y(_6370_)
);

NAND3X1 _16728_ (
    .A(_6130_),
    .B(_6215_),
    .C(_6214_),
    .Y(_6371_)
);

OAI21X1 _16729_ (
    .A(_6211_),
    .B(_6206_),
    .C(_6213_),
    .Y(_6372_)
);

NAND2X1 _16730_ (
    .A(_6371_),
    .B(_6372_),
    .Y(_6373_)
);

OAI21X1 _16731_ (
    .A(_6367_),
    .B(_6368_),
    .C(_6219_),
    .Y(_6375_)
);

NAND3X1 _16732_ (
    .A(_6356_),
    .B(_6362_),
    .C(_6366_),
    .Y(_6376_)
);

NAND3X1 _16733_ (
    .A(_6375_),
    .B(_6376_),
    .C(_6373_),
    .Y(_6377_)
);

NAND3X1 _16734_ (
    .A(_6370_),
    .B(_6377_),
    .C(_6129_),
    .Y(_6378_)
);

NOR3X1 _16735_ (
    .A(_5985_),
    .B(_5986_),
    .C(_5984_),
    .Y(_6379_)
);

AOI21X1 _16736_ (
    .A(_5835_),
    .B(_5987_),
    .C(_6379_),
    .Y(_6380_)
);

AOI21X1 _16737_ (
    .A(_6376_),
    .B(_6375_),
    .C(_6373_),
    .Y(_6381_)
);

AOI21X1 _16738_ (
    .A(_6364_),
    .B(_6369_),
    .C(_6217_),
    .Y(_6382_)
);

OAI21X1 _16739_ (
    .A(_6381_),
    .B(_6382_),
    .C(_6380_),
    .Y(_6383_)
);

NAND3X1 _16740_ (
    .A(_6378_),
    .B(_6383_),
    .C(_6127_),
    .Y(_6384_)
);

NAND3X1 _16741_ (
    .A(_6123_),
    .B(_6124_),
    .C(_6125_),
    .Y(_6386_)
);

NAND3X1 _16742_ (
    .A(_6116_),
    .B(_6048_),
    .C(_6120_),
    .Y(_6387_)
);

NAND2X1 _16743_ (
    .A(_6386_),
    .B(_6387_),
    .Y(_6388_)
);

OAI21X1 _16744_ (
    .A(_6381_),
    .B(_6382_),
    .C(_6129_),
    .Y(_6389_)
);

NAND3X1 _16745_ (
    .A(_6370_),
    .B(_6377_),
    .C(_6380_),
    .Y(_6390_)
);

NAND3X1 _16746_ (
    .A(_6388_),
    .B(_6390_),
    .C(_6389_),
    .Y(_6391_)
);

NAND3X1 _16747_ (
    .A(_6391_),
    .B(_6047_),
    .C(_6384_),
    .Y(_6392_)
);

NOR3X1 _16748_ (
    .A(_5999_),
    .B(_6000_),
    .C(_5998_),
    .Y(_6393_)
);

AOI21X1 _16749_ (
    .A(_5743_),
    .B(_6002_),
    .C(_6393_),
    .Y(_6394_)
);

AOI21X1 _16750_ (
    .A(_6390_),
    .B(_6389_),
    .C(_6388_),
    .Y(_6395_)
);

AOI21X1 _16751_ (
    .A(_6378_),
    .B(_6383_),
    .C(_6127_),
    .Y(_6397_)
);

OAI21X1 _16752_ (
    .A(_6397_),
    .B(_6395_),
    .C(_6394_),
    .Y(_6398_)
);

NAND3X1 _16753_ (
    .A(_6045_),
    .B(_6392_),
    .C(_6398_),
    .Y(_6399_)
);

INVX2 _16754_ (
    .A(_6045_),
    .Y(_6400_)
);

NOR3X1 _16755_ (
    .A(_6397_),
    .B(_6395_),
    .C(_6394_),
    .Y(_6401_)
);

AOI21X1 _16756_ (
    .A(_6391_),
    .B(_6384_),
    .C(_6047_),
    .Y(_6402_)
);

OAI21X1 _16757_ (
    .A(_6401_),
    .B(_6402_),
    .C(_6400_),
    .Y(_6403_)
);

NAND3X1 _16758_ (
    .A(_6043_),
    .B(_6399_),
    .C(_6403_),
    .Y(_6404_)
);

AOI21X1 _16759_ (
    .A(_5666_),
    .B(_6015_),
    .C(_6018_),
    .Y(_6405_)
);

OAI21X1 _16760_ (
    .A(_6397_),
    .B(_6395_),
    .C(_6047_),
    .Y(_6406_)
);

NAND3X1 _16761_ (
    .A(_6391_),
    .B(_6384_),
    .C(_6394_),
    .Y(_6408_)
);

AOI21X1 _16762_ (
    .A(_6408_),
    .B(_6406_),
    .C(_6400_),
    .Y(_6409_)
);

AOI21X1 _16763_ (
    .A(_6392_),
    .B(_6398_),
    .C(_6045_),
    .Y(_6410_)
);

OAI21X1 _16764_ (
    .A(_6409_),
    .B(_6410_),
    .C(_6405_),
    .Y(_6411_)
);

NAND3X1 _16765_ (
    .A(_6404_),
    .B(_6411_),
    .C(_6030_),
    .Y(_6412_)
);

OAI21X1 _16766_ (
    .A(_6409_),
    .B(_6410_),
    .C(_6043_),
    .Y(_6413_)
);

NAND3X1 _16767_ (
    .A(_6405_),
    .B(_6399_),
    .C(_6403_),
    .Y(_6414_)
);

NAND3X1 _16768_ (
    .A(_6413_),
    .B(_6021_),
    .C(_6414_),
    .Y(_6415_)
);

NAND2X1 _16769_ (
    .A(_6415_),
    .B(_6412_),
    .Y(_6416_)
);

XOR2X1 _16770_ (
    .A(_6042_),
    .B(_6416_),
    .Y(_0_[28])
);

OAI21X1 _16771_ (
    .A(_6042_),
    .B(_6416_),
    .C(_6412_),
    .Y(_6418_)
);

NOR3X1 _16772_ (
    .A(_6409_),
    .B(_6410_),
    .C(_6405_),
    .Y(_6419_)
);

OAI21X1 _16773_ (
    .A(_6402_),
    .B(_6400_),
    .C(_6392_),
    .Y(_6420_)
);

NAND2X1 _16774_ (
    .A(_6124_),
    .B(_6386_),
    .Y(_6421_)
);

AOI21X1 _16775_ (
    .A(_6370_),
    .B(_6377_),
    .C(_6129_),
    .Y(_6422_)
);

OAI21X1 _16776_ (
    .A(_6422_),
    .B(_6388_),
    .C(_6378_),
    .Y(_6423_)
);

NAND2X1 _16777_ (
    .A(_6102_),
    .B(_6111_),
    .Y(_6424_)
);

INVX1 _16778_ (
    .A(_6049_),
    .Y(_6425_)
);

NAND2X1 _16779_ (
    .A(_6425_),
    .B(_5669_),
    .Y(_6426_)
);

INVX4 _16780_ (
    .A(breg_29_bF$buf4),
    .Y(_6427_)
);

NOR2X1 _16781_ (
    .A(_2376__bF$buf3),
    .B(_6427_),
    .Y(_6429_)
);

NAND2X1 _16782_ (
    .A(areg_2_bF$buf0),
    .B(breg_28_bF$buf3),
    .Y(_6430_)
);

OAI21X1 _16783_ (
    .A(_2519__bF$buf2),
    .B(_5668__bF$buf4),
    .C(_6049_),
    .Y(_6431_)
);

OAI21X1 _16784_ (
    .A(_6051_),
    .B(_6430_),
    .C(_6431_),
    .Y(_6432_)
);

XNOR2X1 _16785_ (
    .A(_6432_),
    .B(_6429_),
    .Y(_6433_)
);

INVX1 _16786_ (
    .A(_6433_),
    .Y(_6434_)
);

NOR2X1 _16787_ (
    .A(_6426_),
    .B(_6434_),
    .Y(_6435_)
);

INVX1 _16788_ (
    .A(_6435_),
    .Y(_6436_)
);

OAI21X1 _16789_ (
    .A(_5726_),
    .B(_6049_),
    .C(_6434_),
    .Y(_6437_)
);

NAND2X1 _16790_ (
    .A(_6437_),
    .B(_6436_),
    .Y(_6438_)
);

OAI21X1 _16791_ (
    .A(_6097_),
    .B(_6100_),
    .C(_6090_),
    .Y(_6440_)
);

AND2X2 _16792_ (
    .A(_6081_),
    .B(_6073_),
    .Y(_6441_)
);

INVX1 _16793_ (
    .A(_6063_),
    .Y(_6442_)
);

OAI21X1 _16794_ (
    .A(_5685_),
    .B(_6442_),
    .C(_6066_),
    .Y(_6443_)
);

NAND2X1 _16795_ (
    .A(areg_3_bF$buf0),
    .B(breg_26_bF$buf1),
    .Y(_6444_)
);

INVX1 _16796_ (
    .A(_6444_),
    .Y(_6445_)
);

AND2X2 _16797_ (
    .A(areg_4_bF$buf4),
    .B(breg_25_bF$buf3),
    .Y(_6446_)
);

AND2X2 _16798_ (
    .A(areg_5_bF$buf3),
    .B(breg_24_bF$buf4),
    .Y(_6447_)
);

NAND2X1 _16799_ (
    .A(_6446_),
    .B(_6447_),
    .Y(_6448_)
);

OAI22X1 _16800_ (
    .A(_2825__bF$buf3),
    .B(_5315__bF$buf3),
    .C(_2562__bF$buf0),
    .D(_5318_),
    .Y(_6449_)
);

NAND3X1 _16801_ (
    .A(_6445_),
    .B(_6449_),
    .C(_6448_),
    .Y(_6451_)
);

OAI21X1 _16802_ (
    .A(_2562__bF$buf4),
    .B(_5318_),
    .C(_6447_),
    .Y(_6452_)
);

OAI21X1 _16803_ (
    .A(_2825__bF$buf2),
    .B(_5315__bF$buf2),
    .C(_6446_),
    .Y(_6453_)
);

NAND3X1 _16804_ (
    .A(_6444_),
    .B(_6452_),
    .C(_6453_),
    .Y(_6454_)
);

NAND2X1 _16805_ (
    .A(areg_7_bF$buf4),
    .B(breg_22_bF$buf2),
    .Y(_6455_)
);

AND2X2 _16806_ (
    .A(_6070_),
    .B(_6134_),
    .Y(_6456_)
);

OAI22X1 _16807_ (
    .A(_5750_),
    .B(_6455_),
    .C(_6456_),
    .D(_6131_),
    .Y(_6457_)
);

NAND3X1 _16808_ (
    .A(_6451_),
    .B(_6454_),
    .C(_6457_),
    .Y(_6458_)
);

AOI21X1 _16809_ (
    .A(_6452_),
    .B(_6453_),
    .C(_6444_),
    .Y(_6459_)
);

AOI21X1 _16810_ (
    .A(_6449_),
    .B(_6448_),
    .C(_6445_),
    .Y(_6460_)
);

NOR2X1 _16811_ (
    .A(_6070_),
    .B(_6134_),
    .Y(_6462_)
);

OAI21X1 _16812_ (
    .A(_4434__bF$buf3),
    .B(_3781__bF$buf2),
    .C(_6070_),
    .Y(_6463_)
);

AOI21X1 _16813_ (
    .A(_6133_),
    .B(_6463_),
    .C(_6462_),
    .Y(_6464_)
);

OAI21X1 _16814_ (
    .A(_6459_),
    .B(_6460_),
    .C(_6464_),
    .Y(_6465_)
);

NAND3X1 _16815_ (
    .A(_6443_),
    .B(_6458_),
    .C(_6465_),
    .Y(_6466_)
);

AOI21X1 _16816_ (
    .A(_5679_),
    .B(_6446_),
    .C(_6074_),
    .Y(_6467_)
);

NAND3X1 _16817_ (
    .A(_6464_),
    .B(_6451_),
    .C(_6454_),
    .Y(_6468_)
);

OAI21X1 _16818_ (
    .A(_6459_),
    .B(_6460_),
    .C(_6457_),
    .Y(_6469_)
);

NAND3X1 _16819_ (
    .A(_6467_),
    .B(_6468_),
    .C(_6469_),
    .Y(_6470_)
);

NOR3X1 _16820_ (
    .A(_6149_),
    .B(_6151_),
    .C(_6145_),
    .Y(_6471_)
);

AOI21X1 _16821_ (
    .A(_6159_),
    .B(_6157_),
    .C(_6471_),
    .Y(_6473_)
);

NAND3X1 _16822_ (
    .A(_6466_),
    .B(_6470_),
    .C(_6473_),
    .Y(_6474_)
);

AOI21X1 _16823_ (
    .A(_6468_),
    .B(_6469_),
    .C(_6467_),
    .Y(_6475_)
);

AOI21X1 _16824_ (
    .A(_6458_),
    .B(_6465_),
    .C(_6443_),
    .Y(_6476_)
);

AOI21X1 _16825_ (
    .A(_6152_),
    .B(_6153_),
    .C(_6137_),
    .Y(_6477_)
);

OAI21X1 _16826_ (
    .A(_6136_),
    .B(_6477_),
    .C(_6158_),
    .Y(_6478_)
);

OAI21X1 _16827_ (
    .A(_6475_),
    .B(_6476_),
    .C(_6478_),
    .Y(_6479_)
);

AOI21X1 _16828_ (
    .A(_6479_),
    .B(_6474_),
    .C(_6441_),
    .Y(_6480_)
);

NAND2X1 _16829_ (
    .A(_6073_),
    .B(_6081_),
    .Y(_6481_)
);

NAND3X1 _16830_ (
    .A(_6466_),
    .B(_6470_),
    .C(_6478_),
    .Y(_6482_)
);

OAI21X1 _16831_ (
    .A(_6475_),
    .B(_6476_),
    .C(_6473_),
    .Y(_6484_)
);

AOI21X1 _16832_ (
    .A(_6484_),
    .B(_6482_),
    .C(_6481_),
    .Y(_6485_)
);

OAI21X1 _16833_ (
    .A(_6480_),
    .B(_6485_),
    .C(_6440_),
    .Y(_6486_)
);

AOI21X1 _16834_ (
    .A(_6058_),
    .B(_6095_),
    .C(_6098_),
    .Y(_6487_)
);

NAND3X1 _16835_ (
    .A(_6481_),
    .B(_6484_),
    .C(_6482_),
    .Y(_6488_)
);

NAND3X1 _16836_ (
    .A(_6441_),
    .B(_6479_),
    .C(_6474_),
    .Y(_6489_)
);

NAND3X1 _16837_ (
    .A(_6488_),
    .B(_6489_),
    .C(_6487_),
    .Y(_6490_)
);

AOI21X1 _16838_ (
    .A(_6490_),
    .B(_6486_),
    .C(_6438_),
    .Y(_6491_)
);

INVX1 _16839_ (
    .A(_6438_),
    .Y(_6492_)
);

NAND3X1 _16840_ (
    .A(_6488_),
    .B(_6489_),
    .C(_6440_),
    .Y(_6493_)
);

OAI21X1 _16841_ (
    .A(_6480_),
    .B(_6485_),
    .C(_6487_),
    .Y(_6495_)
);

AOI21X1 _16842_ (
    .A(_6493_),
    .B(_6495_),
    .C(_6492_),
    .Y(_6496_)
);

AOI21X1 _16843_ (
    .A(_6130_),
    .B(_6214_),
    .C(_6211_),
    .Y(_6497_)
);

NOR3X1 _16844_ (
    .A(_6491_),
    .B(_6496_),
    .C(_6497_),
    .Y(_6498_)
);

NAND3X1 _16845_ (
    .A(_6492_),
    .B(_6493_),
    .C(_6495_),
    .Y(_6499_)
);

NAND3X1 _16846_ (
    .A(_6438_),
    .B(_6490_),
    .C(_6486_),
    .Y(_6500_)
);

OAI21X1 _16847_ (
    .A(_6213_),
    .B(_6206_),
    .C(_6215_),
    .Y(_6501_)
);

AOI21X1 _16848_ (
    .A(_6499_),
    .B(_6500_),
    .C(_6501_),
    .Y(_6502_)
);

OAI21X1 _16849_ (
    .A(_6498_),
    .B(_6502_),
    .C(_6424_),
    .Y(_6503_)
);

AND2X2 _16850_ (
    .A(_6111_),
    .B(_6102_),
    .Y(_6504_)
);

NAND3X1 _16851_ (
    .A(_6499_),
    .B(_6500_),
    .C(_6501_),
    .Y(_6506_)
);

OAI21X1 _16852_ (
    .A(_6491_),
    .B(_6496_),
    .C(_6497_),
    .Y(_6507_)
);

NAND3X1 _16853_ (
    .A(_6504_),
    .B(_6507_),
    .C(_6506_),
    .Y(_6508_)
);

NAND2X1 _16854_ (
    .A(_6508_),
    .B(_6503_),
    .Y(_6509_)
);

AOI21X1 _16855_ (
    .A(_6356_),
    .B(_6362_),
    .C(_6219_),
    .Y(_6510_)
);

OAI21X1 _16856_ (
    .A(_6373_),
    .B(_6510_),
    .C(_6364_),
    .Y(_6511_)
);

NAND2X1 _16857_ (
    .A(_6192_),
    .B(_6200_),
    .Y(_6512_)
);

NOR2X1 _16858_ (
    .A(_3646__bF$buf1),
    .B(_5369_),
    .Y(_6513_)
);

NAND2X1 _16859_ (
    .A(areg_8_bF$buf3),
    .B(breg_21_bF$buf2),
    .Y(_6514_)
);

XOR2X1 _16860_ (
    .A(_6455_),
    .B(_6514_),
    .Y(_6515_)
);

XNOR2X1 _16861_ (
    .A(_6515_),
    .B(_6513_),
    .Y(_6517_)
);

OAI21X1 _16862_ (
    .A(_6144_),
    .B(_6138_),
    .C(_6147_),
    .Y(_6518_)
);

NOR2X1 _16863_ (
    .A(_6582__bF$buf3),
    .B(_3526_),
    .Y(_6519_)
);

INVX2 _16864_ (
    .A(_6519_),
    .Y(_6520_)
);

AND2X2 _16865_ (
    .A(areg_11_bF$buf4),
    .B(breg_18_bF$buf4),
    .Y(_6521_)
);

OAI21X1 _16866_ (
    .A(_7711__bF$buf3),
    .B(_3253__bF$buf3),
    .C(_6521_),
    .Y(_6522_)
);

AND2X2 _16867_ (
    .A(areg_10_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_6523_)
);

OAI21X1 _16868_ (
    .A(_9104__bF$buf1),
    .B(_3529__bF$buf0),
    .C(_6523_),
    .Y(_6524_)
);

AOI21X1 _16869_ (
    .A(_6522_),
    .B(_6524_),
    .C(_6520_),
    .Y(_6525_)
);

NAND2X1 _16870_ (
    .A(_6523_),
    .B(_6521_),
    .Y(_6526_)
);

OAI22X1 _16871_ (
    .A(_7711__bF$buf2),
    .B(_3253__bF$buf2),
    .C(_9104__bF$buf0),
    .D(_3529__bF$buf4),
    .Y(_6528_)
);

AOI21X1 _16872_ (
    .A(_6528_),
    .B(_6526_),
    .C(_6519_),
    .Y(_6529_)
);

OAI21X1 _16873_ (
    .A(_6525_),
    .B(_6529_),
    .C(_6518_),
    .Y(_6530_)
);

AOI21X1 _16874_ (
    .A(_6146_),
    .B(_6148_),
    .C(_6140_),
    .Y(_6531_)
);

NAND3X1 _16875_ (
    .A(_6519_),
    .B(_6528_),
    .C(_6526_),
    .Y(_6532_)
);

NAND2X1 _16876_ (
    .A(areg_11_bF$buf3),
    .B(breg_19_bF$buf4),
    .Y(_6533_)
);

NOR2X1 _16877_ (
    .A(_6139_),
    .B(_6533_),
    .Y(_6534_)
);

NOR2X1 _16878_ (
    .A(_6523_),
    .B(_6521_),
    .Y(_6535_)
);

OAI21X1 _16879_ (
    .A(_6535_),
    .B(_6534_),
    .C(_6520_),
    .Y(_6536_)
);

NAND3X1 _16880_ (
    .A(_6531_),
    .B(_6532_),
    .C(_6536_),
    .Y(_6537_)
);

AOI21X1 _16881_ (
    .A(_6537_),
    .B(_6530_),
    .C(_6517_),
    .Y(_6539_)
);

INVX2 _16882_ (
    .A(_6513_),
    .Y(_6540_)
);

XNOR2X1 _16883_ (
    .A(_6515_),
    .B(_6540_),
    .Y(_6541_)
);

NAND3X1 _16884_ (
    .A(_6532_),
    .B(_6518_),
    .C(_6536_),
    .Y(_6542_)
);

OAI21X1 _16885_ (
    .A(_6525_),
    .B(_6529_),
    .C(_6531_),
    .Y(_6543_)
);

AOI21X1 _16886_ (
    .A(_6542_),
    .B(_6543_),
    .C(_6541_),
    .Y(_6544_)
);

NOR2X1 _16887_ (
    .A(_6544_),
    .B(_6539_),
    .Y(_6545_)
);

OAI21X1 _16888_ (
    .A(_6190_),
    .B(_6188_),
    .C(_6180_),
    .Y(_6546_)
);

NAND2X1 _16889_ (
    .A(areg_13_bF$buf3),
    .B(breg_16_bF$buf5),
    .Y(_6547_)
);

OAI21X1 _16890_ (
    .A(_6163_),
    .B(_6547_),
    .C(_6172_),
    .Y(_6548_)
);

NAND2X1 _16891_ (
    .A(areg_12_bF$buf0),
    .B(breg_17_bF$buf1),
    .Y(_6550_)
);

INVX1 _16892_ (
    .A(_6550_),
    .Y(_6551_)
);

AND2X2 _16893_ (
    .A(areg_13_bF$buf2),
    .B(breg_16_bF$buf4),
    .Y(_6552_)
);

AND2X2 _16894_ (
    .A(areg_14_bF$buf2),
    .B(breg_15_bF$buf2),
    .Y(_6553_)
);

NAND2X1 _16895_ (
    .A(_6552_),
    .B(_6553_),
    .Y(_6554_)
);

OAI21X1 _16896_ (
    .A(_2287__bF$buf1),
    .B(_2362__bF$buf3),
    .C(_6547_),
    .Y(_6555_)
);

NAND3X1 _16897_ (
    .A(_6551_),
    .B(_6555_),
    .C(_6554_),
    .Y(_6556_)
);

OAI21X1 _16898_ (
    .A(_549__bF$buf0),
    .B(_2560__bF$buf3),
    .C(_6553_),
    .Y(_6557_)
);

OAI21X1 _16899_ (
    .A(_2287__bF$buf0),
    .B(_2362__bF$buf2),
    .C(_6552_),
    .Y(_6558_)
);

NAND3X1 _16900_ (
    .A(_6550_),
    .B(_6557_),
    .C(_6558_),
    .Y(_6559_)
);

NAND2X1 _16901_ (
    .A(breg_13_bF$buf3),
    .B(areg_16_bF$buf2),
    .Y(_6561_)
);

AND2X2 _16902_ (
    .A(_5842_),
    .B(_6223_),
    .Y(_6562_)
);

OAI22X1 _16903_ (
    .A(_6177_),
    .B(_6561_),
    .C(_6562_),
    .D(_6222_),
    .Y(_6563_)
);

NAND3X1 _16904_ (
    .A(_6556_),
    .B(_6559_),
    .C(_6563_),
    .Y(_6564_)
);

AOI21X1 _16905_ (
    .A(_6557_),
    .B(_6558_),
    .C(_6550_),
    .Y(_6565_)
);

AOI21X1 _16906_ (
    .A(_6555_),
    .B(_6554_),
    .C(_6551_),
    .Y(_6566_)
);

NOR2X1 _16907_ (
    .A(_5842_),
    .B(_6223_),
    .Y(_6567_)
);

OAI21X1 _16908_ (
    .A(_2586__bF$buf2),
    .B(_2669__bF$buf3),
    .C(_5842_),
    .Y(_6568_)
);

AOI21X1 _16909_ (
    .A(_6245_),
    .B(_6568_),
    .C(_6567_),
    .Y(_6569_)
);

OAI21X1 _16910_ (
    .A(_6565_),
    .B(_6566_),
    .C(_6569_),
    .Y(_6570_)
);

NAND3X1 _16911_ (
    .A(_6548_),
    .B(_6564_),
    .C(_6570_),
    .Y(_6572_)
);

AOI21X1 _16912_ (
    .A(_5786_),
    .B(_6552_),
    .C(_6181_),
    .Y(_6573_)
);

NAND3X1 _16913_ (
    .A(_6569_),
    .B(_6556_),
    .C(_6559_),
    .Y(_6574_)
);

OAI21X1 _16914_ (
    .A(_6565_),
    .B(_6566_),
    .C(_6563_),
    .Y(_6575_)
);

NAND3X1 _16915_ (
    .A(_6573_),
    .B(_6574_),
    .C(_6575_),
    .Y(_6576_)
);

NAND3X1 _16916_ (
    .A(_6572_),
    .B(_6546_),
    .C(_6576_),
    .Y(_6577_)
);

AOI21X1 _16917_ (
    .A(_6164_),
    .B(_6185_),
    .C(_6189_),
    .Y(_6578_)
);

AOI21X1 _16918_ (
    .A(_6574_),
    .B(_6575_),
    .C(_6573_),
    .Y(_6579_)
);

AOI21X1 _16919_ (
    .A(_6564_),
    .B(_6570_),
    .C(_6548_),
    .Y(_6580_)
);

OAI21X1 _16920_ (
    .A(_6579_),
    .B(_6580_),
    .C(_6578_),
    .Y(_6581_)
);

NAND3X1 _16921_ (
    .A(_6577_),
    .B(_6581_),
    .C(_6545_),
    .Y(_6583_)
);

OR2X2 _16922_ (
    .A(_6539_),
    .B(_6544_),
    .Y(_6584_)
);

OAI21X1 _16923_ (
    .A(_6579_),
    .B(_6580_),
    .C(_6546_),
    .Y(_6585_)
);

NAND3X1 _16924_ (
    .A(_6572_),
    .B(_6576_),
    .C(_6578_),
    .Y(_6586_)
);

NAND3X1 _16925_ (
    .A(_6585_),
    .B(_6586_),
    .C(_6584_),
    .Y(_6587_)
);

OAI21X1 _16926_ (
    .A(_6251_),
    .B(_6258_),
    .C(_6260_),
    .Y(_6588_)
);

AOI21X1 _16927_ (
    .A(_6583_),
    .B(_6587_),
    .C(_6588_),
    .Y(_6589_)
);

AOI21X1 _16928_ (
    .A(_6585_),
    .B(_6586_),
    .C(_6584_),
    .Y(_6590_)
);

AOI21X1 _16929_ (
    .A(_6577_),
    .B(_6581_),
    .C(_6545_),
    .Y(_6591_)
);

AOI21X1 _16930_ (
    .A(_6221_),
    .B(_6259_),
    .C(_6256_),
    .Y(_6592_)
);

NOR3X1 _16931_ (
    .A(_6590_),
    .B(_6591_),
    .C(_6592_),
    .Y(_6594_)
);

OAI21X1 _16932_ (
    .A(_6594_),
    .B(_6589_),
    .C(_6512_),
    .Y(_6595_)
);

AND2X2 _16933_ (
    .A(_6200_),
    .B(_6192_),
    .Y(_6596_)
);

OAI21X1 _16934_ (
    .A(_6590_),
    .B(_6591_),
    .C(_6592_),
    .Y(_6597_)
);

NAND3X1 _16935_ (
    .A(_6583_),
    .B(_6588_),
    .C(_6587_),
    .Y(_6598_)
);

NAND3X1 _16936_ (
    .A(_6596_),
    .B(_6598_),
    .C(_6597_),
    .Y(_6599_)
);

NAND2X1 _16937_ (
    .A(_6599_),
    .B(_6595_),
    .Y(_6600_)
);

AOI21X1 _16938_ (
    .A(_6342_),
    .B(_6348_),
    .C(_6265_),
    .Y(_6601_)
);

OAI21X1 _16939_ (
    .A(_6359_),
    .B(_6601_),
    .C(_6349_),
    .Y(_6602_)
);

NAND2X1 _16940_ (
    .A(_6238_),
    .B(_6244_),
    .Y(_6603_)
);

NOR2X1 _16941_ (
    .A(_2379_),
    .B(_2465__bF$buf3),
    .Y(_6605_)
);

NAND2X1 _16942_ (
    .A(breg_13_bF$buf2),
    .B(areg_17_bF$buf1),
    .Y(_6606_)
);

OAI21X1 _16943_ (
    .A(_2586__bF$buf1),
    .B(_2884__bF$buf2),
    .C(_6561_),
    .Y(_6607_)
);

OAI21X1 _16944_ (
    .A(_6223_),
    .B(_6606_),
    .C(_6607_),
    .Y(_6608_)
);

XNOR2X1 _16945_ (
    .A(_6608_),
    .B(_6605_),
    .Y(_6609_)
);

OAI21X1 _16946_ (
    .A(_6236_),
    .B(_6227_),
    .C(_6230_),
    .Y(_6610_)
);

NAND2X1 _16947_ (
    .A(breg_11_bF$buf3),
    .B(areg_18_bF$buf2),
    .Y(_6611_)
);

INVX2 _16948_ (
    .A(_6611_),
    .Y(_6612_)
);

AND2X2 _16949_ (
    .A(breg_9_bF$buf1),
    .B(areg_20_bF$buf2),
    .Y(_6613_)
);

NAND2X1 _16950_ (
    .A(_6229_),
    .B(_6613_),
    .Y(_6614_)
);

OAI22X1 _16951_ (
    .A(_6044__bF$buf5),
    .B(_3958__bF$buf1),
    .C(_7217__bF$buf2),
    .D(_3402__bF$buf0),
    .Y(_6616_)
);

NAND3X1 _16952_ (
    .A(_6612_),
    .B(_6616_),
    .C(_6614_),
    .Y(_6617_)
);

NAND2X1 _16953_ (
    .A(breg_10_bF$buf3),
    .B(areg_20_bF$buf1),
    .Y(_6618_)
);

NOR2X1 _16954_ (
    .A(_6234_),
    .B(_6618_),
    .Y(_6619_)
);

NOR2X1 _16955_ (
    .A(_6229_),
    .B(_6613_),
    .Y(_6620_)
);

OAI21X1 _16956_ (
    .A(_6620_),
    .B(_6619_),
    .C(_6611_),
    .Y(_6621_)
);

NAND3X1 _16957_ (
    .A(_6610_),
    .B(_6617_),
    .C(_6621_),
    .Y(_6622_)
);

AOI21X1 _16958_ (
    .A(_6228_),
    .B(_6232_),
    .C(_6235_),
    .Y(_6623_)
);

OAI21X1 _16959_ (
    .A(_7217__bF$buf1),
    .B(_3402__bF$buf3),
    .C(_6613_),
    .Y(_6624_)
);

OAI21X1 _16960_ (
    .A(_6044__bF$buf4),
    .B(_3958__bF$buf0),
    .C(_6229_),
    .Y(_6625_)
);

AOI21X1 _16961_ (
    .A(_6624_),
    .B(_6625_),
    .C(_6611_),
    .Y(_6627_)
);

AOI21X1 _16962_ (
    .A(_6616_),
    .B(_6614_),
    .C(_6612_),
    .Y(_6628_)
);

OAI21X1 _16963_ (
    .A(_6627_),
    .B(_6628_),
    .C(_6623_),
    .Y(_6629_)
);

NAND3X1 _16964_ (
    .A(_6622_),
    .B(_6629_),
    .C(_6609_),
    .Y(_6630_)
);

INVX2 _16965_ (
    .A(_6605_),
    .Y(_6631_)
);

XNOR2X1 _16966_ (
    .A(_6608_),
    .B(_6631_),
    .Y(_6632_)
);

OAI21X1 _16967_ (
    .A(_6627_),
    .B(_6628_),
    .C(_6610_),
    .Y(_6633_)
);

NAND3X1 _16968_ (
    .A(_6623_),
    .B(_6617_),
    .C(_6621_),
    .Y(_6634_)
);

NAND3X1 _16969_ (
    .A(_6633_),
    .B(_6634_),
    .C(_6632_),
    .Y(_6635_)
);

OAI21X1 _16970_ (
    .A(_6281_),
    .B(_6287_),
    .C(_6289_),
    .Y(_6636_)
);

AOI21X1 _16971_ (
    .A(_6635_),
    .B(_6630_),
    .C(_6636_),
    .Y(_6638_)
);

AOI21X1 _16972_ (
    .A(_6633_),
    .B(_6634_),
    .C(_6632_),
    .Y(_6639_)
);

AOI21X1 _16973_ (
    .A(_6629_),
    .B(_6622_),
    .C(_6609_),
    .Y(_6640_)
);

AOI21X1 _16974_ (
    .A(_6267_),
    .B(_6288_),
    .C(_6284_),
    .Y(_6641_)
);

NOR3X1 _16975_ (
    .A(_6639_),
    .B(_6640_),
    .C(_6641_),
    .Y(_6642_)
);

OAI21X1 _16976_ (
    .A(_6642_),
    .B(_6638_),
    .C(_6603_),
    .Y(_6643_)
);

AND2X2 _16977_ (
    .A(_6244_),
    .B(_6238_),
    .Y(_6644_)
);

OAI21X1 _16978_ (
    .A(_6639_),
    .B(_6640_),
    .C(_6641_),
    .Y(_6645_)
);

NAND3X1 _16979_ (
    .A(_6630_),
    .B(_6635_),
    .C(_6636_),
    .Y(_6646_)
);

NAND3X1 _16980_ (
    .A(_6644_),
    .B(_6645_),
    .C(_6646_),
    .Y(_6647_)
);

NAND2X1 _16981_ (
    .A(_6647_),
    .B(_6643_),
    .Y(_6648_)
);

AOI21X1 _16982_ (
    .A(_6334_),
    .B(_6329_),
    .C(_6293_),
    .Y(_6649_)
);

OAI21X1 _16983_ (
    .A(_6345_),
    .B(_6649_),
    .C(_6335_),
    .Y(_6650_)
);

NAND2X1 _16984_ (
    .A(breg_7_bF$buf0),
    .B(areg_22_bF$buf0),
    .Y(_6651_)
);

OAI21X1 _16985_ (
    .A(_6266_),
    .B(_6651_),
    .C(_6273_),
    .Y(_6652_)
);

NOR2X1 _16986_ (
    .A(_5420__bF$buf0),
    .B(_3961__bF$buf3),
    .Y(_6653_)
);

AND2X2 _16987_ (
    .A(breg_7_bF$buf5),
    .B(areg_22_bF$buf4),
    .Y(_6654_)
);

AND2X2 _16988_ (
    .A(breg_6_bF$buf4),
    .B(areg_23_bF$buf1),
    .Y(_6655_)
);

NAND2X1 _16989_ (
    .A(_6654_),
    .B(_6655_),
    .Y(_6656_)
);

OAI21X1 _16990_ (
    .A(_5453__bF$buf5),
    .B(_4541__bF$buf1),
    .C(_6651_),
    .Y(_6657_)
);

NAND3X1 _16991_ (
    .A(_6653_),
    .B(_6657_),
    .C(_6656_),
    .Y(_6660_)
);

INVX1 _16992_ (
    .A(_6653_),
    .Y(_6661_)
);

OAI21X1 _16993_ (
    .A(_4116__bF$buf1),
    .B(_4551__bF$buf0),
    .C(_6655_),
    .Y(_6662_)
);

OAI21X1 _16994_ (
    .A(_5453__bF$buf4),
    .B(_4541__bF$buf0),
    .C(_6654_),
    .Y(_6663_)
);

NAND3X1 _16995_ (
    .A(_6662_),
    .B(_6663_),
    .C(_6661_),
    .Y(_6664_)
);

OAI21X1 _16996_ (
    .A(_6304_),
    .B(_6294_),
    .C(_6299_),
    .Y(_6665_)
);

AOI21X1 _16997_ (
    .A(_6660_),
    .B(_6664_),
    .C(_6665_),
    .Y(_6666_)
);

AOI21X1 _16998_ (
    .A(_6662_),
    .B(_6663_),
    .C(_6661_),
    .Y(_6667_)
);

AOI21X1 _16999_ (
    .A(_6657_),
    .B(_6656_),
    .C(_6653_),
    .Y(_6668_)
);

AOI21X1 _17000_ (
    .A(_6295_),
    .B(_6301_),
    .C(_6303_),
    .Y(_6669_)
);

NOR3X1 _17001_ (
    .A(_6668_),
    .B(_6669_),
    .C(_6667_),
    .Y(_6671_)
);

OAI21X1 _17002_ (
    .A(_6671_),
    .B(_6666_),
    .C(_6652_),
    .Y(_6672_)
);

AND2X2 _17003_ (
    .A(_6273_),
    .B(_6271_),
    .Y(_6673_)
);

OAI21X1 _17004_ (
    .A(_6667_),
    .B(_6668_),
    .C(_6669_),
    .Y(_6674_)
);

NAND3X1 _17005_ (
    .A(_6665_),
    .B(_6660_),
    .C(_6664_),
    .Y(_6675_)
);

NAND3X1 _17006_ (
    .A(_6673_),
    .B(_6675_),
    .C(_6674_),
    .Y(_6676_)
);

NAND2X1 _17007_ (
    .A(_6676_),
    .B(_6672_),
    .Y(_6677_)
);

AOI21X1 _17008_ (
    .A(_6321_),
    .B(_6316_),
    .C(_6307_),
    .Y(_6678_)
);

OAI21X1 _17009_ (
    .A(_6678_),
    .B(_6331_),
    .C(_6322_),
    .Y(_6679_)
);

NAND2X1 _17010_ (
    .A(breg_5_bF$buf0),
    .B(areg_24_bF$buf1),
    .Y(_6680_)
);

INVX1 _17011_ (
    .A(_6680_),
    .Y(_6682_)
);

NAND2X1 _17012_ (
    .A(breg_4_bF$buf3),
    .B(areg_25_bF$buf2),
    .Y(_6683_)
);

NAND2X1 _17013_ (
    .A(breg_3_bF$buf5),
    .B(areg_26_bF$buf4),
    .Y(_6684_)
);

OR2X2 _17014_ (
    .A(_6683_),
    .B(_6684_),
    .Y(_6685_)
);

INVX8 _17015_ (
    .A(areg_26_bF$buf3),
    .Y(_6686_)
);

OAI21X1 _17016_ (
    .A(_2365_),
    .B(_6686__bF$buf3),
    .C(_6683_),
    .Y(_6687_)
);

NAND3X1 _17017_ (
    .A(_6682_),
    .B(_6687_),
    .C(_6685_),
    .Y(_6688_)
);

NOR2X1 _17018_ (
    .A(_6683_),
    .B(_6684_),
    .Y(_6689_)
);

AND2X2 _17019_ (
    .A(_6683_),
    .B(_6684_),
    .Y(_6690_)
);

OAI21X1 _17020_ (
    .A(_6690_),
    .B(_6689_),
    .C(_6680_),
    .Y(_6691_)
);

AND2X2 _17021_ (
    .A(_6688_),
    .B(_6691_),
    .Y(_6693_)
);

OAI21X1 _17022_ (
    .A(_6309_),
    .B(_6314_),
    .C(_6313_),
    .Y(_6694_)
);

NAND2X1 _17023_ (
    .A(breg_2_bF$buf4),
    .B(areg_27_bF$buf5),
    .Y(_6695_)
);

INVX2 _17024_ (
    .A(_6695_),
    .Y(_6696_)
);

AND2X2 _17025_ (
    .A(breg_1_bF$buf2),
    .B(areg_28_bF$buf2),
    .Y(_6697_)
);

AND2X2 _17026_ (
    .A(breg_0_bF$buf1),
    .B(areg_29_bF$buf5),
    .Y(_6698_)
);

NAND2X1 _17027_ (
    .A(_6697_),
    .B(_6698_),
    .Y(_6699_)
);

AOI22X1 _17028_ (
    .A(breg_0_bF$buf0),
    .B(areg_29_bF$buf4),
    .C(breg_1_bF$buf1),
    .D(areg_28_bF$buf1),
    .Y(_6700_)
);

INVX2 _17029_ (
    .A(_6700_),
    .Y(_6701_)
);

NAND3X1 _17030_ (
    .A(_6696_),
    .B(_6701_),
    .C(_6699_),
    .Y(_6702_)
);

NAND2X1 _17031_ (
    .A(breg_1_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_6704_)
);

NAND2X1 _17032_ (
    .A(breg_0_bF$buf6),
    .B(areg_29_bF$buf3),
    .Y(_6705_)
);

NOR2X1 _17033_ (
    .A(_6704_),
    .B(_6705_),
    .Y(_6706_)
);

OAI21X1 _17034_ (
    .A(_6706_),
    .B(_6700_),
    .C(_6695_),
    .Y(_6707_)
);

NAND3X1 _17035_ (
    .A(_6694_),
    .B(_6707_),
    .C(_6702_),
    .Y(_6708_)
);

AOI21X1 _17036_ (
    .A(_6310_),
    .B(_6315_),
    .C(_6320_),
    .Y(_6709_)
);

NAND3X1 _17037_ (
    .A(breg_0_bF$buf5),
    .B(areg_29_bF$buf2),
    .C(_6704_),
    .Y(_6710_)
);

NAND2X1 _17038_ (
    .A(_6705_),
    .B(_6697_),
    .Y(_6711_)
);

AOI21X1 _17039_ (
    .A(_6710_),
    .B(_6711_),
    .C(_6695_),
    .Y(_6712_)
);

AOI21X1 _17040_ (
    .A(_6701_),
    .B(_6699_),
    .C(_6696_),
    .Y(_6713_)
);

OAI21X1 _17041_ (
    .A(_6713_),
    .B(_6712_),
    .C(_6709_),
    .Y(_6715_)
);

NAND3X1 _17042_ (
    .A(_6708_),
    .B(_6715_),
    .C(_6693_),
    .Y(_6716_)
);

NAND2X1 _17043_ (
    .A(_6691_),
    .B(_6688_),
    .Y(_6717_)
);

OAI21X1 _17044_ (
    .A(_6713_),
    .B(_6712_),
    .C(_6694_),
    .Y(_6718_)
);

NAND3X1 _17045_ (
    .A(_6707_),
    .B(_6709_),
    .C(_6702_),
    .Y(_6719_)
);

NAND3X1 _17046_ (
    .A(_6717_),
    .B(_6719_),
    .C(_6718_),
    .Y(_6720_)
);

NAND3X1 _17047_ (
    .A(_6679_),
    .B(_6720_),
    .C(_6716_),
    .Y(_6721_)
);

NOR3X1 _17048_ (
    .A(_6326_),
    .B(_6323_),
    .C(_6327_),
    .Y(_6722_)
);

AOI21X1 _17049_ (
    .A(_6306_),
    .B(_6328_),
    .C(_6722_),
    .Y(_6723_)
);

AOI21X1 _17050_ (
    .A(_6719_),
    .B(_6718_),
    .C(_6717_),
    .Y(_6724_)
);

AOI21X1 _17051_ (
    .A(_6708_),
    .B(_6715_),
    .C(_6693_),
    .Y(_6726_)
);

OAI21X1 _17052_ (
    .A(_6724_),
    .B(_6726_),
    .C(_6723_),
    .Y(_6727_)
);

NAND3X1 _17053_ (
    .A(_6721_),
    .B(_6727_),
    .C(_6677_),
    .Y(_6728_)
);

NAND3X1 _17054_ (
    .A(_6652_),
    .B(_6675_),
    .C(_6674_),
    .Y(_6729_)
);

OAI21X1 _17055_ (
    .A(_6671_),
    .B(_6666_),
    .C(_6673_),
    .Y(_6730_)
);

NAND2X1 _17056_ (
    .A(_6729_),
    .B(_6730_),
    .Y(_6731_)
);

OAI21X1 _17057_ (
    .A(_6724_),
    .B(_6726_),
    .C(_6679_),
    .Y(_6732_)
);

NAND3X1 _17058_ (
    .A(_6716_),
    .B(_6720_),
    .C(_6723_),
    .Y(_6733_)
);

NAND3X1 _17059_ (
    .A(_6733_),
    .B(_6732_),
    .C(_6731_),
    .Y(_6734_)
);

NAND3X1 _17060_ (
    .A(_6728_),
    .B(_6734_),
    .C(_6650_),
    .Y(_6735_)
);

NOR3X1 _17061_ (
    .A(_6338_),
    .B(_6339_),
    .C(_6337_),
    .Y(_6737_)
);

AOI21X1 _17062_ (
    .A(_6291_),
    .B(_6340_),
    .C(_6737_),
    .Y(_6738_)
);

AOI21X1 _17063_ (
    .A(_6733_),
    .B(_6732_),
    .C(_6731_),
    .Y(_6739_)
);

AOI21X1 _17064_ (
    .A(_6721_),
    .B(_6727_),
    .C(_6677_),
    .Y(_6740_)
);

OAI21X1 _17065_ (
    .A(_6739_),
    .B(_6740_),
    .C(_6738_),
    .Y(_6741_)
);

NAND3X1 _17066_ (
    .A(_6735_),
    .B(_6741_),
    .C(_6648_),
    .Y(_6742_)
);

NAND3X1 _17067_ (
    .A(_6603_),
    .B(_6645_),
    .C(_6646_),
    .Y(_6743_)
);

OAI21X1 _17068_ (
    .A(_6642_),
    .B(_6638_),
    .C(_6644_),
    .Y(_6744_)
);

NAND2X1 _17069_ (
    .A(_6743_),
    .B(_6744_),
    .Y(_6745_)
);

OAI21X1 _17070_ (
    .A(_6739_),
    .B(_6740_),
    .C(_6650_),
    .Y(_6746_)
);

NAND3X1 _17071_ (
    .A(_6728_),
    .B(_6734_),
    .C(_6738_),
    .Y(_6748_)
);

NAND3X1 _17072_ (
    .A(_6748_),
    .B(_6745_),
    .C(_6746_),
    .Y(_6749_)
);

NAND3X1 _17073_ (
    .A(_6742_),
    .B(_6749_),
    .C(_6602_),
    .Y(_6750_)
);

NOR3X1 _17074_ (
    .A(_6353_),
    .B(_6354_),
    .C(_6351_),
    .Y(_6751_)
);

AOI21X1 _17075_ (
    .A(_6262_),
    .B(_6355_),
    .C(_6751_),
    .Y(_6752_)
);

AOI21X1 _17076_ (
    .A(_6748_),
    .B(_6746_),
    .C(_6745_),
    .Y(_6753_)
);

AOI21X1 _17077_ (
    .A(_6735_),
    .B(_6741_),
    .C(_6648_),
    .Y(_6754_)
);

OAI21X1 _17078_ (
    .A(_6753_),
    .B(_6754_),
    .C(_6752_),
    .Y(_6755_)
);

NAND3X1 _17079_ (
    .A(_6750_),
    .B(_6755_),
    .C(_6600_),
    .Y(_6756_)
);

NAND3X1 _17080_ (
    .A(_6512_),
    .B(_6598_),
    .C(_6597_),
    .Y(_6757_)
);

OAI21X1 _17081_ (
    .A(_6594_),
    .B(_6589_),
    .C(_6596_),
    .Y(_6759_)
);

NAND2X1 _17082_ (
    .A(_6757_),
    .B(_6759_),
    .Y(_6760_)
);

OAI21X1 _17083_ (
    .A(_6753_),
    .B(_6754_),
    .C(_6602_),
    .Y(_6761_)
);

NAND3X1 _17084_ (
    .A(_6742_),
    .B(_6749_),
    .C(_6752_),
    .Y(_6762_)
);

NAND3X1 _17085_ (
    .A(_6761_),
    .B(_6762_),
    .C(_6760_),
    .Y(_6763_)
);

NAND3X1 _17086_ (
    .A(_6756_),
    .B(_6763_),
    .C(_6511_),
    .Y(_6764_)
);

NOR3X1 _17087_ (
    .A(_6367_),
    .B(_6368_),
    .C(_6366_),
    .Y(_6765_)
);

AOI21X1 _17088_ (
    .A(_6217_),
    .B(_6369_),
    .C(_6765_),
    .Y(_6766_)
);

AOI21X1 _17089_ (
    .A(_6762_),
    .B(_6761_),
    .C(_6760_),
    .Y(_6767_)
);

AOI21X1 _17090_ (
    .A(_6750_),
    .B(_6755_),
    .C(_6600_),
    .Y(_6768_)
);

OAI21X1 _17091_ (
    .A(_6767_),
    .B(_6768_),
    .C(_6766_),
    .Y(_6770_)
);

NAND3X1 _17092_ (
    .A(_6764_),
    .B(_6770_),
    .C(_6509_),
    .Y(_6771_)
);

NAND3X1 _17093_ (
    .A(_6424_),
    .B(_6507_),
    .C(_6506_),
    .Y(_6772_)
);

OAI21X1 _17094_ (
    .A(_6498_),
    .B(_6502_),
    .C(_6504_),
    .Y(_6773_)
);

NAND2X1 _17095_ (
    .A(_6772_),
    .B(_6773_),
    .Y(_6774_)
);

NOR3X1 _17096_ (
    .A(_6767_),
    .B(_6768_),
    .C(_6766_),
    .Y(_6775_)
);

AOI21X1 _17097_ (
    .A(_6756_),
    .B(_6763_),
    .C(_6511_),
    .Y(_6776_)
);

OAI21X1 _17098_ (
    .A(_6775_),
    .B(_6776_),
    .C(_6774_),
    .Y(_6777_)
);

NAND3X1 _17099_ (
    .A(_6423_),
    .B(_6771_),
    .C(_6777_),
    .Y(_6778_)
);

NOR3X1 _17100_ (
    .A(_6381_),
    .B(_6382_),
    .C(_6380_),
    .Y(_6779_)
);

AOI21X1 _17101_ (
    .A(_6383_),
    .B(_6127_),
    .C(_6779_),
    .Y(_6781_)
);

OAI21X1 _17102_ (
    .A(_6767_),
    .B(_6768_),
    .C(_6511_),
    .Y(_6782_)
);

NAND3X1 _17103_ (
    .A(_6756_),
    .B(_6763_),
    .C(_6766_),
    .Y(_6783_)
);

AOI21X1 _17104_ (
    .A(_6783_),
    .B(_6782_),
    .C(_6774_),
    .Y(_6784_)
);

AOI21X1 _17105_ (
    .A(_6764_),
    .B(_6770_),
    .C(_6509_),
    .Y(_6785_)
);

OAI21X1 _17106_ (
    .A(_6784_),
    .B(_6785_),
    .C(_6781_),
    .Y(_6786_)
);

NAND3X1 _17107_ (
    .A(_6786_),
    .B(_6421_),
    .C(_6778_),
    .Y(_6787_)
);

INVX1 _17108_ (
    .A(_6421_),
    .Y(_6788_)
);

OAI21X1 _17109_ (
    .A(_6784_),
    .B(_6785_),
    .C(_6423_),
    .Y(_6789_)
);

NAND3X1 _17110_ (
    .A(_6771_),
    .B(_6781_),
    .C(_6777_),
    .Y(_6790_)
);

NAND3X1 _17111_ (
    .A(_6788_),
    .B(_6789_),
    .C(_6790_),
    .Y(_6792_)
);

NAND3X1 _17112_ (
    .A(_6787_),
    .B(_6420_),
    .C(_6792_),
    .Y(_6793_)
);

AOI21X1 _17113_ (
    .A(_6045_),
    .B(_6398_),
    .C(_6401_),
    .Y(_6794_)
);

AOI21X1 _17114_ (
    .A(_6789_),
    .B(_6790_),
    .C(_6788_),
    .Y(_6795_)
);

AOI21X1 _17115_ (
    .A(_6786_),
    .B(_6778_),
    .C(_6421_),
    .Y(_6796_)
);

OAI21X1 _17116_ (
    .A(_6795_),
    .B(_6796_),
    .C(_6794_),
    .Y(_6797_)
);

NAND3X1 _17117_ (
    .A(_6793_),
    .B(_6797_),
    .C(_6419_),
    .Y(_6798_)
);

OAI21X1 _17118_ (
    .A(_6795_),
    .B(_6796_),
    .C(_6420_),
    .Y(_6799_)
);

NAND3X1 _17119_ (
    .A(_6787_),
    .B(_6792_),
    .C(_6794_),
    .Y(_6800_)
);

NAND3X1 _17120_ (
    .A(_6800_),
    .B(_6799_),
    .C(_6404_),
    .Y(_6801_)
);

NAND2X1 _17121_ (
    .A(_6801_),
    .B(_6798_),
    .Y(_6803_)
);

XNOR2X1 _17122_ (
    .A(_6418_),
    .B(_6803_),
    .Y(_0_[29])
);

OAI21X1 _17123_ (
    .A(_6803_),
    .B(_6412_),
    .C(_6798_),
    .Y(_6804_)
);

NOR2X1 _17124_ (
    .A(_6416_),
    .B(_6803_),
    .Y(_6805_)
);

INVX1 _17125_ (
    .A(_6805_),
    .Y(_6806_)
);

NOR2X1 _17126_ (
    .A(_6806_),
    .B(_6042_),
    .Y(_6807_)
);

NOR2X1 _17127_ (
    .A(_6804_),
    .B(_6807_),
    .Y(_6808_)
);

INVX1 _17128_ (
    .A(_6793_),
    .Y(_6809_)
);

NAND2X1 _17129_ (
    .A(_6778_),
    .B(_6787_),
    .Y(_6810_)
);

OAI21X1 _17130_ (
    .A(_6502_),
    .B(_6504_),
    .C(_6506_),
    .Y(_6811_)
);

OAI21X1 _17131_ (
    .A(_6774_),
    .B(_6776_),
    .C(_6764_),
    .Y(_6813_)
);

AND2X2 _17132_ (
    .A(_6499_),
    .B(_6493_),
    .Y(_6814_)
);

INVX8 _17133_ (
    .A(breg[30]),
    .Y(_6815_)
);

NOR2X1 _17134_ (
    .A(_2376__bF$buf2),
    .B(_6815__bF$buf4),
    .Y(_6816_)
);

INVX2 _17135_ (
    .A(_6816_),
    .Y(_6817_)
);

NOR2X1 _17136_ (
    .A(_6051_),
    .B(_6430_),
    .Y(_6818_)
);

AOI21X1 _17137_ (
    .A(_6429_),
    .B(_6431_),
    .C(_6818_),
    .Y(_6819_)
);

NAND2X1 _17138_ (
    .A(areg_1_bF$buf2),
    .B(breg_29_bF$buf3),
    .Y(_6820_)
);

NAND2X1 _17139_ (
    .A(areg_3_bF$buf4),
    .B(breg_27_bF$buf3),
    .Y(_6821_)
);

NOR2X1 _17140_ (
    .A(_6430_),
    .B(_6821_),
    .Y(_6822_)
);

AND2X2 _17141_ (
    .A(areg_2_bF$buf4),
    .B(breg_28_bF$buf2),
    .Y(_6824_)
);

AND2X2 _17142_ (
    .A(areg_3_bF$buf3),
    .B(breg_27_bF$buf2),
    .Y(_6825_)
);

NOR2X1 _17143_ (
    .A(_6824_),
    .B(_6825_),
    .Y(_6826_)
);

NOR3X1 _17144_ (
    .A(_6820_),
    .B(_6822_),
    .C(_6826_),
    .Y(_6827_)
);

INVX2 _17145_ (
    .A(_6820_),
    .Y(_6828_)
);

NAND2X1 _17146_ (
    .A(_6824_),
    .B(_6825_),
    .Y(_6829_)
);

OAI21X1 _17147_ (
    .A(_2792_),
    .B(_5668__bF$buf3),
    .C(_6430_),
    .Y(_6830_)
);

AOI21X1 _17148_ (
    .A(_6830_),
    .B(_6829_),
    .C(_6828_),
    .Y(_6831_)
);

NOR3X1 _17149_ (
    .A(_6819_),
    .B(_6831_),
    .C(_6827_),
    .Y(_6832_)
);

INVX1 _17150_ (
    .A(_6819_),
    .Y(_6833_)
);

NAND3X1 _17151_ (
    .A(_6828_),
    .B(_6830_),
    .C(_6829_),
    .Y(_6835_)
);

INVX1 _17152_ (
    .A(_6831_),
    .Y(_6836_)
);

AOI21X1 _17153_ (
    .A(_6835_),
    .B(_6836_),
    .C(_6833_),
    .Y(_6837_)
);

NOR3X1 _17154_ (
    .A(_6817_),
    .B(_6832_),
    .C(_6837_),
    .Y(_6838_)
);

OAI21X1 _17155_ (
    .A(_6837_),
    .B(_6832_),
    .C(_6817_),
    .Y(_6839_)
);

INVX1 _17156_ (
    .A(_6839_),
    .Y(_6840_)
);

OAI21X1 _17157_ (
    .A(_6840_),
    .B(_6838_),
    .C(_6436_),
    .Y(_6841_)
);

INVX1 _17158_ (
    .A(_6838_),
    .Y(_6842_)
);

NAND3X1 _17159_ (
    .A(_6435_),
    .B(_6839_),
    .C(_6842_),
    .Y(_6843_)
);

AND2X2 _17160_ (
    .A(_6843_),
    .B(_6841_),
    .Y(_6844_)
);

AOI21X1 _17161_ (
    .A(_6466_),
    .B(_6470_),
    .C(_6478_),
    .Y(_6846_)
);

OAI21X1 _17162_ (
    .A(_6846_),
    .B(_6441_),
    .C(_6482_),
    .Y(_6847_)
);

NAND2X1 _17163_ (
    .A(_6458_),
    .B(_6466_),
    .Y(_6848_)
);

NAND2X1 _17164_ (
    .A(areg_5_bF$buf2),
    .B(breg_25_bF$buf2),
    .Y(_6849_)
);

OAI21X1 _17165_ (
    .A(_6442_),
    .B(_6849_),
    .C(_6451_),
    .Y(_6850_)
);

NAND2X1 _17166_ (
    .A(areg_4_bF$buf3),
    .B(breg_26_bF$buf0),
    .Y(_6851_)
);

INVX1 _17167_ (
    .A(_6851_),
    .Y(_6852_)
);

AND2X2 _17168_ (
    .A(areg_5_bF$buf1),
    .B(breg_25_bF$buf1),
    .Y(_6853_)
);

AND2X2 _17169_ (
    .A(areg_6_bF$buf3),
    .B(breg_24_bF$buf3),
    .Y(_6854_)
);

NAND2X1 _17170_ (
    .A(_6853_),
    .B(_6854_),
    .Y(_6855_)
);

NAND2X1 _17171_ (
    .A(areg_6_bF$buf2),
    .B(breg_24_bF$buf2),
    .Y(_6857_)
);

OAI21X1 _17172_ (
    .A(_2825__bF$buf1),
    .B(_5318_),
    .C(_6857_),
    .Y(_6858_)
);

NAND3X1 _17173_ (
    .A(_6852_),
    .B(_6858_),
    .C(_6855_),
    .Y(_6859_)
);

NOR2X1 _17174_ (
    .A(_6849_),
    .B(_6857_),
    .Y(_6860_)
);

NOR2X1 _17175_ (
    .A(_6853_),
    .B(_6854_),
    .Y(_6861_)
);

OAI21X1 _17176_ (
    .A(_6861_),
    .B(_6860_),
    .C(_6851_),
    .Y(_6862_)
);

NAND2X1 _17177_ (
    .A(areg_8_bF$buf2),
    .B(breg_22_bF$buf1),
    .Y(_6863_)
);

AND2X2 _17178_ (
    .A(_6455_),
    .B(_6514_),
    .Y(_6864_)
);

OAI22X1 _17179_ (
    .A(_6134_),
    .B(_6863_),
    .C(_6540_),
    .D(_6864_),
    .Y(_6865_)
);

NAND3X1 _17180_ (
    .A(_6859_),
    .B(_6862_),
    .C(_6865_),
    .Y(_6866_)
);

NOR3X1 _17181_ (
    .A(_6851_),
    .B(_6860_),
    .C(_6861_),
    .Y(_6868_)
);

AOI21X1 _17182_ (
    .A(_6858_),
    .B(_6855_),
    .C(_6852_),
    .Y(_6869_)
);

NOR2X1 _17183_ (
    .A(_6455_),
    .B(_6514_),
    .Y(_6870_)
);

OAI21X1 _17184_ (
    .A(_5190__bF$buf2),
    .B(_3781__bF$buf1),
    .C(_6455_),
    .Y(_6871_)
);

AOI21X1 _17185_ (
    .A(_6513_),
    .B(_6871_),
    .C(_6870_),
    .Y(_6872_)
);

OAI21X1 _17186_ (
    .A(_6868_),
    .B(_6869_),
    .C(_6872_),
    .Y(_6873_)
);

NAND3X1 _17187_ (
    .A(_6850_),
    .B(_6873_),
    .C(_6866_),
    .Y(_6874_)
);

INVX1 _17188_ (
    .A(_6850_),
    .Y(_6875_)
);

NAND3X1 _17189_ (
    .A(_6859_),
    .B(_6872_),
    .C(_6862_),
    .Y(_6876_)
);

OAI21X1 _17190_ (
    .A(_6868_),
    .B(_6869_),
    .C(_6865_),
    .Y(_6877_)
);

NAND3X1 _17191_ (
    .A(_6876_),
    .B(_6877_),
    .C(_6875_),
    .Y(_6879_)
);

AOI21X1 _17192_ (
    .A(_6532_),
    .B(_6536_),
    .C(_6518_),
    .Y(_6880_)
);

OAI21X1 _17193_ (
    .A(_6517_),
    .B(_6880_),
    .C(_6542_),
    .Y(_6881_)
);

NAND3X1 _17194_ (
    .A(_6874_),
    .B(_6881_),
    .C(_6879_),
    .Y(_6882_)
);

AOI21X1 _17195_ (
    .A(_6876_),
    .B(_6877_),
    .C(_6875_),
    .Y(_6883_)
);

AOI21X1 _17196_ (
    .A(_6873_),
    .B(_6866_),
    .C(_6850_),
    .Y(_6884_)
);

NOR3X1 _17197_ (
    .A(_6529_),
    .B(_6531_),
    .C(_6525_),
    .Y(_6885_)
);

AOI21X1 _17198_ (
    .A(_6543_),
    .B(_6541_),
    .C(_6885_),
    .Y(_6886_)
);

OAI21X1 _17199_ (
    .A(_6884_),
    .B(_6883_),
    .C(_6886_),
    .Y(_6887_)
);

NAND3X1 _17200_ (
    .A(_6848_),
    .B(_6882_),
    .C(_6887_),
    .Y(_6888_)
);

INVX2 _17201_ (
    .A(_6848_),
    .Y(_6890_)
);

NAND3X1 _17202_ (
    .A(_6874_),
    .B(_6879_),
    .C(_6886_),
    .Y(_6891_)
);

OAI21X1 _17203_ (
    .A(_6884_),
    .B(_6883_),
    .C(_6881_),
    .Y(_6892_)
);

NAND3X1 _17204_ (
    .A(_6891_),
    .B(_6892_),
    .C(_6890_),
    .Y(_6893_)
);

NAND3X1 _17205_ (
    .A(_6847_),
    .B(_6888_),
    .C(_6893_),
    .Y(_6894_)
);

NAND2X1 _17206_ (
    .A(_6466_),
    .B(_6470_),
    .Y(_6895_)
);

NOR2X1 _17207_ (
    .A(_6473_),
    .B(_6895_),
    .Y(_6896_)
);

AOI21X1 _17208_ (
    .A(_6481_),
    .B(_6484_),
    .C(_6896_),
    .Y(_6897_)
);

AOI21X1 _17209_ (
    .A(_6891_),
    .B(_6892_),
    .C(_6890_),
    .Y(_6898_)
);

AOI21X1 _17210_ (
    .A(_6882_),
    .B(_6887_),
    .C(_6848_),
    .Y(_6899_)
);

OAI21X1 _17211_ (
    .A(_6899_),
    .B(_6898_),
    .C(_6897_),
    .Y(_6901_)
);

NAND3X1 _17212_ (
    .A(_6894_),
    .B(_6844_),
    .C(_6901_),
    .Y(_6902_)
);

NAND2X1 _17213_ (
    .A(_6841_),
    .B(_6843_),
    .Y(_6903_)
);

OAI21X1 _17214_ (
    .A(_6899_),
    .B(_6898_),
    .C(_6847_),
    .Y(_6904_)
);

NAND3X1 _17215_ (
    .A(_6888_),
    .B(_6893_),
    .C(_6897_),
    .Y(_6905_)
);

NAND3X1 _17216_ (
    .A(_6903_),
    .B(_6904_),
    .C(_6905_),
    .Y(_6906_)
);

OAI21X1 _17217_ (
    .A(_6589_),
    .B(_6596_),
    .C(_6598_),
    .Y(_6907_)
);

NAND3X1 _17218_ (
    .A(_6902_),
    .B(_6907_),
    .C(_6906_),
    .Y(_6908_)
);

AOI21X1 _17219_ (
    .A(_6904_),
    .B(_6905_),
    .C(_6903_),
    .Y(_6909_)
);

AOI21X1 _17220_ (
    .A(_6894_),
    .B(_6901_),
    .C(_6844_),
    .Y(_6910_)
);

AOI21X1 _17221_ (
    .A(_6512_),
    .B(_6597_),
    .C(_6594_),
    .Y(_6912_)
);

OAI21X1 _17222_ (
    .A(_6909_),
    .B(_6910_),
    .C(_6912_),
    .Y(_6913_)
);

NAND3X1 _17223_ (
    .A(_6814_),
    .B(_6908_),
    .C(_6913_),
    .Y(_6914_)
);

NAND2X1 _17224_ (
    .A(_6493_),
    .B(_6499_),
    .Y(_6915_)
);

NAND3X1 _17225_ (
    .A(_6902_),
    .B(_6912_),
    .C(_6906_),
    .Y(_6916_)
);

OAI21X1 _17226_ (
    .A(_6909_),
    .B(_6910_),
    .C(_6907_),
    .Y(_6917_)
);

NAND3X1 _17227_ (
    .A(_6915_),
    .B(_6916_),
    .C(_6917_),
    .Y(_6918_)
);

NAND2X1 _17228_ (
    .A(_6914_),
    .B(_6918_),
    .Y(_6919_)
);

AOI21X1 _17229_ (
    .A(_6742_),
    .B(_6749_),
    .C(_6602_),
    .Y(_6920_)
);

OAI21X1 _17230_ (
    .A(_6760_),
    .B(_6920_),
    .C(_6750_),
    .Y(_6921_)
);

NAND2X1 _17231_ (
    .A(_6577_),
    .B(_6583_),
    .Y(_6923_)
);

INVX2 _17232_ (
    .A(_6923_),
    .Y(_6924_)
);

NAND2X1 _17233_ (
    .A(areg_7_bF$buf3),
    .B(breg_23_bF$buf0),
    .Y(_6925_)
);

INVX2 _17234_ (
    .A(_6925_),
    .Y(_6926_)
);

NAND2X1 _17235_ (
    .A(areg_9_bF$buf2),
    .B(breg_21_bF$buf1),
    .Y(_6927_)
);

NOR2X1 _17236_ (
    .A(_6863_),
    .B(_6927_),
    .Y(_6928_)
);

AND2X2 _17237_ (
    .A(_6863_),
    .B(_6927_),
    .Y(_6929_)
);

NOR2X1 _17238_ (
    .A(_6928_),
    .B(_6929_),
    .Y(_6930_)
);

XNOR2X1 _17239_ (
    .A(_6930_),
    .B(_6926_),
    .Y(_6931_)
);

OAI21X1 _17240_ (
    .A(_6520_),
    .B(_6535_),
    .C(_6526_),
    .Y(_6932_)
);

NAND2X1 _17241_ (
    .A(areg_10_bF$buf2),
    .B(breg_20_bF$buf1),
    .Y(_6934_)
);

NAND2X1 _17242_ (
    .A(areg_12_bF$buf4),
    .B(breg_18_bF$buf3),
    .Y(_6935_)
);

NOR2X1 _17243_ (
    .A(_6533_),
    .B(_6935_),
    .Y(_6936_)
);

AND2X2 _17244_ (
    .A(areg_11_bF$buf2),
    .B(breg_19_bF$buf3),
    .Y(_6937_)
);

AND2X2 _17245_ (
    .A(areg_12_bF$buf3),
    .B(breg_18_bF$buf2),
    .Y(_6938_)
);

NOR2X1 _17246_ (
    .A(_6937_),
    .B(_6938_),
    .Y(_6939_)
);

NOR3X1 _17247_ (
    .A(_6934_),
    .B(_6936_),
    .C(_6939_),
    .Y(_6940_)
);

INVX2 _17248_ (
    .A(_6934_),
    .Y(_6941_)
);

NAND2X1 _17249_ (
    .A(_6937_),
    .B(_6938_),
    .Y(_6942_)
);

OAI21X1 _17250_ (
    .A(_10869__bF$buf1),
    .B(_3529__bF$buf3),
    .C(_6533_),
    .Y(_6943_)
);

AOI21X1 _17251_ (
    .A(_6943_),
    .B(_6942_),
    .C(_6941_),
    .Y(_6945_)
);

OAI21X1 _17252_ (
    .A(_6940_),
    .B(_6945_),
    .C(_6932_),
    .Y(_6946_)
);

AOI21X1 _17253_ (
    .A(_6519_),
    .B(_6528_),
    .C(_6534_),
    .Y(_6947_)
);

NAND3X1 _17254_ (
    .A(_6941_),
    .B(_6943_),
    .C(_6942_),
    .Y(_6948_)
);

OAI21X1 _17255_ (
    .A(_6939_),
    .B(_6936_),
    .C(_6934_),
    .Y(_6949_)
);

NAND3X1 _17256_ (
    .A(_6947_),
    .B(_6948_),
    .C(_6949_),
    .Y(_6950_)
);

AOI21X1 _17257_ (
    .A(_6946_),
    .B(_6950_),
    .C(_6931_),
    .Y(_6951_)
);

XNOR2X1 _17258_ (
    .A(_6930_),
    .B(_6925_),
    .Y(_6952_)
);

NAND3X1 _17259_ (
    .A(_6948_),
    .B(_6949_),
    .C(_6932_),
    .Y(_6953_)
);

OAI21X1 _17260_ (
    .A(_6940_),
    .B(_6945_),
    .C(_6947_),
    .Y(_6954_)
);

AOI21X1 _17261_ (
    .A(_6954_),
    .B(_6953_),
    .C(_6952_),
    .Y(_6956_)
);

NOR2X1 _17262_ (
    .A(_6951_),
    .B(_6956_),
    .Y(_6957_)
);

AOI21X1 _17263_ (
    .A(_6556_),
    .B(_6559_),
    .C(_6563_),
    .Y(_6958_)
);

OAI21X1 _17264_ (
    .A(_6958_),
    .B(_6573_),
    .C(_6564_),
    .Y(_6959_)
);

NAND2X1 _17265_ (
    .A(_6554_),
    .B(_6556_),
    .Y(_6960_)
);

NAND2X1 _17266_ (
    .A(areg_13_bF$buf1),
    .B(breg_17_bF$buf0),
    .Y(_6961_)
);

INVX1 _17267_ (
    .A(_6961_),
    .Y(_6962_)
);

AND2X2 _17268_ (
    .A(areg_14_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_6963_)
);

AND2X2 _17269_ (
    .A(areg_15_bF$buf0),
    .B(breg_15_bF$buf1),
    .Y(_6964_)
);

NAND2X1 _17270_ (
    .A(_6963_),
    .B(_6964_),
    .Y(_6965_)
);

NAND2X1 _17271_ (
    .A(areg_14_bF$buf0),
    .B(breg_16_bF$buf2),
    .Y(_6967_)
);

OAI21X1 _17272_ (
    .A(_2465__bF$buf2),
    .B(_2362__bF$buf1),
    .C(_6967_),
    .Y(_6968_)
);

NAND3X1 _17273_ (
    .A(_6962_),
    .B(_6968_),
    .C(_6965_),
    .Y(_6969_)
);

NAND2X1 _17274_ (
    .A(areg_15_bF$buf4),
    .B(breg_15_bF$buf0),
    .Y(_6970_)
);

NOR2X1 _17275_ (
    .A(_6967_),
    .B(_6970_),
    .Y(_6971_)
);

NOR2X1 _17276_ (
    .A(_6963_),
    .B(_6964_),
    .Y(_6972_)
);

OAI21X1 _17277_ (
    .A(_6972_),
    .B(_6971_),
    .C(_6961_),
    .Y(_6973_)
);

NAND2X1 _17278_ (
    .A(breg_12_bF$buf1),
    .B(areg_17_bF$buf0),
    .Y(_6974_)
);

AND2X2 _17279_ (
    .A(_6561_),
    .B(_6974_),
    .Y(_6975_)
);

OAI22X1 _17280_ (
    .A(_6223_),
    .B(_6606_),
    .C(_6631_),
    .D(_6975_),
    .Y(_6976_)
);

NAND3X1 _17281_ (
    .A(_6969_),
    .B(_6973_),
    .C(_6976_),
    .Y(_6978_)
);

NOR3X1 _17282_ (
    .A(_6961_),
    .B(_6971_),
    .C(_6972_),
    .Y(_6979_)
);

AOI21X1 _17283_ (
    .A(_6968_),
    .B(_6965_),
    .C(_6962_),
    .Y(_6980_)
);

NOR2X1 _17284_ (
    .A(_6561_),
    .B(_6974_),
    .Y(_6981_)
);

AOI21X1 _17285_ (
    .A(_6605_),
    .B(_6607_),
    .C(_6981_),
    .Y(_6982_)
);

OAI21X1 _17286_ (
    .A(_6979_),
    .B(_6980_),
    .C(_6982_),
    .Y(_6983_)
);

NAND3X1 _17287_ (
    .A(_6960_),
    .B(_6983_),
    .C(_6978_),
    .Y(_6984_)
);

INVX2 _17288_ (
    .A(_6960_),
    .Y(_6985_)
);

NOR3X1 _17289_ (
    .A(_6980_),
    .B(_6982_),
    .C(_6979_),
    .Y(_6986_)
);

AOI21X1 _17290_ (
    .A(_6969_),
    .B(_6973_),
    .C(_6976_),
    .Y(_6987_)
);

OAI21X1 _17291_ (
    .A(_6986_),
    .B(_6987_),
    .C(_6985_),
    .Y(_6989_)
);

NAND3X1 _17292_ (
    .A(_6959_),
    .B(_6984_),
    .C(_6989_),
    .Y(_6990_)
);

INVX1 _17293_ (
    .A(_6959_),
    .Y(_6991_)
);

NAND3X1 _17294_ (
    .A(_6969_),
    .B(_6982_),
    .C(_6973_),
    .Y(_6992_)
);

OAI21X1 _17295_ (
    .A(_6979_),
    .B(_6980_),
    .C(_6976_),
    .Y(_6993_)
);

AOI21X1 _17296_ (
    .A(_6992_),
    .B(_6993_),
    .C(_6985_),
    .Y(_6994_)
);

AOI21X1 _17297_ (
    .A(_6983_),
    .B(_6978_),
    .C(_6960_),
    .Y(_6995_)
);

OAI21X1 _17298_ (
    .A(_6995_),
    .B(_6994_),
    .C(_6991_),
    .Y(_6996_)
);

NAND3X1 _17299_ (
    .A(_6957_),
    .B(_6990_),
    .C(_6996_),
    .Y(_6997_)
);

OR2X2 _17300_ (
    .A(_6951_),
    .B(_6956_),
    .Y(_6998_)
);

OAI21X1 _17301_ (
    .A(_6995_),
    .B(_6994_),
    .C(_6959_),
    .Y(_7000_)
);

NAND3X1 _17302_ (
    .A(_6989_),
    .B(_6984_),
    .C(_6991_),
    .Y(_7001_)
);

NAND3X1 _17303_ (
    .A(_7000_),
    .B(_6998_),
    .C(_7001_),
    .Y(_7002_)
);

OAI21X1 _17304_ (
    .A(_6638_),
    .B(_6644_),
    .C(_6646_),
    .Y(_7003_)
);

NAND3X1 _17305_ (
    .A(_6997_),
    .B(_7003_),
    .C(_7002_),
    .Y(_7004_)
);

AOI21X1 _17306_ (
    .A(_7000_),
    .B(_7001_),
    .C(_6998_),
    .Y(_7005_)
);

AOI21X1 _17307_ (
    .A(_6990_),
    .B(_6996_),
    .C(_6957_),
    .Y(_7006_)
);

AOI21X1 _17308_ (
    .A(_6603_),
    .B(_6645_),
    .C(_6642_),
    .Y(_7007_)
);

OAI21X1 _17309_ (
    .A(_7005_),
    .B(_7006_),
    .C(_7007_),
    .Y(_7008_)
);

NAND3X1 _17310_ (
    .A(_6924_),
    .B(_7004_),
    .C(_7008_),
    .Y(_7009_)
);

NAND3X1 _17311_ (
    .A(_6997_),
    .B(_7007_),
    .C(_7002_),
    .Y(_7010_)
);

OAI21X1 _17312_ (
    .A(_7005_),
    .B(_7006_),
    .C(_7003_),
    .Y(_7011_)
);

NAND3X1 _17313_ (
    .A(_6923_),
    .B(_7010_),
    .C(_7011_),
    .Y(_7012_)
);

NAND2X1 _17314_ (
    .A(_7009_),
    .B(_7012_),
    .Y(_7013_)
);

AOI21X1 _17315_ (
    .A(_6728_),
    .B(_6734_),
    .C(_6650_),
    .Y(_7014_)
);

OAI21X1 _17316_ (
    .A(_6745_),
    .B(_7014_),
    .C(_6735_),
    .Y(_7015_)
);

AND2X2 _17317_ (
    .A(_6630_),
    .B(_6622_),
    .Y(_7016_)
);

NAND2X1 _17318_ (
    .A(breg_14_bF$buf1),
    .B(areg_16_bF$buf1),
    .Y(_7017_)
);

NAND2X1 _17319_ (
    .A(breg_12_bF$buf0),
    .B(areg_18_bF$buf1),
    .Y(_7018_)
);

NOR2X1 _17320_ (
    .A(_6606_),
    .B(_7018_),
    .Y(_7019_)
);

AND2X2 _17321_ (
    .A(_6606_),
    .B(_7018_),
    .Y(_7021_)
);

NOR2X1 _17322_ (
    .A(_7019_),
    .B(_7021_),
    .Y(_7022_)
);

XNOR2X1 _17323_ (
    .A(_7022_),
    .B(_7017_),
    .Y(_7023_)
);

OAI21X1 _17324_ (
    .A(_6620_),
    .B(_6611_),
    .C(_6614_),
    .Y(_7024_)
);

NAND2X1 _17325_ (
    .A(breg_11_bF$buf2),
    .B(areg_19_bF$buf2),
    .Y(_7025_)
);

INVX2 _17326_ (
    .A(_7025_),
    .Y(_7026_)
);

AND2X2 _17327_ (
    .A(breg_10_bF$buf2),
    .B(areg_20_bF$buf0),
    .Y(_7027_)
);

AND2X2 _17328_ (
    .A(breg_9_bF$buf0),
    .B(areg_21_bF$buf3),
    .Y(_7028_)
);

NAND2X1 _17329_ (
    .A(_7027_),
    .B(_7028_),
    .Y(_7029_)
);

OAI21X1 _17330_ (
    .A(_6044__bF$buf3),
    .B(_3961__bF$buf2),
    .C(_6618_),
    .Y(_7030_)
);

NAND3X1 _17331_ (
    .A(_7026_),
    .B(_7030_),
    .C(_7029_),
    .Y(_7033_)
);

NAND2X1 _17332_ (
    .A(breg_9_bF$buf5),
    .B(areg_21_bF$buf2),
    .Y(_7034_)
);

NOR2X1 _17333_ (
    .A(_6618_),
    .B(_7034_),
    .Y(_7035_)
);

NOR2X1 _17334_ (
    .A(_7027_),
    .B(_7028_),
    .Y(_7036_)
);

OAI21X1 _17335_ (
    .A(_7036_),
    .B(_7035_),
    .C(_7025_),
    .Y(_7037_)
);

NAND3X1 _17336_ (
    .A(_7033_),
    .B(_7024_),
    .C(_7037_),
    .Y(_7038_)
);

AOI21X1 _17337_ (
    .A(_6612_),
    .B(_6616_),
    .C(_6619_),
    .Y(_7039_)
);

NOR3X1 _17338_ (
    .A(_7025_),
    .B(_7035_),
    .C(_7036_),
    .Y(_7040_)
);

AOI21X1 _17339_ (
    .A(_7030_),
    .B(_7029_),
    .C(_7026_),
    .Y(_7041_)
);

OAI21X1 _17340_ (
    .A(_7040_),
    .B(_7041_),
    .C(_7039_),
    .Y(_7042_)
);

NAND3X1 _17341_ (
    .A(_7038_),
    .B(_7042_),
    .C(_7023_),
    .Y(_7044_)
);

INVX2 _17342_ (
    .A(_7017_),
    .Y(_7045_)
);

XNOR2X1 _17343_ (
    .A(_7022_),
    .B(_7045_),
    .Y(_7046_)
);

OAI21X1 _17344_ (
    .A(_7040_),
    .B(_7041_),
    .C(_7024_),
    .Y(_7047_)
);

NAND3X1 _17345_ (
    .A(_7039_),
    .B(_7033_),
    .C(_7037_),
    .Y(_7048_)
);

NAND3X1 _17346_ (
    .A(_7048_),
    .B(_7047_),
    .C(_7046_),
    .Y(_7049_)
);

OAI21X1 _17347_ (
    .A(_6666_),
    .B(_6673_),
    .C(_6675_),
    .Y(_7050_)
);

NAND3X1 _17348_ (
    .A(_7050_),
    .B(_7044_),
    .C(_7049_),
    .Y(_7051_)
);

AOI21X1 _17349_ (
    .A(_7048_),
    .B(_7047_),
    .C(_7046_),
    .Y(_7052_)
);

AOI21X1 _17350_ (
    .A(_7038_),
    .B(_7042_),
    .C(_7023_),
    .Y(_7053_)
);

AOI21X1 _17351_ (
    .A(_6652_),
    .B(_6674_),
    .C(_6671_),
    .Y(_7055_)
);

OAI21X1 _17352_ (
    .A(_7052_),
    .B(_7053_),
    .C(_7055_),
    .Y(_7056_)
);

NAND3X1 _17353_ (
    .A(_7016_),
    .B(_7051_),
    .C(_7056_),
    .Y(_7057_)
);

NAND2X1 _17354_ (
    .A(_6622_),
    .B(_6630_),
    .Y(_7058_)
);

NAND3X1 _17355_ (
    .A(_7055_),
    .B(_7044_),
    .C(_7049_),
    .Y(_7059_)
);

OAI21X1 _17356_ (
    .A(_7052_),
    .B(_7053_),
    .C(_7050_),
    .Y(_7060_)
);

NAND3X1 _17357_ (
    .A(_7058_),
    .B(_7059_),
    .C(_7060_),
    .Y(_7061_)
);

NAND2X1 _17358_ (
    .A(_7057_),
    .B(_7061_),
    .Y(_7062_)
);

AOI21X1 _17359_ (
    .A(_6720_),
    .B(_6716_),
    .C(_6679_),
    .Y(_7063_)
);

OAI21X1 _17360_ (
    .A(_6731_),
    .B(_7063_),
    .C(_6721_),
    .Y(_7064_)
);

AND2X2 _17361_ (
    .A(_6660_),
    .B(_6656_),
    .Y(_7066_)
);

NAND2X1 _17362_ (
    .A(breg[8]),
    .B(areg_22_bF$buf3),
    .Y(_7067_)
);

INVX1 _17363_ (
    .A(_7067_),
    .Y(_7068_)
);

AND2X2 _17364_ (
    .A(breg_7_bF$buf4),
    .B(areg_23_bF$buf0),
    .Y(_7069_)
);

AND2X2 _17365_ (
    .A(breg_6_bF$buf3),
    .B(areg_24_bF$buf0),
    .Y(_7070_)
);

NAND2X1 _17366_ (
    .A(_7069_),
    .B(_7070_),
    .Y(_7071_)
);

OAI22X1 _17367_ (
    .A(_5453__bF$buf3),
    .B(_5921__bF$buf2),
    .C(_4116__bF$buf0),
    .D(_4541__bF$buf4),
    .Y(_7072_)
);

NAND3X1 _17368_ (
    .A(_7068_),
    .B(_7072_),
    .C(_7071_),
    .Y(_7073_)
);

OAI21X1 _17369_ (
    .A(_4116__bF$buf4),
    .B(_4541__bF$buf3),
    .C(_7070_),
    .Y(_7074_)
);

OAI21X1 _17370_ (
    .A(_5453__bF$buf2),
    .B(_5921__bF$buf1),
    .C(_7069_),
    .Y(_7075_)
);

NAND3X1 _17371_ (
    .A(_7067_),
    .B(_7074_),
    .C(_7075_),
    .Y(_7077_)
);

OAI21X1 _17372_ (
    .A(_6690_),
    .B(_6680_),
    .C(_6685_),
    .Y(_7078_)
);

NAND3X1 _17373_ (
    .A(_7073_),
    .B(_7077_),
    .C(_7078_),
    .Y(_7079_)
);

AOI21X1 _17374_ (
    .A(_7074_),
    .B(_7075_),
    .C(_7067_),
    .Y(_7080_)
);

AOI21X1 _17375_ (
    .A(_7072_),
    .B(_7071_),
    .C(_7068_),
    .Y(_7081_)
);

AOI21X1 _17376_ (
    .A(_6682_),
    .B(_6687_),
    .C(_6689_),
    .Y(_7082_)
);

OAI21X1 _17377_ (
    .A(_7080_),
    .B(_7081_),
    .C(_7082_),
    .Y(_7083_)
);

NAND3X1 _17378_ (
    .A(_7066_),
    .B(_7079_),
    .C(_7083_),
    .Y(_7084_)
);

INVX1 _17379_ (
    .A(_6655_),
    .Y(_7085_)
);

OAI21X1 _17380_ (
    .A(_6651_),
    .B(_7085_),
    .C(_6660_),
    .Y(_7086_)
);

NOR3X1 _17381_ (
    .A(_7081_),
    .B(_7082_),
    .C(_7080_),
    .Y(_7088_)
);

AOI21X1 _17382_ (
    .A(_7073_),
    .B(_7077_),
    .C(_7078_),
    .Y(_7089_)
);

OAI21X1 _17383_ (
    .A(_7088_),
    .B(_7089_),
    .C(_7086_),
    .Y(_7090_)
);

NAND2X1 _17384_ (
    .A(_7084_),
    .B(_7090_),
    .Y(_7091_)
);

AOI21X1 _17385_ (
    .A(_6707_),
    .B(_6702_),
    .C(_6694_),
    .Y(_7092_)
);

OAI21X1 _17386_ (
    .A(_7092_),
    .B(_6717_),
    .C(_6708_),
    .Y(_7093_)
);

NAND2X1 _17387_ (
    .A(breg_5_bF$buf3),
    .B(areg_25_bF$buf1),
    .Y(_7094_)
);

INVX1 _17388_ (
    .A(_7094_),
    .Y(_7095_)
);

NAND2X1 _17389_ (
    .A(breg_4_bF$buf2),
    .B(areg_26_bF$buf2),
    .Y(_7096_)
);

NAND2X1 _17390_ (
    .A(breg_3_bF$buf4),
    .B(areg_27_bF$buf4),
    .Y(_7097_)
);

OR2X2 _17391_ (
    .A(_7096_),
    .B(_7097_),
    .Y(_7099_)
);

INVX8 _17392_ (
    .A(areg_27_bF$buf3),
    .Y(_7100_)
);

OAI21X1 _17393_ (
    .A(_2365_),
    .B(_7100__bF$buf3),
    .C(_7096_),
    .Y(_7101_)
);

NAND3X1 _17394_ (
    .A(_7095_),
    .B(_7101_),
    .C(_7099_),
    .Y(_7102_)
);

NOR2X1 _17395_ (
    .A(_7096_),
    .B(_7097_),
    .Y(_7103_)
);

AND2X2 _17396_ (
    .A(_7096_),
    .B(_7097_),
    .Y(_7104_)
);

OAI21X1 _17397_ (
    .A(_7104_),
    .B(_7103_),
    .C(_7094_),
    .Y(_7105_)
);

AND2X2 _17398_ (
    .A(_7102_),
    .B(_7105_),
    .Y(_7106_)
);

OAI21X1 _17399_ (
    .A(_6695_),
    .B(_6700_),
    .C(_6699_),
    .Y(_7107_)
);

NAND2X1 _17400_ (
    .A(breg_2_bF$buf3),
    .B(areg_28_bF$buf5),
    .Y(_7108_)
);

INVX2 _17401_ (
    .A(_7108_),
    .Y(_7110_)
);

AND2X2 _17402_ (
    .A(breg_1_bF$buf6),
    .B(areg_30_bF$buf5),
    .Y(_7111_)
);

NAND2X1 _17403_ (
    .A(_6698_),
    .B(_7111_),
    .Y(_7112_)
);

AOI22X1 _17404_ (
    .A(breg_0_bF$buf4),
    .B(areg_30_bF$buf4),
    .C(breg_1_bF$buf5),
    .D(areg_29_bF$buf1),
    .Y(_7113_)
);

INVX2 _17405_ (
    .A(_7113_),
    .Y(_7114_)
);

NAND3X1 _17406_ (
    .A(_7110_),
    .B(_7114_),
    .C(_7112_),
    .Y(_7115_)
);

NAND2X1 _17407_ (
    .A(breg_1_bF$buf4),
    .B(areg_30_bF$buf3),
    .Y(_7116_)
);

NOR2X1 _17408_ (
    .A(_6705_),
    .B(_7116_),
    .Y(_7117_)
);

OAI21X1 _17409_ (
    .A(_7117_),
    .B(_7113_),
    .C(_7108_),
    .Y(_7118_)
);

NAND3X1 _17410_ (
    .A(_7107_),
    .B(_7118_),
    .C(_7115_),
    .Y(_7119_)
);

AOI21X1 _17411_ (
    .A(_6696_),
    .B(_6701_),
    .C(_6706_),
    .Y(_7121_)
);

NAND2X1 _17412_ (
    .A(breg_1_bF$buf3),
    .B(areg_29_bF$buf0),
    .Y(_7122_)
);

NAND3X1 _17413_ (
    .A(breg_0_bF$buf3),
    .B(areg_30_bF$buf2),
    .C(_7122_),
    .Y(_7123_)
);

NAND2X1 _17414_ (
    .A(breg_0_bF$buf2),
    .B(areg_30_bF$buf1),
    .Y(_7124_)
);

NAND3X1 _17415_ (
    .A(breg_1_bF$buf2),
    .B(areg_29_bF$buf5),
    .C(_7124_),
    .Y(_7125_)
);

AOI21X1 _17416_ (
    .A(_7123_),
    .B(_7125_),
    .C(_7108_),
    .Y(_7126_)
);

AOI21X1 _17417_ (
    .A(_7114_),
    .B(_7112_),
    .C(_7110_),
    .Y(_7127_)
);

OAI21X1 _17418_ (
    .A(_7127_),
    .B(_7126_),
    .C(_7121_),
    .Y(_7128_)
);

NAND3X1 _17419_ (
    .A(_7119_),
    .B(_7128_),
    .C(_7106_),
    .Y(_7129_)
);

NAND2X1 _17420_ (
    .A(_7105_),
    .B(_7102_),
    .Y(_7130_)
);

OAI21X1 _17421_ (
    .A(_7127_),
    .B(_7126_),
    .C(_7107_),
    .Y(_7132_)
);

NAND3X1 _17422_ (
    .A(_7118_),
    .B(_7121_),
    .C(_7115_),
    .Y(_7133_)
);

NAND3X1 _17423_ (
    .A(_7130_),
    .B(_7133_),
    .C(_7132_),
    .Y(_7134_)
);

NAND3X1 _17424_ (
    .A(_7093_),
    .B(_7134_),
    .C(_7129_),
    .Y(_7135_)
);

NOR3X1 _17425_ (
    .A(_6712_),
    .B(_6709_),
    .C(_6713_),
    .Y(_7136_)
);

AOI21X1 _17426_ (
    .A(_6693_),
    .B(_6715_),
    .C(_7136_),
    .Y(_7137_)
);

AOI21X1 _17427_ (
    .A(_7133_),
    .B(_7132_),
    .C(_7130_),
    .Y(_7138_)
);

AOI21X1 _17428_ (
    .A(_7119_),
    .B(_7128_),
    .C(_7106_),
    .Y(_7139_)
);

OAI21X1 _17429_ (
    .A(_7138_),
    .B(_7139_),
    .C(_7137_),
    .Y(_7140_)
);

NAND3X1 _17430_ (
    .A(_7135_),
    .B(_7091_),
    .C(_7140_),
    .Y(_7141_)
);

NAND3X1 _17431_ (
    .A(_7086_),
    .B(_7079_),
    .C(_7083_),
    .Y(_7143_)
);

OAI21X1 _17432_ (
    .A(_7088_),
    .B(_7089_),
    .C(_7066_),
    .Y(_7144_)
);

NAND2X1 _17433_ (
    .A(_7143_),
    .B(_7144_),
    .Y(_7145_)
);

OAI21X1 _17434_ (
    .A(_7138_),
    .B(_7139_),
    .C(_7093_),
    .Y(_7146_)
);

NAND3X1 _17435_ (
    .A(_7129_),
    .B(_7134_),
    .C(_7137_),
    .Y(_7147_)
);

NAND3X1 _17436_ (
    .A(_7145_),
    .B(_7147_),
    .C(_7146_),
    .Y(_7148_)
);

NAND3X1 _17437_ (
    .A(_7141_),
    .B(_7148_),
    .C(_7064_),
    .Y(_7149_)
);

NOR3X1 _17438_ (
    .A(_6724_),
    .B(_6726_),
    .C(_6723_),
    .Y(_7150_)
);

AOI21X1 _17439_ (
    .A(_6677_),
    .B(_6727_),
    .C(_7150_),
    .Y(_7151_)
);

AOI21X1 _17440_ (
    .A(_7147_),
    .B(_7146_),
    .C(_7145_),
    .Y(_7152_)
);

AOI21X1 _17441_ (
    .A(_7135_),
    .B(_7140_),
    .C(_7091_),
    .Y(_7154_)
);

OAI21X1 _17442_ (
    .A(_7152_),
    .B(_7154_),
    .C(_7151_),
    .Y(_7155_)
);

NAND3X1 _17443_ (
    .A(_7149_),
    .B(_7062_),
    .C(_7155_),
    .Y(_7156_)
);

NAND3X1 _17444_ (
    .A(_7058_),
    .B(_7051_),
    .C(_7056_),
    .Y(_7157_)
);

NAND3X1 _17445_ (
    .A(_7016_),
    .B(_7059_),
    .C(_7060_),
    .Y(_7158_)
);

NAND2X1 _17446_ (
    .A(_7157_),
    .B(_7158_),
    .Y(_7159_)
);

OAI21X1 _17447_ (
    .A(_7152_),
    .B(_7154_),
    .C(_7064_),
    .Y(_7160_)
);

NAND3X1 _17448_ (
    .A(_7141_),
    .B(_7148_),
    .C(_7151_),
    .Y(_7161_)
);

NAND3X1 _17449_ (
    .A(_7159_),
    .B(_7161_),
    .C(_7160_),
    .Y(_7162_)
);

NAND3X1 _17450_ (
    .A(_7156_),
    .B(_7162_),
    .C(_7015_),
    .Y(_7163_)
);

NOR3X1 _17451_ (
    .A(_6739_),
    .B(_6740_),
    .C(_6738_),
    .Y(_7165_)
);

AOI21X1 _17452_ (
    .A(_6648_),
    .B(_6741_),
    .C(_7165_),
    .Y(_7166_)
);

AOI21X1 _17453_ (
    .A(_7161_),
    .B(_7160_),
    .C(_7159_),
    .Y(_7167_)
);

AOI21X1 _17454_ (
    .A(_7149_),
    .B(_7155_),
    .C(_7062_),
    .Y(_7168_)
);

OAI21X1 _17455_ (
    .A(_7167_),
    .B(_7168_),
    .C(_7166_),
    .Y(_7169_)
);

NAND3X1 _17456_ (
    .A(_7163_),
    .B(_7169_),
    .C(_7013_),
    .Y(_7170_)
);

NAND3X1 _17457_ (
    .A(_6923_),
    .B(_7004_),
    .C(_7008_),
    .Y(_7171_)
);

NAND3X1 _17458_ (
    .A(_6924_),
    .B(_7010_),
    .C(_7011_),
    .Y(_7172_)
);

NAND2X1 _17459_ (
    .A(_7171_),
    .B(_7172_),
    .Y(_7173_)
);

OAI21X1 _17460_ (
    .A(_7167_),
    .B(_7168_),
    .C(_7015_),
    .Y(_7174_)
);

NAND3X1 _17461_ (
    .A(_7156_),
    .B(_7162_),
    .C(_7166_),
    .Y(_7175_)
);

NAND3X1 _17462_ (
    .A(_7174_),
    .B(_7175_),
    .C(_7173_),
    .Y(_7176_)
);

NAND3X1 _17463_ (
    .A(_7170_),
    .B(_7176_),
    .C(_6921_),
    .Y(_7177_)
);

NOR3X1 _17464_ (
    .A(_6753_),
    .B(_6754_),
    .C(_6752_),
    .Y(_7178_)
);

AOI21X1 _17465_ (
    .A(_6600_),
    .B(_6755_),
    .C(_7178_),
    .Y(_7179_)
);

AOI21X1 _17466_ (
    .A(_7175_),
    .B(_7174_),
    .C(_7173_),
    .Y(_7180_)
);

AOI21X1 _17467_ (
    .A(_7163_),
    .B(_7169_),
    .C(_7013_),
    .Y(_7181_)
);

OAI21X1 _17468_ (
    .A(_7180_),
    .B(_7181_),
    .C(_7179_),
    .Y(_7182_)
);

NAND3X1 _17469_ (
    .A(_7177_),
    .B(_6919_),
    .C(_7182_),
    .Y(_7183_)
);

NAND3X1 _17470_ (
    .A(_6915_),
    .B(_6908_),
    .C(_6913_),
    .Y(_7184_)
);

NAND3X1 _17471_ (
    .A(_6814_),
    .B(_6916_),
    .C(_6917_),
    .Y(_7186_)
);

NAND2X1 _17472_ (
    .A(_7184_),
    .B(_7186_),
    .Y(_7187_)
);

OAI21X1 _17473_ (
    .A(_7180_),
    .B(_7181_),
    .C(_6921_),
    .Y(_7188_)
);

NAND3X1 _17474_ (
    .A(_7170_),
    .B(_7176_),
    .C(_7179_),
    .Y(_7189_)
);

NAND3X1 _17475_ (
    .A(_7189_),
    .B(_7187_),
    .C(_7188_),
    .Y(_7190_)
);

NAND3X1 _17476_ (
    .A(_7183_),
    .B(_7190_),
    .C(_6813_),
    .Y(_7191_)
);

AOI21X1 _17477_ (
    .A(_6509_),
    .B(_6770_),
    .C(_6775_),
    .Y(_7192_)
);

AOI21X1 _17478_ (
    .A(_7189_),
    .B(_7188_),
    .C(_7187_),
    .Y(_7193_)
);

AOI21X1 _17479_ (
    .A(_7177_),
    .B(_7182_),
    .C(_6919_),
    .Y(_7194_)
);

OAI21X1 _17480_ (
    .A(_7193_),
    .B(_7194_),
    .C(_7192_),
    .Y(_7195_)
);

NAND3X1 _17481_ (
    .A(_6811_),
    .B(_7191_),
    .C(_7195_),
    .Y(_7197_)
);

INVX1 _17482_ (
    .A(_6811_),
    .Y(_7198_)
);

NOR3X1 _17483_ (
    .A(_7193_),
    .B(_7194_),
    .C(_7192_),
    .Y(_7199_)
);

AOI21X1 _17484_ (
    .A(_7183_),
    .B(_7190_),
    .C(_6813_),
    .Y(_7200_)
);

OAI21X1 _17485_ (
    .A(_7199_),
    .B(_7200_),
    .C(_7198_),
    .Y(_7201_)
);

NAND3X1 _17486_ (
    .A(_7197_),
    .B(_7201_),
    .C(_6810_),
    .Y(_7202_)
);

INVX1 _17487_ (
    .A(_6778_),
    .Y(_7203_)
);

AOI21X1 _17488_ (
    .A(_6421_),
    .B(_6786_),
    .C(_7203_),
    .Y(_7204_)
);

INVX1 _17489_ (
    .A(_7197_),
    .Y(_7205_)
);

AOI21X1 _17490_ (
    .A(_7191_),
    .B(_7195_),
    .C(_6811_),
    .Y(_7206_)
);

OAI21X1 _17491_ (
    .A(_7205_),
    .B(_7206_),
    .C(_7204_),
    .Y(_7208_)
);

NAND3X1 _17492_ (
    .A(_7208_),
    .B(_6809_),
    .C(_7202_),
    .Y(_7209_)
);

OAI21X1 _17493_ (
    .A(_7205_),
    .B(_7206_),
    .C(_6810_),
    .Y(_7210_)
);

NAND3X1 _17494_ (
    .A(_7197_),
    .B(_7201_),
    .C(_7204_),
    .Y(_7211_)
);

NAND3X1 _17495_ (
    .A(_6793_),
    .B(_7211_),
    .C(_7210_),
    .Y(_7212_)
);

AND2X2 _17496_ (
    .A(_7209_),
    .B(_7212_),
    .Y(_7213_)
);

XNOR2X1 _17497_ (
    .A(_6808_),
    .B(_7213_),
    .Y(_0_[30])
);

NAND2X1 _17498_ (
    .A(_7212_),
    .B(_7209_),
    .Y(_7214_)
);

OAI21X1 _17499_ (
    .A(_6808_),
    .B(_7214_),
    .C(_7209_),
    .Y(_7215_)
);

NAND2X1 _17500_ (
    .A(_7197_),
    .B(_7201_),
    .Y(_7216_)
);

NOR2X1 _17501_ (
    .A(_7204_),
    .B(_7216_),
    .Y(_7218_)
);

INVX2 _17502_ (
    .A(_6843_),
    .Y(_7219_)
);

OAI21X1 _17503_ (
    .A(_7200_),
    .B(_7198_),
    .C(_7191_),
    .Y(_7220_)
);

NAND2X1 _17504_ (
    .A(_6908_),
    .B(_7184_),
    .Y(_7221_)
);

AOI21X1 _17505_ (
    .A(_7170_),
    .B(_7176_),
    .C(_6921_),
    .Y(_7222_)
);

OAI21X1 _17506_ (
    .A(_7187_),
    .B(_7222_),
    .C(_7177_),
    .Y(_7223_)
);

AND2X2 _17507_ (
    .A(_6902_),
    .B(_6894_),
    .Y(_7224_)
);

INVX8 _17508_ (
    .A(breg[31]),
    .Y(_7225_)
);

NOR2X1 _17509_ (
    .A(_2376__bF$buf1),
    .B(_7225__bF$buf4),
    .Y(_7226_)
);

INVX1 _17510_ (
    .A(_7226_),
    .Y(_7227_)
);

NOR2X1 _17511_ (
    .A(_6831_),
    .B(_6827_),
    .Y(_7229_)
);

NAND2X1 _17512_ (
    .A(_6833_),
    .B(_7229_),
    .Y(_7230_)
);

OAI21X1 _17513_ (
    .A(_6837_),
    .B(_6817_),
    .C(_7230_),
    .Y(_7231_)
);

NOR2X1 _17514_ (
    .A(_2661_),
    .B(_6815__bF$buf3),
    .Y(_7232_)
);

INVX2 _17515_ (
    .A(_7232_),
    .Y(_7233_)
);

OAI21X1 _17516_ (
    .A(_6826_),
    .B(_6820_),
    .C(_6829_),
    .Y(_7234_)
);

NAND2X1 _17517_ (
    .A(areg_2_bF$buf3),
    .B(breg_29_bF$buf2),
    .Y(_7235_)
);

INVX2 _17518_ (
    .A(_7235_),
    .Y(_7236_)
);

AND2X2 _17519_ (
    .A(areg_3_bF$buf2),
    .B(breg_28_bF$buf1),
    .Y(_7237_)
);

AND2X2 _17520_ (
    .A(areg_4_bF$buf2),
    .B(breg_27_bF$buf1),
    .Y(_7238_)
);

NAND2X1 _17521_ (
    .A(_7237_),
    .B(_7238_),
    .Y(_7240_)
);

OAI22X1 _17522_ (
    .A(_2562__bF$buf3),
    .B(_5668__bF$buf2),
    .C(_2792_),
    .D(_6050__bF$buf2),
    .Y(_7241_)
);

NAND3X1 _17523_ (
    .A(_7236_),
    .B(_7241_),
    .C(_7240_),
    .Y(_7242_)
);

NAND2X1 _17524_ (
    .A(areg_4_bF$buf1),
    .B(breg_28_bF$buf0),
    .Y(_7243_)
);

NOR2X1 _17525_ (
    .A(_6821_),
    .B(_7243_),
    .Y(_7244_)
);

NOR2X1 _17526_ (
    .A(_7237_),
    .B(_7238_),
    .Y(_7245_)
);

OAI21X1 _17527_ (
    .A(_7245_),
    .B(_7244_),
    .C(_7235_),
    .Y(_7246_)
);

AOI21X1 _17528_ (
    .A(_7242_),
    .B(_7246_),
    .C(_7234_),
    .Y(_7247_)
);

AOI21X1 _17529_ (
    .A(_6828_),
    .B(_6830_),
    .C(_6822_),
    .Y(_7248_)
);

OAI21X1 _17530_ (
    .A(_2792_),
    .B(_6050__bF$buf1),
    .C(_7238_),
    .Y(_7249_)
);

OAI21X1 _17531_ (
    .A(_2562__bF$buf2),
    .B(_5668__bF$buf1),
    .C(_7237_),
    .Y(_7251_)
);

AOI21X1 _17532_ (
    .A(_7249_),
    .B(_7251_),
    .C(_7235_),
    .Y(_7252_)
);

AOI21X1 _17533_ (
    .A(_7241_),
    .B(_7240_),
    .C(_7236_),
    .Y(_7253_)
);

NOR3X1 _17534_ (
    .A(_7253_),
    .B(_7248_),
    .C(_7252_),
    .Y(_7254_)
);

OAI21X1 _17535_ (
    .A(_7254_),
    .B(_7247_),
    .C(_7233_),
    .Y(_7255_)
);

OAI21X1 _17536_ (
    .A(_7252_),
    .B(_7253_),
    .C(_7248_),
    .Y(_7256_)
);

NAND3X1 _17537_ (
    .A(_7242_),
    .B(_7234_),
    .C(_7246_),
    .Y(_7257_)
);

NAND3X1 _17538_ (
    .A(_7232_),
    .B(_7256_),
    .C(_7257_),
    .Y(_7258_)
);

AOI21X1 _17539_ (
    .A(_7255_),
    .B(_7258_),
    .C(_7231_),
    .Y(_7259_)
);

OAI21X1 _17540_ (
    .A(_6827_),
    .B(_6831_),
    .C(_6819_),
    .Y(_7260_)
);

AOI21X1 _17541_ (
    .A(_6816_),
    .B(_7260_),
    .C(_6832_),
    .Y(_7262_)
);

AOI21X1 _17542_ (
    .A(_7256_),
    .B(_7257_),
    .C(_7232_),
    .Y(_7263_)
);

NOR3X1 _17543_ (
    .A(_7247_),
    .B(_7233_),
    .C(_7254_),
    .Y(_7264_)
);

NOR3X1 _17544_ (
    .A(_7262_),
    .B(_7263_),
    .C(_7264_),
    .Y(_7265_)
);

OAI21X1 _17545_ (
    .A(_7259_),
    .B(_7265_),
    .C(_7227_),
    .Y(_7266_)
);

OAI21X1 _17546_ (
    .A(_7264_),
    .B(_7263_),
    .C(_7262_),
    .Y(_7267_)
);

NAND3X1 _17547_ (
    .A(_7255_),
    .B(_7258_),
    .C(_7231_),
    .Y(_7268_)
);

NAND3X1 _17548_ (
    .A(_7226_),
    .B(_7267_),
    .C(_7268_),
    .Y(_7269_)
);

AND2X2 _17549_ (
    .A(_7266_),
    .B(_7269_),
    .Y(_7270_)
);

AOI21X1 _17550_ (
    .A(_6874_),
    .B(_6879_),
    .C(_6881_),
    .Y(_7271_)
);

OAI21X1 _17551_ (
    .A(_6890_),
    .B(_7271_),
    .C(_6882_),
    .Y(_7273_)
);

NAND2X1 _17552_ (
    .A(_6866_),
    .B(_6874_),
    .Y(_7274_)
);

OAI21X1 _17553_ (
    .A(_6861_),
    .B(_6851_),
    .C(_6855_),
    .Y(_7275_)
);

NAND2X1 _17554_ (
    .A(areg_5_bF$buf0),
    .B(breg_26_bF$buf4),
    .Y(_7276_)
);

AOI22X1 _17555_ (
    .A(areg_6_bF$buf1),
    .B(breg_25_bF$buf0),
    .C(areg_7_bF$buf2),
    .D(breg_24_bF$buf1),
    .Y(_7277_)
);

NAND2X1 _17556_ (
    .A(areg_7_bF$buf1),
    .B(breg_25_bF$buf5),
    .Y(_7278_)
);

NOR2X1 _17557_ (
    .A(_6857_),
    .B(_7278_),
    .Y(_7279_)
);

OAI21X1 _17558_ (
    .A(_7279_),
    .B(_7277_),
    .C(_7276_),
    .Y(_7280_)
);

INVX1 _17559_ (
    .A(_7276_),
    .Y(_7281_)
);

INVX1 _17560_ (
    .A(_7277_),
    .Y(_7282_)
);

OR2X2 _17561_ (
    .A(_6857_),
    .B(_7278_),
    .Y(_7284_)
);

NAND3X1 _17562_ (
    .A(_7281_),
    .B(_7282_),
    .C(_7284_),
    .Y(_7285_)
);

NAND2X1 _17563_ (
    .A(areg_9_bF$buf1),
    .B(breg_22_bF$buf0),
    .Y(_7286_)
);

OAI22X1 _17564_ (
    .A(_6514_),
    .B(_7286_),
    .C(_6929_),
    .D(_6925_),
    .Y(_7287_)
);

NAND3X1 _17565_ (
    .A(_7280_),
    .B(_7285_),
    .C(_7287_),
    .Y(_7288_)
);

AOI21X1 _17566_ (
    .A(_7282_),
    .B(_7284_),
    .C(_7281_),
    .Y(_7289_)
);

NOR3X1 _17567_ (
    .A(_7276_),
    .B(_7277_),
    .C(_7279_),
    .Y(_7290_)
);

OAI21X1 _17568_ (
    .A(_6582__bF$buf2),
    .B(_3781__bF$buf0),
    .C(_6863_),
    .Y(_7291_)
);

AOI21X1 _17569_ (
    .A(_6926_),
    .B(_7291_),
    .C(_6928_),
    .Y(_7292_)
);

OAI21X1 _17570_ (
    .A(_7289_),
    .B(_7290_),
    .C(_7292_),
    .Y(_7293_)
);

NAND3X1 _17571_ (
    .A(_7275_),
    .B(_7288_),
    .C(_7293_),
    .Y(_7295_)
);

INVX1 _17572_ (
    .A(_7275_),
    .Y(_7296_)
);

NAND3X1 _17573_ (
    .A(_7292_),
    .B(_7280_),
    .C(_7285_),
    .Y(_7297_)
);

OAI21X1 _17574_ (
    .A(_7289_),
    .B(_7290_),
    .C(_7287_),
    .Y(_7298_)
);

NAND3X1 _17575_ (
    .A(_7296_),
    .B(_7297_),
    .C(_7298_),
    .Y(_7299_)
);

AOI21X1 _17576_ (
    .A(_6948_),
    .B(_6949_),
    .C(_6932_),
    .Y(_7300_)
);

OAI21X1 _17577_ (
    .A(_6931_),
    .B(_7300_),
    .C(_6953_),
    .Y(_7301_)
);

NAND3X1 _17578_ (
    .A(_7295_),
    .B(_7299_),
    .C(_7301_),
    .Y(_7302_)
);

AOI21X1 _17579_ (
    .A(_7297_),
    .B(_7298_),
    .C(_7296_),
    .Y(_7303_)
);

AOI21X1 _17580_ (
    .A(_7288_),
    .B(_7293_),
    .C(_7275_),
    .Y(_7304_)
);

NOR3X1 _17581_ (
    .A(_6947_),
    .B(_6945_),
    .C(_6940_),
    .Y(_7306_)
);

AOI21X1 _17582_ (
    .A(_6954_),
    .B(_6952_),
    .C(_7306_),
    .Y(_7307_)
);

OAI21X1 _17583_ (
    .A(_7303_),
    .B(_7304_),
    .C(_7307_),
    .Y(_7308_)
);

NAND3X1 _17584_ (
    .A(_7274_),
    .B(_7308_),
    .C(_7302_),
    .Y(_7309_)
);

AND2X2 _17585_ (
    .A(_6874_),
    .B(_6866_),
    .Y(_7310_)
);

NAND3X1 _17586_ (
    .A(_7295_),
    .B(_7299_),
    .C(_7307_),
    .Y(_7311_)
);

OAI21X1 _17587_ (
    .A(_7303_),
    .B(_7304_),
    .C(_7301_),
    .Y(_7312_)
);

NAND3X1 _17588_ (
    .A(_7310_),
    .B(_7312_),
    .C(_7311_),
    .Y(_7313_)
);

NAND3X1 _17589_ (
    .A(_7309_),
    .B(_7313_),
    .C(_7273_),
    .Y(_7314_)
);

NOR3X1 _17590_ (
    .A(_6886_),
    .B(_6883_),
    .C(_6884_),
    .Y(_7315_)
);

AOI21X1 _17591_ (
    .A(_6848_),
    .B(_6887_),
    .C(_7315_),
    .Y(_7317_)
);

AOI21X1 _17592_ (
    .A(_7312_),
    .B(_7311_),
    .C(_7310_),
    .Y(_7318_)
);

AOI21X1 _17593_ (
    .A(_7308_),
    .B(_7302_),
    .C(_7274_),
    .Y(_7319_)
);

OAI21X1 _17594_ (
    .A(_7318_),
    .B(_7319_),
    .C(_7317_),
    .Y(_7320_)
);

NAND3X1 _17595_ (
    .A(_7314_),
    .B(_7320_),
    .C(_7270_),
    .Y(_7321_)
);

NAND2X1 _17596_ (
    .A(_7269_),
    .B(_7266_),
    .Y(_7322_)
);

OAI21X1 _17597_ (
    .A(_7318_),
    .B(_7319_),
    .C(_7273_),
    .Y(_7323_)
);

NAND3X1 _17598_ (
    .A(_7309_),
    .B(_7313_),
    .C(_7317_),
    .Y(_7324_)
);

NAND3X1 _17599_ (
    .A(_7322_),
    .B(_7324_),
    .C(_7323_),
    .Y(_7325_)
);

AOI21X1 _17600_ (
    .A(_6997_),
    .B(_7002_),
    .C(_7003_),
    .Y(_7326_)
);

OAI21X1 _17601_ (
    .A(_7326_),
    .B(_6924_),
    .C(_7004_),
    .Y(_7328_)
);

NAND3X1 _17602_ (
    .A(_7325_),
    .B(_7328_),
    .C(_7321_),
    .Y(_7329_)
);

AOI21X1 _17603_ (
    .A(_7324_),
    .B(_7323_),
    .C(_7322_),
    .Y(_7330_)
);

AOI21X1 _17604_ (
    .A(_7314_),
    .B(_7320_),
    .C(_7270_),
    .Y(_7331_)
);

NOR3X1 _17605_ (
    .A(_7006_),
    .B(_7007_),
    .C(_7005_),
    .Y(_7332_)
);

AOI21X1 _17606_ (
    .A(_6923_),
    .B(_7008_),
    .C(_7332_),
    .Y(_7333_)
);

OAI21X1 _17607_ (
    .A(_7331_),
    .B(_7330_),
    .C(_7333_),
    .Y(_7334_)
);

NAND3X1 _17608_ (
    .A(_7224_),
    .B(_7329_),
    .C(_7334_),
    .Y(_7335_)
);

NAND2X1 _17609_ (
    .A(_6894_),
    .B(_6902_),
    .Y(_7336_)
);

NAND3X1 _17610_ (
    .A(_7325_),
    .B(_7321_),
    .C(_7333_),
    .Y(_7337_)
);

OAI21X1 _17611_ (
    .A(_7331_),
    .B(_7330_),
    .C(_7328_),
    .Y(_7339_)
);

NAND3X1 _17612_ (
    .A(_7336_),
    .B(_7339_),
    .C(_7337_),
    .Y(_7340_)
);

NAND2X1 _17613_ (
    .A(_7335_),
    .B(_7340_),
    .Y(_7341_)
);

AOI21X1 _17614_ (
    .A(_7156_),
    .B(_7162_),
    .C(_7015_),
    .Y(_7342_)
);

OAI21X1 _17615_ (
    .A(_7173_),
    .B(_7342_),
    .C(_7163_),
    .Y(_7343_)
);

AND2X2 _17616_ (
    .A(_6997_),
    .B(_6990_),
    .Y(_7344_)
);

NOR2X1 _17617_ (
    .A(_5190__bF$buf1),
    .B(_5369_),
    .Y(_7345_)
);

NAND2X1 _17618_ (
    .A(areg_10_bF$buf1),
    .B(breg_21_bF$buf0),
    .Y(_7346_)
);

NOR2X1 _17619_ (
    .A(_7286_),
    .B(_7346_),
    .Y(_7347_)
);

AND2X2 _17620_ (
    .A(_7286_),
    .B(_7346_),
    .Y(_7348_)
);

NOR2X1 _17621_ (
    .A(_7347_),
    .B(_7348_),
    .Y(_7350_)
);

XNOR2X1 _17622_ (
    .A(_7350_),
    .B(_7345_),
    .Y(_7351_)
);

OAI21X1 _17623_ (
    .A(_6939_),
    .B(_6934_),
    .C(_6942_),
    .Y(_7352_)
);

NAND2X1 _17624_ (
    .A(areg_11_bF$buf1),
    .B(breg_20_bF$buf0),
    .Y(_7353_)
);

NAND2X1 _17625_ (
    .A(areg_12_bF$buf2),
    .B(breg_19_bF$buf2),
    .Y(_7354_)
);

NAND2X1 _17626_ (
    .A(areg_13_bF$buf0),
    .B(breg_18_bF$buf1),
    .Y(_7355_)
);

NOR2X1 _17627_ (
    .A(_7354_),
    .B(_7355_),
    .Y(_7356_)
);

AND2X2 _17628_ (
    .A(areg_12_bF$buf1),
    .B(breg_19_bF$buf1),
    .Y(_7357_)
);

AND2X2 _17629_ (
    .A(areg_13_bF$buf4),
    .B(breg_18_bF$buf0),
    .Y(_7358_)
);

NOR2X1 _17630_ (
    .A(_7357_),
    .B(_7358_),
    .Y(_7359_)
);

NOR3X1 _17631_ (
    .A(_7353_),
    .B(_7356_),
    .C(_7359_),
    .Y(_7361_)
);

INVX2 _17632_ (
    .A(_7353_),
    .Y(_7362_)
);

NAND2X1 _17633_ (
    .A(_7357_),
    .B(_7358_),
    .Y(_7363_)
);

OAI21X1 _17634_ (
    .A(_549__bF$buf4),
    .B(_3529__bF$buf2),
    .C(_7354_),
    .Y(_7364_)
);

AOI21X1 _17635_ (
    .A(_7364_),
    .B(_7363_),
    .C(_7362_),
    .Y(_7365_)
);

OAI21X1 _17636_ (
    .A(_7361_),
    .B(_7365_),
    .C(_7352_),
    .Y(_7366_)
);

AOI21X1 _17637_ (
    .A(_6941_),
    .B(_6943_),
    .C(_6936_),
    .Y(_7367_)
);

NAND3X1 _17638_ (
    .A(_7362_),
    .B(_7364_),
    .C(_7363_),
    .Y(_7368_)
);

OAI21X1 _17639_ (
    .A(_7359_),
    .B(_7356_),
    .C(_7353_),
    .Y(_7369_)
);

NAND3X1 _17640_ (
    .A(_7367_),
    .B(_7368_),
    .C(_7369_),
    .Y(_7370_)
);

AOI21X1 _17641_ (
    .A(_7366_),
    .B(_7370_),
    .C(_7351_),
    .Y(_7372_)
);

INVX2 _17642_ (
    .A(_7345_),
    .Y(_7373_)
);

XNOR2X1 _17643_ (
    .A(_7350_),
    .B(_7373_),
    .Y(_7374_)
);

NAND3X1 _17644_ (
    .A(_7368_),
    .B(_7352_),
    .C(_7369_),
    .Y(_7375_)
);

OAI21X1 _17645_ (
    .A(_7361_),
    .B(_7365_),
    .C(_7367_),
    .Y(_7376_)
);

AOI21X1 _17646_ (
    .A(_7376_),
    .B(_7375_),
    .C(_7374_),
    .Y(_7377_)
);

NOR2X1 _17647_ (
    .A(_7372_),
    .B(_7377_),
    .Y(_7378_)
);

OAI21X1 _17648_ (
    .A(_6985_),
    .B(_6987_),
    .C(_6978_),
    .Y(_7379_)
);

OAI21X1 _17649_ (
    .A(_6972_),
    .B(_6961_),
    .C(_6965_),
    .Y(_7380_)
);

NAND2X1 _17650_ (
    .A(areg_14_bF$buf4),
    .B(breg_17_bF$buf4),
    .Y(_7381_)
);

INVX1 _17651_ (
    .A(_7381_),
    .Y(_7383_)
);

AND2X2 _17652_ (
    .A(areg_15_bF$buf3),
    .B(breg_16_bF$buf1),
    .Y(_7384_)
);

AND2X2 _17653_ (
    .A(breg_15_bF$buf5),
    .B(areg_16_bF$buf0),
    .Y(_7385_)
);

NAND2X1 _17654_ (
    .A(_7384_),
    .B(_7385_),
    .Y(_7386_)
);

OAI22X1 _17655_ (
    .A(_2465__bF$buf1),
    .B(_2560__bF$buf2),
    .C(_2362__bF$buf0),
    .D(_2669__bF$buf2),
    .Y(_7387_)
);

NAND3X1 _17656_ (
    .A(_7383_),
    .B(_7387_),
    .C(_7386_),
    .Y(_7388_)
);

OAI21X1 _17657_ (
    .A(_2465__bF$buf0),
    .B(_2560__bF$buf1),
    .C(_7385_),
    .Y(_7389_)
);

OAI21X1 _17658_ (
    .A(_2362__bF$buf5),
    .B(_2669__bF$buf1),
    .C(_7384_),
    .Y(_7390_)
);

NAND3X1 _17659_ (
    .A(_7381_),
    .B(_7389_),
    .C(_7390_),
    .Y(_7391_)
);

NAND2X1 _17660_ (
    .A(breg_13_bF$buf1),
    .B(areg_18_bF$buf0),
    .Y(_7392_)
);

OAI22X1 _17661_ (
    .A(_6974_),
    .B(_7392_),
    .C(_7021_),
    .D(_7017_),
    .Y(_7394_)
);

NAND3X1 _17662_ (
    .A(_7388_),
    .B(_7391_),
    .C(_7394_),
    .Y(_7395_)
);

AOI21X1 _17663_ (
    .A(_7389_),
    .B(_7390_),
    .C(_7381_),
    .Y(_7396_)
);

AOI21X1 _17664_ (
    .A(_7387_),
    .B(_7386_),
    .C(_7383_),
    .Y(_7397_)
);

OAI21X1 _17665_ (
    .A(_2586__bF$buf0),
    .B(_3146__bF$buf1),
    .C(_6606_),
    .Y(_7398_)
);

AOI21X1 _17666_ (
    .A(_7045_),
    .B(_7398_),
    .C(_7019_),
    .Y(_7399_)
);

OAI21X1 _17667_ (
    .A(_7396_),
    .B(_7397_),
    .C(_7399_),
    .Y(_7400_)
);

NAND3X1 _17668_ (
    .A(_7380_),
    .B(_7395_),
    .C(_7400_),
    .Y(_7401_)
);

INVX2 _17669_ (
    .A(_7380_),
    .Y(_7402_)
);

NOR3X1 _17670_ (
    .A(_7397_),
    .B(_7399_),
    .C(_7396_),
    .Y(_7403_)
);

AOI21X1 _17671_ (
    .A(_7388_),
    .B(_7391_),
    .C(_7394_),
    .Y(_7405_)
);

OAI21X1 _17672_ (
    .A(_7403_),
    .B(_7405_),
    .C(_7402_),
    .Y(_7406_)
);

NAND3X1 _17673_ (
    .A(_7401_),
    .B(_7406_),
    .C(_7379_),
    .Y(_7407_)
);

AOI21X1 _17674_ (
    .A(_6960_),
    .B(_6983_),
    .C(_6986_),
    .Y(_7408_)
);

NAND3X1 _17675_ (
    .A(_7399_),
    .B(_7388_),
    .C(_7391_),
    .Y(_7409_)
);

OAI21X1 _17676_ (
    .A(_7396_),
    .B(_7397_),
    .C(_7394_),
    .Y(_7410_)
);

AOI21X1 _17677_ (
    .A(_7409_),
    .B(_7410_),
    .C(_7402_),
    .Y(_7411_)
);

AOI21X1 _17678_ (
    .A(_7395_),
    .B(_7400_),
    .C(_7380_),
    .Y(_7412_)
);

OAI21X1 _17679_ (
    .A(_7412_),
    .B(_7411_),
    .C(_7408_),
    .Y(_7413_)
);

NAND3X1 _17680_ (
    .A(_7413_),
    .B(_7378_),
    .C(_7407_),
    .Y(_7414_)
);

OR2X2 _17681_ (
    .A(_7372_),
    .B(_7377_),
    .Y(_7416_)
);

OAI21X1 _17682_ (
    .A(_7412_),
    .B(_7411_),
    .C(_7379_),
    .Y(_7417_)
);

NAND3X1 _17683_ (
    .A(_7401_),
    .B(_7406_),
    .C(_7408_),
    .Y(_7418_)
);

NAND3X1 _17684_ (
    .A(_7417_),
    .B(_7418_),
    .C(_7416_),
    .Y(_7419_)
);

AOI21X1 _17685_ (
    .A(_7044_),
    .B(_7049_),
    .C(_7050_),
    .Y(_7420_)
);

OAI21X1 _17686_ (
    .A(_7420_),
    .B(_7016_),
    .C(_7051_),
    .Y(_7421_)
);

NAND3X1 _17687_ (
    .A(_7414_),
    .B(_7421_),
    .C(_7419_),
    .Y(_7422_)
);

AOI21X1 _17688_ (
    .A(_7417_),
    .B(_7418_),
    .C(_7416_),
    .Y(_7423_)
);

AOI21X1 _17689_ (
    .A(_7413_),
    .B(_7407_),
    .C(_7378_),
    .Y(_7424_)
);

NOR3X1 _17690_ (
    .A(_7053_),
    .B(_7055_),
    .C(_7052_),
    .Y(_7425_)
);

AOI21X1 _17691_ (
    .A(_7058_),
    .B(_7056_),
    .C(_7425_),
    .Y(_7427_)
);

OAI21X1 _17692_ (
    .A(_7423_),
    .B(_7424_),
    .C(_7427_),
    .Y(_7428_)
);

NAND3X1 _17693_ (
    .A(_7422_),
    .B(_7344_),
    .C(_7428_),
    .Y(_7429_)
);

NAND2X1 _17694_ (
    .A(_6990_),
    .B(_6997_),
    .Y(_7430_)
);

NAND3X1 _17695_ (
    .A(_7414_),
    .B(_7419_),
    .C(_7427_),
    .Y(_7431_)
);

OAI21X1 _17696_ (
    .A(_7423_),
    .B(_7424_),
    .C(_7421_),
    .Y(_7432_)
);

NAND3X1 _17697_ (
    .A(_7430_),
    .B(_7432_),
    .C(_7431_),
    .Y(_7433_)
);

NAND2X1 _17698_ (
    .A(_7433_),
    .B(_7429_),
    .Y(_7434_)
);

AOI21X1 _17699_ (
    .A(_7141_),
    .B(_7148_),
    .C(_7064_),
    .Y(_7435_)
);

OAI21X1 _17700_ (
    .A(_7159_),
    .B(_7435_),
    .C(_7149_),
    .Y(_7436_)
);

AND2X2 _17701_ (
    .A(_7044_),
    .B(_7038_),
    .Y(_7438_)
);

NAND2X1 _17702_ (
    .A(breg_14_bF$buf0),
    .B(areg_17_bF$buf5),
    .Y(_7439_)
);

NAND2X1 _17703_ (
    .A(breg_12_bF$buf4),
    .B(areg_19_bF$buf1),
    .Y(_7440_)
);

XOR2X1 _17704_ (
    .A(_7392_),
    .B(_7440_),
    .Y(_7441_)
);

XNOR2X1 _17705_ (
    .A(_7441_),
    .B(_7439_),
    .Y(_7442_)
);

OAI21X1 _17706_ (
    .A(_7036_),
    .B(_7025_),
    .C(_7029_),
    .Y(_7443_)
);

NAND2X1 _17707_ (
    .A(breg_11_bF$buf1),
    .B(areg_20_bF$buf4),
    .Y(_7444_)
);

INVX2 _17708_ (
    .A(_7444_),
    .Y(_7445_)
);

AND2X2 _17709_ (
    .A(breg_10_bF$buf1),
    .B(areg_21_bF$buf1),
    .Y(_7446_)
);

AND2X2 _17710_ (
    .A(breg_9_bF$buf4),
    .B(areg_22_bF$buf2),
    .Y(_7447_)
);

NAND2X1 _17711_ (
    .A(_7446_),
    .B(_7447_),
    .Y(_7449_)
);

OAI22X1 _17712_ (
    .A(_6044__bF$buf2),
    .B(_4551__bF$buf4),
    .C(_7217__bF$buf0),
    .D(_3961__bF$buf1),
    .Y(_7450_)
);

NAND3X1 _17713_ (
    .A(_7445_),
    .B(_7450_),
    .C(_7449_),
    .Y(_7451_)
);

NAND2X1 _17714_ (
    .A(breg_10_bF$buf0),
    .B(areg_22_bF$buf1),
    .Y(_7452_)
);

NOR2X1 _17715_ (
    .A(_7034_),
    .B(_7452_),
    .Y(_7453_)
);

NOR2X1 _17716_ (
    .A(_7446_),
    .B(_7447_),
    .Y(_7454_)
);

OAI21X1 _17717_ (
    .A(_7454_),
    .B(_7453_),
    .C(_7444_),
    .Y(_7455_)
);

NAND3X1 _17718_ (
    .A(_7451_),
    .B(_7443_),
    .C(_7455_),
    .Y(_7456_)
);

AOI21X1 _17719_ (
    .A(_7026_),
    .B(_7030_),
    .C(_7035_),
    .Y(_7457_)
);

OAI21X1 _17720_ (
    .A(_7217__bF$buf4),
    .B(_3961__bF$buf0),
    .C(_7447_),
    .Y(_7458_)
);

OAI21X1 _17721_ (
    .A(_6044__bF$buf1),
    .B(_4551__bF$buf3),
    .C(_7446_),
    .Y(_7460_)
);

AOI21X1 _17722_ (
    .A(_7458_),
    .B(_7460_),
    .C(_7444_),
    .Y(_7461_)
);

AOI21X1 _17723_ (
    .A(_7450_),
    .B(_7449_),
    .C(_7445_),
    .Y(_7462_)
);

OAI21X1 _17724_ (
    .A(_7461_),
    .B(_7462_),
    .C(_7457_),
    .Y(_7463_)
);

NAND3X1 _17725_ (
    .A(_7456_),
    .B(_7463_),
    .C(_7442_),
    .Y(_7464_)
);

INVX2 _17726_ (
    .A(_7439_),
    .Y(_7465_)
);

XNOR2X1 _17727_ (
    .A(_7441_),
    .B(_7465_),
    .Y(_7466_)
);

OAI21X1 _17728_ (
    .A(_7461_),
    .B(_7462_),
    .C(_7443_),
    .Y(_7467_)
);

NAND3X1 _17729_ (
    .A(_7457_),
    .B(_7451_),
    .C(_7455_),
    .Y(_7468_)
);

NAND3X1 _17730_ (
    .A(_7467_),
    .B(_7468_),
    .C(_7466_),
    .Y(_7469_)
);

OAI21X1 _17731_ (
    .A(_7089_),
    .B(_7066_),
    .C(_7079_),
    .Y(_7471_)
);

NAND3X1 _17732_ (
    .A(_7471_),
    .B(_7464_),
    .C(_7469_),
    .Y(_7472_)
);

AOI21X1 _17733_ (
    .A(_7467_),
    .B(_7468_),
    .C(_7466_),
    .Y(_7473_)
);

AOI21X1 _17734_ (
    .A(_7456_),
    .B(_7463_),
    .C(_7442_),
    .Y(_7474_)
);

AOI21X1 _17735_ (
    .A(_7086_),
    .B(_7083_),
    .C(_7088_),
    .Y(_7475_)
);

OAI21X1 _17736_ (
    .A(_7473_),
    .B(_7474_),
    .C(_7475_),
    .Y(_7476_)
);

NAND3X1 _17737_ (
    .A(_7472_),
    .B(_7476_),
    .C(_7438_),
    .Y(_7477_)
);

NAND2X1 _17738_ (
    .A(_7038_),
    .B(_7044_),
    .Y(_7478_)
);

NOR3X1 _17739_ (
    .A(_7474_),
    .B(_7475_),
    .C(_7473_),
    .Y(_7479_)
);

AOI21X1 _17740_ (
    .A(_7464_),
    .B(_7469_),
    .C(_7471_),
    .Y(_7480_)
);

OAI21X1 _17741_ (
    .A(_7479_),
    .B(_7480_),
    .C(_7478_),
    .Y(_7482_)
);

NAND2X1 _17742_ (
    .A(_7477_),
    .B(_7482_),
    .Y(_7483_)
);

AOI21X1 _17743_ (
    .A(_7134_),
    .B(_7129_),
    .C(_7093_),
    .Y(_7484_)
);

OAI21X1 _17744_ (
    .A(_7145_),
    .B(_7484_),
    .C(_7135_),
    .Y(_7485_)
);

AND2X2 _17745_ (
    .A(breg_7_bF$buf3),
    .B(areg_24_bF$buf4),
    .Y(_7486_)
);

AOI21X1 _17746_ (
    .A(_6655_),
    .B(_7486_),
    .C(_7080_),
    .Y(_7487_)
);

NAND2X1 _17747_ (
    .A(breg[8]),
    .B(areg_23_bF$buf4),
    .Y(_7488_)
);

INVX1 _17748_ (
    .A(_7488_),
    .Y(_7489_)
);

AND2X2 _17749_ (
    .A(breg_6_bF$buf2),
    .B(areg_25_bF$buf0),
    .Y(_7490_)
);

NAND2X1 _17750_ (
    .A(_7486_),
    .B(_7490_),
    .Y(_7491_)
);

NAND2X1 _17751_ (
    .A(breg_7_bF$buf2),
    .B(areg_24_bF$buf3),
    .Y(_7493_)
);

OAI21X1 _17752_ (
    .A(_5453__bF$buf1),
    .B(_6300__bF$buf2),
    .C(_7493_),
    .Y(_7494_)
);

NAND3X1 _17753_ (
    .A(_7489_),
    .B(_7494_),
    .C(_7491_),
    .Y(_7495_)
);

OAI21X1 _17754_ (
    .A(_4116__bF$buf3),
    .B(_5921__bF$buf0),
    .C(_7490_),
    .Y(_7496_)
);

OAI21X1 _17755_ (
    .A(_5453__bF$buf0),
    .B(_6300__bF$buf1),
    .C(_7486_),
    .Y(_7497_)
);

NAND3X1 _17756_ (
    .A(_7488_),
    .B(_7496_),
    .C(_7497_),
    .Y(_7498_)
);

OAI21X1 _17757_ (
    .A(_7104_),
    .B(_7094_),
    .C(_7099_),
    .Y(_7499_)
);

NAND3X1 _17758_ (
    .A(_7495_),
    .B(_7498_),
    .C(_7499_),
    .Y(_7500_)
);

AOI21X1 _17759_ (
    .A(_7496_),
    .B(_7497_),
    .C(_7488_),
    .Y(_7501_)
);

AOI21X1 _17760_ (
    .A(_7494_),
    .B(_7491_),
    .C(_7489_),
    .Y(_7502_)
);

AOI21X1 _17761_ (
    .A(_7095_),
    .B(_7101_),
    .C(_7103_),
    .Y(_7504_)
);

OAI21X1 _17762_ (
    .A(_7501_),
    .B(_7502_),
    .C(_7504_),
    .Y(_7505_)
);

NAND3X1 _17763_ (
    .A(_7487_),
    .B(_7500_),
    .C(_7505_),
    .Y(_7506_)
);

OAI21X1 _17764_ (
    .A(_7085_),
    .B(_7493_),
    .C(_7073_),
    .Y(_7507_)
);

NOR3X1 _17765_ (
    .A(_7502_),
    .B(_7504_),
    .C(_7501_),
    .Y(_7508_)
);

AOI21X1 _17766_ (
    .A(_7495_),
    .B(_7498_),
    .C(_7499_),
    .Y(_7509_)
);

OAI21X1 _17767_ (
    .A(_7508_),
    .B(_7509_),
    .C(_7507_),
    .Y(_7510_)
);

NAND2X1 _17768_ (
    .A(_7506_),
    .B(_7510_),
    .Y(_7511_)
);

AOI21X1 _17769_ (
    .A(_7118_),
    .B(_7115_),
    .C(_7107_),
    .Y(_7512_)
);

OAI21X1 _17770_ (
    .A(_7512_),
    .B(_7130_),
    .C(_7119_),
    .Y(_7513_)
);

NAND2X1 _17771_ (
    .A(breg_5_bF$buf2),
    .B(areg_26_bF$buf1),
    .Y(_7515_)
);

INVX1 _17772_ (
    .A(_7515_),
    .Y(_7516_)
);

NAND2X1 _17773_ (
    .A(breg_4_bF$buf1),
    .B(areg_27_bF$buf2),
    .Y(_7517_)
);

NAND2X1 _17774_ (
    .A(breg_3_bF$buf3),
    .B(areg_28_bF$buf4),
    .Y(_7518_)
);

OR2X2 _17775_ (
    .A(_7517_),
    .B(_7518_),
    .Y(_7519_)
);

INVX8 _17776_ (
    .A(areg_28_bF$buf3),
    .Y(_7520_)
);

OAI21X1 _17777_ (
    .A(_2365_),
    .B(_7520__bF$buf3),
    .C(_7517_),
    .Y(_7521_)
);

NAND3X1 _17778_ (
    .A(_7516_),
    .B(_7521_),
    .C(_7519_),
    .Y(_7522_)
);

NOR2X1 _17779_ (
    .A(_7517_),
    .B(_7518_),
    .Y(_7523_)
);

AND2X2 _17780_ (
    .A(_7517_),
    .B(_7518_),
    .Y(_7524_)
);

OAI21X1 _17781_ (
    .A(_7524_),
    .B(_7523_),
    .C(_7515_),
    .Y(_7526_)
);

AND2X2 _17782_ (
    .A(_7522_),
    .B(_7526_),
    .Y(_7527_)
);

OAI21X1 _17783_ (
    .A(_7108_),
    .B(_7113_),
    .C(_7112_),
    .Y(_7528_)
);

NAND2X1 _17784_ (
    .A(breg_2_bF$buf2),
    .B(areg_29_bF$buf4),
    .Y(_7529_)
);

INVX1 _17785_ (
    .A(_7529_),
    .Y(_7530_)
);

AND2X2 _17786_ (
    .A(breg_0_bF$buf1),
    .B(areg_31_bF$buf4),
    .Y(_7531_)
);

NAND2X1 _17787_ (
    .A(_7111_),
    .B(_7531_),
    .Y(_7532_)
);

AOI22X1 _17788_ (
    .A(breg_0_bF$buf0),
    .B(areg_31_bF$buf3),
    .C(breg_1_bF$buf1),
    .D(areg_30_bF$buf0),
    .Y(_7533_)
);

INVX1 _17789_ (
    .A(_7533_),
    .Y(_7534_)
);

NAND3X1 _17790_ (
    .A(_7530_),
    .B(_7534_),
    .C(_7532_),
    .Y(_7535_)
);

NAND3X1 _17791_ (
    .A(breg_0_bF$buf6),
    .B(areg_31_bF$buf2),
    .C(_7116_),
    .Y(_7537_)
);

NAND2X1 _17792_ (
    .A(breg_0_bF$buf5),
    .B(areg_31_bF$buf1),
    .Y(_7538_)
);

NAND2X1 _17793_ (
    .A(_7538_),
    .B(_7111_),
    .Y(_7539_)
);

NAND3X1 _17794_ (
    .A(_7529_),
    .B(_7537_),
    .C(_7539_),
    .Y(_7540_)
);

NAND3X1 _17795_ (
    .A(_7528_),
    .B(_7540_),
    .C(_7535_),
    .Y(_7541_)
);

AOI21X1 _17796_ (
    .A(_7110_),
    .B(_7114_),
    .C(_7117_),
    .Y(_7542_)
);

AOI21X1 _17797_ (
    .A(_7537_),
    .B(_7539_),
    .C(_7529_),
    .Y(_7543_)
);

AOI21X1 _17798_ (
    .A(_7534_),
    .B(_7532_),
    .C(_7530_),
    .Y(_7544_)
);

OAI21X1 _17799_ (
    .A(_7544_),
    .B(_7543_),
    .C(_7542_),
    .Y(_7545_)
);

NAND3X1 _17800_ (
    .A(_7541_),
    .B(_7545_),
    .C(_7527_),
    .Y(_7546_)
);

NAND2X1 _17801_ (
    .A(_7526_),
    .B(_7522_),
    .Y(_7548_)
);

OAI21X1 _17802_ (
    .A(_7544_),
    .B(_7543_),
    .C(_7528_),
    .Y(_7549_)
);

NAND3X1 _17803_ (
    .A(_7540_),
    .B(_7542_),
    .C(_7535_),
    .Y(_7550_)
);

NAND3X1 _17804_ (
    .A(_7548_),
    .B(_7550_),
    .C(_7549_),
    .Y(_7551_)
);

NAND3X1 _17805_ (
    .A(_7513_),
    .B(_7551_),
    .C(_7546_),
    .Y(_7552_)
);

NOR3X1 _17806_ (
    .A(_7121_),
    .B(_7126_),
    .C(_7127_),
    .Y(_7553_)
);

AOI21X1 _17807_ (
    .A(_7128_),
    .B(_7106_),
    .C(_7553_),
    .Y(_7554_)
);

AOI21X1 _17808_ (
    .A(_7550_),
    .B(_7549_),
    .C(_7548_),
    .Y(_7555_)
);

AOI21X1 _17809_ (
    .A(_7541_),
    .B(_7545_),
    .C(_7527_),
    .Y(_7556_)
);

OAI21X1 _17810_ (
    .A(_7555_),
    .B(_7556_),
    .C(_7554_),
    .Y(_7557_)
);

NAND3X1 _17811_ (
    .A(_7552_),
    .B(_7511_),
    .C(_7557_),
    .Y(_7559_)
);

NAND3X1 _17812_ (
    .A(_7507_),
    .B(_7500_),
    .C(_7505_),
    .Y(_7560_)
);

OAI21X1 _17813_ (
    .A(_7508_),
    .B(_7509_),
    .C(_7487_),
    .Y(_7561_)
);

NAND2X1 _17814_ (
    .A(_7560_),
    .B(_7561_),
    .Y(_7562_)
);

OAI21X1 _17815_ (
    .A(_7555_),
    .B(_7556_),
    .C(_7513_),
    .Y(_7563_)
);

NAND3X1 _17816_ (
    .A(_7551_),
    .B(_7546_),
    .C(_7554_),
    .Y(_7564_)
);

NAND3X1 _17817_ (
    .A(_7564_),
    .B(_7562_),
    .C(_7563_),
    .Y(_7565_)
);

NAND3X1 _17818_ (
    .A(_7559_),
    .B(_7485_),
    .C(_7565_),
    .Y(_7566_)
);

NOR3X1 _17819_ (
    .A(_7138_),
    .B(_7139_),
    .C(_7137_),
    .Y(_7567_)
);

AOI21X1 _17820_ (
    .A(_7091_),
    .B(_7140_),
    .C(_7567_),
    .Y(_7568_)
);

AOI21X1 _17821_ (
    .A(_7564_),
    .B(_7563_),
    .C(_7562_),
    .Y(_7570_)
);

AOI21X1 _17822_ (
    .A(_7552_),
    .B(_7557_),
    .C(_7511_),
    .Y(_7571_)
);

OAI21X1 _17823_ (
    .A(_7570_),
    .B(_7571_),
    .C(_7568_),
    .Y(_7572_)
);

NAND3X1 _17824_ (
    .A(_7566_),
    .B(_7572_),
    .C(_7483_),
    .Y(_7573_)
);

NAND3X1 _17825_ (
    .A(_7478_),
    .B(_7472_),
    .C(_7476_),
    .Y(_7574_)
);

NAND3X1 _17826_ (
    .A(_7475_),
    .B(_7464_),
    .C(_7469_),
    .Y(_7575_)
);

OAI21X1 _17827_ (
    .A(_7473_),
    .B(_7474_),
    .C(_7471_),
    .Y(_7576_)
);

NAND3X1 _17828_ (
    .A(_7575_),
    .B(_7576_),
    .C(_7438_),
    .Y(_7577_)
);

NAND2X1 _17829_ (
    .A(_7574_),
    .B(_7577_),
    .Y(_7578_)
);

OAI21X1 _17830_ (
    .A(_7570_),
    .B(_7571_),
    .C(_7485_),
    .Y(_7579_)
);

NAND3X1 _17831_ (
    .A(_7559_),
    .B(_7565_),
    .C(_7568_),
    .Y(_7581_)
);

NAND3X1 _17832_ (
    .A(_7578_),
    .B(_7581_),
    .C(_7579_),
    .Y(_7582_)
);

NAND3X1 _17833_ (
    .A(_7582_),
    .B(_7436_),
    .C(_7573_),
    .Y(_7583_)
);

NOR3X1 _17834_ (
    .A(_7152_),
    .B(_7154_),
    .C(_7151_),
    .Y(_7584_)
);

AOI21X1 _17835_ (
    .A(_7062_),
    .B(_7155_),
    .C(_7584_),
    .Y(_7585_)
);

AOI21X1 _17836_ (
    .A(_7581_),
    .B(_7579_),
    .C(_7578_),
    .Y(_7586_)
);

AOI21X1 _17837_ (
    .A(_7566_),
    .B(_7572_),
    .C(_7483_),
    .Y(_7587_)
);

OAI21X1 _17838_ (
    .A(_7586_),
    .B(_7587_),
    .C(_7585_),
    .Y(_7588_)
);

NAND3X1 _17839_ (
    .A(_7583_),
    .B(_7434_),
    .C(_7588_),
    .Y(_7589_)
);

NAND3X1 _17840_ (
    .A(_7430_),
    .B(_7422_),
    .C(_7428_),
    .Y(_7590_)
);

NAND3X1 _17841_ (
    .A(_7432_),
    .B(_7344_),
    .C(_7431_),
    .Y(_7592_)
);

NAND2X1 _17842_ (
    .A(_7590_),
    .B(_7592_),
    .Y(_7593_)
);

OAI21X1 _17843_ (
    .A(_7586_),
    .B(_7587_),
    .C(_7436_),
    .Y(_7594_)
);

NAND3X1 _17844_ (
    .A(_7573_),
    .B(_7582_),
    .C(_7585_),
    .Y(_7595_)
);

NAND3X1 _17845_ (
    .A(_7593_),
    .B(_7595_),
    .C(_7594_),
    .Y(_7596_)
);

NAND3X1 _17846_ (
    .A(_7589_),
    .B(_7596_),
    .C(_7343_),
    .Y(_7597_)
);

NOR3X1 _17847_ (
    .A(_7167_),
    .B(_7168_),
    .C(_7166_),
    .Y(_7598_)
);

AOI21X1 _17848_ (
    .A(_7169_),
    .B(_7013_),
    .C(_7598_),
    .Y(_7599_)
);

AOI21X1 _17849_ (
    .A(_7595_),
    .B(_7594_),
    .C(_7593_),
    .Y(_7600_)
);

AOI21X1 _17850_ (
    .A(_7583_),
    .B(_7588_),
    .C(_7434_),
    .Y(_7601_)
);

OAI21X1 _17851_ (
    .A(_7600_),
    .B(_7601_),
    .C(_7599_),
    .Y(_7603_)
);

NAND3X1 _17852_ (
    .A(_7597_),
    .B(_7341_),
    .C(_7603_),
    .Y(_7604_)
);

NAND3X1 _17853_ (
    .A(_7336_),
    .B(_7329_),
    .C(_7334_),
    .Y(_7605_)
);

NAND3X1 _17854_ (
    .A(_7224_),
    .B(_7339_),
    .C(_7337_),
    .Y(_7606_)
);

NAND2X1 _17855_ (
    .A(_7605_),
    .B(_7606_),
    .Y(_7607_)
);

OAI21X1 _17856_ (
    .A(_7600_),
    .B(_7601_),
    .C(_7343_),
    .Y(_7608_)
);

NAND3X1 _17857_ (
    .A(_7589_),
    .B(_7596_),
    .C(_7599_),
    .Y(_7609_)
);

NAND3X1 _17858_ (
    .A(_7609_),
    .B(_7607_),
    .C(_7608_),
    .Y(_7610_)
);

NAND3X1 _17859_ (
    .A(_7604_),
    .B(_7610_),
    .C(_7223_),
    .Y(_7611_)
);

NOR3X1 _17860_ (
    .A(_7180_),
    .B(_7181_),
    .C(_7179_),
    .Y(_7612_)
);

AOI21X1 _17861_ (
    .A(_6919_),
    .B(_7182_),
    .C(_7612_),
    .Y(_7613_)
);

AOI21X1 _17862_ (
    .A(_7609_),
    .B(_7608_),
    .C(_7607_),
    .Y(_7614_)
);

AOI21X1 _17863_ (
    .A(_7597_),
    .B(_7603_),
    .C(_7341_),
    .Y(_7615_)
);

OAI21X1 _17864_ (
    .A(_7614_),
    .B(_7615_),
    .C(_7613_),
    .Y(_7616_)
);

NAND3X1 _17865_ (
    .A(_7221_),
    .B(_7611_),
    .C(_7616_),
    .Y(_7617_)
);

INVX2 _17866_ (
    .A(_7221_),
    .Y(_7618_)
);

OAI21X1 _17867_ (
    .A(_7614_),
    .B(_7615_),
    .C(_7223_),
    .Y(_7619_)
);

NAND3X1 _17868_ (
    .A(_7604_),
    .B(_7610_),
    .C(_7613_),
    .Y(_7620_)
);

NAND3X1 _17869_ (
    .A(_7618_),
    .B(_7620_),
    .C(_7619_),
    .Y(_7621_)
);

NAND3X1 _17870_ (
    .A(_7617_),
    .B(_7220_),
    .C(_7621_),
    .Y(_7622_)
);

AOI21X1 _17871_ (
    .A(_6811_),
    .B(_7195_),
    .C(_7199_),
    .Y(_7625_)
);

AOI21X1 _17872_ (
    .A(_7620_),
    .B(_7619_),
    .C(_7618_),
    .Y(_7626_)
);

AOI21X1 _17873_ (
    .A(_7611_),
    .B(_7616_),
    .C(_7221_),
    .Y(_7627_)
);

OAI21X1 _17874_ (
    .A(_7626_),
    .B(_7627_),
    .C(_7625_),
    .Y(_7628_)
);

NAND3X1 _17875_ (
    .A(_7219_),
    .B(_7622_),
    .C(_7628_),
    .Y(_7629_)
);

OAI21X1 _17876_ (
    .A(_7626_),
    .B(_7627_),
    .C(_7220_),
    .Y(_7630_)
);

NAND3X1 _17877_ (
    .A(_7617_),
    .B(_7621_),
    .C(_7625_),
    .Y(_7631_)
);

NAND3X1 _17878_ (
    .A(_6843_),
    .B(_7631_),
    .C(_7630_),
    .Y(_7632_)
);

NAND3X1 _17879_ (
    .A(_7218_),
    .B(_7629_),
    .C(_7632_),
    .Y(_7633_)
);

NAND3X1 _17880_ (
    .A(_6843_),
    .B(_7622_),
    .C(_7628_),
    .Y(_7634_)
);

NAND3X1 _17881_ (
    .A(_7219_),
    .B(_7631_),
    .C(_7630_),
    .Y(_7636_)
);

NAND3X1 _17882_ (
    .A(_7202_),
    .B(_7634_),
    .C(_7636_),
    .Y(_7637_)
);

NAND2X1 _17883_ (
    .A(_7633_),
    .B(_7637_),
    .Y(_7638_)
);

XNOR2X1 _17884_ (
    .A(_7215_),
    .B(_7638_),
    .Y(_0_[31])
);

OAI21X1 _17885_ (
    .A(_5660_),
    .B(_6033_),
    .C(_6029_),
    .Y(_7639_)
);

AOI21X1 _17886_ (
    .A(_6039_),
    .B(_5300_),
    .C(_7639_),
    .Y(_7640_)
);

AOI21X1 _17887_ (
    .A(_7634_),
    .B(_7636_),
    .C(_7202_),
    .Y(_7641_)
);

AOI21X1 _17888_ (
    .A(_7629_),
    .B(_7632_),
    .C(_7218_),
    .Y(_7642_)
);

NOR2X1 _17889_ (
    .A(_7641_),
    .B(_7642_),
    .Y(_7643_)
);

NAND3X1 _17890_ (
    .A(_7213_),
    .B(_6805_),
    .C(_7643_),
    .Y(_7644_)
);

NOR2X1 _17891_ (
    .A(_7214_),
    .B(_7638_),
    .Y(_7646_)
);

OAI21X1 _17892_ (
    .A(_7642_),
    .B(_7209_),
    .C(_7633_),
    .Y(_7647_)
);

AOI21X1 _17893_ (
    .A(_6804_),
    .B(_7646_),
    .C(_7647_),
    .Y(_7648_)
);

OAI21X1 _17894_ (
    .A(_7640_),
    .B(_7644_),
    .C(_7648_),
    .Y(_7649_)
);

NOR2X1 _17895_ (
    .A(_6040_),
    .B(_7644_),
    .Y(_7650_)
);

AOI21X1 _17896_ (
    .A(_7650_),
    .B(_4648_),
    .C(_7649_),
    .Y(_7651_)
);

INVX2 _17897_ (
    .A(_7651_),
    .Y(_7652_)
);

AOI21X1 _17898_ (
    .A(_7617_),
    .B(_7621_),
    .C(_7220_),
    .Y(_7653_)
);

OAI21X1 _17899_ (
    .A(_7653_),
    .B(_6843_),
    .C(_7622_),
    .Y(_7654_)
);

OAI21X1 _17900_ (
    .A(_7259_),
    .B(_7227_),
    .C(_7268_),
    .Y(_7655_)
);

INVX2 _17901_ (
    .A(_7655_),
    .Y(_7657_)
);

AOI21X1 _17902_ (
    .A(_7604_),
    .B(_7610_),
    .C(_7223_),
    .Y(_7658_)
);

OAI21X1 _17903_ (
    .A(_7658_),
    .B(_7618_),
    .C(_7611_),
    .Y(_7659_)
);

NAND2X1 _17904_ (
    .A(_7329_),
    .B(_7605_),
    .Y(_7660_)
);

INVX2 _17905_ (
    .A(_7660_),
    .Y(_7661_)
);

AOI21X1 _17906_ (
    .A(_7589_),
    .B(_7596_),
    .C(_7343_),
    .Y(_7662_)
);

OAI21X1 _17907_ (
    .A(_7607_),
    .B(_7662_),
    .C(_7597_),
    .Y(_7663_)
);

NAND2X1 _17908_ (
    .A(_7314_),
    .B(_7321_),
    .Y(_7664_)
);

NOR2X1 _17909_ (
    .A(_2661_),
    .B(_7225__bF$buf3),
    .Y(_7665_)
);

INVX1 _17910_ (
    .A(_7665_),
    .Y(_7666_)
);

OAI21X1 _17911_ (
    .A(_7247_),
    .B(_7233_),
    .C(_7257_),
    .Y(_7668_)
);

NOR2X1 _17912_ (
    .A(_2519__bF$buf1),
    .B(_6815__bF$buf2),
    .Y(_7669_)
);

INVX2 _17913_ (
    .A(_7669_),
    .Y(_7670_)
);

OAI21X1 _17914_ (
    .A(_7245_),
    .B(_7235_),
    .C(_7240_),
    .Y(_7671_)
);

NAND2X1 _17915_ (
    .A(areg_3_bF$buf1),
    .B(breg_29_bF$buf1),
    .Y(_7672_)
);

INVX2 _17916_ (
    .A(_7672_),
    .Y(_7673_)
);

AND2X2 _17917_ (
    .A(areg_4_bF$buf0),
    .B(breg_28_bF$buf5),
    .Y(_7674_)
);

AND2X2 _17918_ (
    .A(areg_5_bF$buf4),
    .B(breg_27_bF$buf0),
    .Y(_7675_)
);

NAND2X1 _17919_ (
    .A(_7674_),
    .B(_7675_),
    .Y(_7676_)
);

OAI21X1 _17920_ (
    .A(_2825__bF$buf0),
    .B(_5668__bF$buf0),
    .C(_7243_),
    .Y(_7677_)
);

NAND3X1 _17921_ (
    .A(_7673_),
    .B(_7677_),
    .C(_7676_),
    .Y(_7679_)
);

NAND2X1 _17922_ (
    .A(areg_5_bF$buf3),
    .B(breg_27_bF$buf5),
    .Y(_7680_)
);

NOR2X1 _17923_ (
    .A(_7243_),
    .B(_7680_),
    .Y(_7681_)
);

NOR2X1 _17924_ (
    .A(_7674_),
    .B(_7675_),
    .Y(_7682_)
);

OAI21X1 _17925_ (
    .A(_7682_),
    .B(_7681_),
    .C(_7672_),
    .Y(_7683_)
);

AOI21X1 _17926_ (
    .A(_7679_),
    .B(_7683_),
    .C(_7671_),
    .Y(_7684_)
);

AOI21X1 _17927_ (
    .A(_7236_),
    .B(_7241_),
    .C(_7244_),
    .Y(_7685_)
);

OAI21X1 _17928_ (
    .A(_2562__bF$buf1),
    .B(_6050__bF$buf0),
    .C(_7675_),
    .Y(_7686_)
);

OAI21X1 _17929_ (
    .A(_2825__bF$buf4),
    .B(_5668__bF$buf5),
    .C(_7674_),
    .Y(_7687_)
);

AOI21X1 _17930_ (
    .A(_7686_),
    .B(_7687_),
    .C(_7672_),
    .Y(_7688_)
);

AOI21X1 _17931_ (
    .A(_7677_),
    .B(_7676_),
    .C(_7673_),
    .Y(_7690_)
);

NOR3X1 _17932_ (
    .A(_7690_),
    .B(_7685_),
    .C(_7688_),
    .Y(_7691_)
);

OAI21X1 _17933_ (
    .A(_7691_),
    .B(_7684_),
    .C(_7670_),
    .Y(_7692_)
);

OAI21X1 _17934_ (
    .A(_7688_),
    .B(_7690_),
    .C(_7685_),
    .Y(_7693_)
);

NAND3X1 _17935_ (
    .A(_7679_),
    .B(_7671_),
    .C(_7683_),
    .Y(_7694_)
);

NAND3X1 _17936_ (
    .A(_7669_),
    .B(_7693_),
    .C(_7694_),
    .Y(_7695_)
);

AOI21X1 _17937_ (
    .A(_7695_),
    .B(_7692_),
    .C(_7668_),
    .Y(_7696_)
);

AOI21X1 _17938_ (
    .A(_7232_),
    .B(_7256_),
    .C(_7254_),
    .Y(_7697_)
);

AOI21X1 _17939_ (
    .A(_7693_),
    .B(_7694_),
    .C(_7669_),
    .Y(_7698_)
);

NOR3X1 _17940_ (
    .A(_7684_),
    .B(_7670_),
    .C(_7691_),
    .Y(_7699_)
);

NOR3X1 _17941_ (
    .A(_7697_),
    .B(_7698_),
    .C(_7699_),
    .Y(_7701_)
);

OAI21X1 _17942_ (
    .A(_7701_),
    .B(_7696_),
    .C(_7666_),
    .Y(_7702_)
);

OAI21X1 _17943_ (
    .A(_7699_),
    .B(_7698_),
    .C(_7697_),
    .Y(_7703_)
);

NAND3X1 _17944_ (
    .A(_7668_),
    .B(_7695_),
    .C(_7692_),
    .Y(_7704_)
);

NAND3X1 _17945_ (
    .A(_7665_),
    .B(_7704_),
    .C(_7703_),
    .Y(_7705_)
);

AND2X2 _17946_ (
    .A(_7702_),
    .B(_7705_),
    .Y(_7706_)
);

AOI21X1 _17947_ (
    .A(_7295_),
    .B(_7299_),
    .C(_7301_),
    .Y(_7707_)
);

OAI21X1 _17948_ (
    .A(_7707_),
    .B(_7310_),
    .C(_7302_),
    .Y(_7708_)
);

NAND2X1 _17949_ (
    .A(_7288_),
    .B(_7295_),
    .Y(_7709_)
);

OAI21X1 _17950_ (
    .A(_7276_),
    .B(_7277_),
    .C(_7284_),
    .Y(_7710_)
);

NAND2X1 _17951_ (
    .A(areg_6_bF$buf0),
    .B(breg_26_bF$buf3),
    .Y(_7712_)
);

NAND2X1 _17952_ (
    .A(areg_8_bF$buf1),
    .B(breg_24_bF$buf0),
    .Y(_7713_)
);

NOR2X1 _17953_ (
    .A(_7278_),
    .B(_7713_),
    .Y(_7714_)
);

AND2X2 _17954_ (
    .A(_7278_),
    .B(_7713_),
    .Y(_7715_)
);

OAI21X1 _17955_ (
    .A(_7715_),
    .B(_7714_),
    .C(_7712_),
    .Y(_7716_)
);

INVX1 _17956_ (
    .A(_7712_),
    .Y(_7717_)
);

OR2X2 _17957_ (
    .A(_7278_),
    .B(_7713_),
    .Y(_7718_)
);

OAI21X1 _17958_ (
    .A(_5190__bF$buf0),
    .B(_5315__bF$buf1),
    .C(_7278_),
    .Y(_7719_)
);

NAND3X1 _17959_ (
    .A(_7717_),
    .B(_7719_),
    .C(_7718_),
    .Y(_7720_)
);

NAND2X1 _17960_ (
    .A(areg_10_bF$buf0),
    .B(breg_22_bF$buf4),
    .Y(_7721_)
);

OAI22X1 _17961_ (
    .A(_6927_),
    .B(_7721_),
    .C(_7373_),
    .D(_7348_),
    .Y(_7723_)
);

NAND3X1 _17962_ (
    .A(_7716_),
    .B(_7720_),
    .C(_7723_),
    .Y(_7724_)
);

AOI21X1 _17963_ (
    .A(_7719_),
    .B(_7718_),
    .C(_7717_),
    .Y(_7725_)
);

NOR3X1 _17964_ (
    .A(_7712_),
    .B(_7714_),
    .C(_7715_),
    .Y(_7726_)
);

OAI21X1 _17965_ (
    .A(_7711__bF$buf1),
    .B(_3781__bF$buf3),
    .C(_7286_),
    .Y(_7727_)
);

AOI21X1 _17966_ (
    .A(_7345_),
    .B(_7727_),
    .C(_7347_),
    .Y(_7728_)
);

OAI21X1 _17967_ (
    .A(_7726_),
    .B(_7725_),
    .C(_7728_),
    .Y(_7729_)
);

NAND3X1 _17968_ (
    .A(_7710_),
    .B(_7729_),
    .C(_7724_),
    .Y(_7730_)
);

INVX1 _17969_ (
    .A(_7710_),
    .Y(_7731_)
);

NAND3X1 _17970_ (
    .A(_7728_),
    .B(_7716_),
    .C(_7720_),
    .Y(_7732_)
);

OAI21X1 _17971_ (
    .A(_7726_),
    .B(_7725_),
    .C(_7723_),
    .Y(_7734_)
);

NAND3X1 _17972_ (
    .A(_7731_),
    .B(_7732_),
    .C(_7734_),
    .Y(_7735_)
);

AOI21X1 _17973_ (
    .A(_7368_),
    .B(_7369_),
    .C(_7352_),
    .Y(_7736_)
);

OAI21X1 _17974_ (
    .A(_7351_),
    .B(_7736_),
    .C(_7375_),
    .Y(_7737_)
);

NAND3X1 _17975_ (
    .A(_7730_),
    .B(_7735_),
    .C(_7737_),
    .Y(_7738_)
);

AOI21X1 _17976_ (
    .A(_7732_),
    .B(_7734_),
    .C(_7731_),
    .Y(_7739_)
);

AOI21X1 _17977_ (
    .A(_7729_),
    .B(_7724_),
    .C(_7710_),
    .Y(_7740_)
);

NOR3X1 _17978_ (
    .A(_7367_),
    .B(_7365_),
    .C(_7361_),
    .Y(_7741_)
);

AOI21X1 _17979_ (
    .A(_7376_),
    .B(_7374_),
    .C(_7741_),
    .Y(_7742_)
);

OAI21X1 _17980_ (
    .A(_7740_),
    .B(_7739_),
    .C(_7742_),
    .Y(_7743_)
);

NAND3X1 _17981_ (
    .A(_7709_),
    .B(_7743_),
    .C(_7738_),
    .Y(_7745_)
);

INVX2 _17982_ (
    .A(_7709_),
    .Y(_7746_)
);

NOR3X1 _17983_ (
    .A(_7740_),
    .B(_7739_),
    .C(_7742_),
    .Y(_7747_)
);

AOI21X1 _17984_ (
    .A(_7730_),
    .B(_7735_),
    .C(_7737_),
    .Y(_7748_)
);

OAI21X1 _17985_ (
    .A(_7747_),
    .B(_7748_),
    .C(_7746_),
    .Y(_7749_)
);

NAND3X1 _17986_ (
    .A(_7708_),
    .B(_7745_),
    .C(_7749_),
    .Y(_7750_)
);

NAND2X1 _17987_ (
    .A(_7295_),
    .B(_7299_),
    .Y(_7751_)
);

NOR2X1 _17988_ (
    .A(_7307_),
    .B(_7751_),
    .Y(_7752_)
);

AOI21X1 _17989_ (
    .A(_7274_),
    .B(_7308_),
    .C(_7752_),
    .Y(_7753_)
);

NAND3X1 _17990_ (
    .A(_7730_),
    .B(_7735_),
    .C(_7742_),
    .Y(_7754_)
);

OAI21X1 _17991_ (
    .A(_7740_),
    .B(_7739_),
    .C(_7737_),
    .Y(_7756_)
);

AOI21X1 _17992_ (
    .A(_7756_),
    .B(_7754_),
    .C(_7746_),
    .Y(_7757_)
);

AOI21X1 _17993_ (
    .A(_7743_),
    .B(_7738_),
    .C(_7709_),
    .Y(_7758_)
);

OAI21X1 _17994_ (
    .A(_7757_),
    .B(_7758_),
    .C(_7753_),
    .Y(_7759_)
);

NAND3X1 _17995_ (
    .A(_7759_),
    .B(_7750_),
    .C(_7706_),
    .Y(_7760_)
);

NAND2X1 _17996_ (
    .A(_7705_),
    .B(_7702_),
    .Y(_7761_)
);

OAI21X1 _17997_ (
    .A(_7757_),
    .B(_7758_),
    .C(_7708_),
    .Y(_7762_)
);

NAND3X1 _17998_ (
    .A(_7745_),
    .B(_7749_),
    .C(_7753_),
    .Y(_7763_)
);

NAND3X1 _17999_ (
    .A(_7761_),
    .B(_7762_),
    .C(_7763_),
    .Y(_7764_)
);

AOI21X1 _18000_ (
    .A(_7414_),
    .B(_7419_),
    .C(_7421_),
    .Y(_7765_)
);

OAI21X1 _18001_ (
    .A(_7765_),
    .B(_7344_),
    .C(_7422_),
    .Y(_7767_)
);

NAND3X1 _18002_ (
    .A(_7767_),
    .B(_7760_),
    .C(_7764_),
    .Y(_7768_)
);

AOI21X1 _18003_ (
    .A(_7762_),
    .B(_7763_),
    .C(_7761_),
    .Y(_7769_)
);

AOI21X1 _18004_ (
    .A(_7759_),
    .B(_7750_),
    .C(_7706_),
    .Y(_7770_)
);

NOR3X1 _18005_ (
    .A(_7423_),
    .B(_7424_),
    .C(_7427_),
    .Y(_7771_)
);

AOI21X1 _18006_ (
    .A(_7430_),
    .B(_7428_),
    .C(_7771_),
    .Y(_7772_)
);

OAI21X1 _18007_ (
    .A(_7769_),
    .B(_7770_),
    .C(_7772_),
    .Y(_7773_)
);

NAND3X1 _18008_ (
    .A(_7664_),
    .B(_7768_),
    .C(_7773_),
    .Y(_7774_)
);

AND2X2 _18009_ (
    .A(_7321_),
    .B(_7314_),
    .Y(_7775_)
);

NAND3X1 _18010_ (
    .A(_7760_),
    .B(_7764_),
    .C(_7772_),
    .Y(_7776_)
);

OAI21X1 _18011_ (
    .A(_7769_),
    .B(_7770_),
    .C(_7767_),
    .Y(_7778_)
);

NAND3X1 _18012_ (
    .A(_7776_),
    .B(_7778_),
    .C(_7775_),
    .Y(_7779_)
);

NAND2X1 _18013_ (
    .A(_7774_),
    .B(_7779_),
    .Y(_7780_)
);

AOI21X1 _18014_ (
    .A(_7582_),
    .B(_7573_),
    .C(_7436_),
    .Y(_7781_)
);

OAI21X1 _18015_ (
    .A(_7781_),
    .B(_7593_),
    .C(_7583_),
    .Y(_7782_)
);

NAND2X1 _18016_ (
    .A(_7407_),
    .B(_7414_),
    .Y(_7783_)
);

NOR2X1 _18017_ (
    .A(_6582__bF$buf1),
    .B(_5369_),
    .Y(_7784_)
);

INVX1 _18018_ (
    .A(_7784_),
    .Y(_7785_)
);

NAND2X1 _18019_ (
    .A(areg_11_bF$buf0),
    .B(breg_21_bF$buf4),
    .Y(_7786_)
);

NOR2X1 _18020_ (
    .A(_7721_),
    .B(_7786_),
    .Y(_7787_)
);

AND2X2 _18021_ (
    .A(_7721_),
    .B(_7786_),
    .Y(_7789_)
);

NOR2X1 _18022_ (
    .A(_7787_),
    .B(_7789_),
    .Y(_7790_)
);

XNOR2X1 _18023_ (
    .A(_7790_),
    .B(_7785_),
    .Y(_7791_)
);

AOI21X1 _18024_ (
    .A(_7362_),
    .B(_7364_),
    .C(_7356_),
    .Y(_7792_)
);

INVX2 _18025_ (
    .A(_7792_),
    .Y(_7793_)
);

NAND2X1 _18026_ (
    .A(areg_12_bF$buf0),
    .B(breg_20_bF$buf4),
    .Y(_7794_)
);

INVX2 _18027_ (
    .A(_7794_),
    .Y(_7795_)
);

AND2X2 _18028_ (
    .A(areg_13_bF$buf3),
    .B(breg_19_bF$buf0),
    .Y(_7796_)
);

AND2X2 _18029_ (
    .A(areg_14_bF$buf3),
    .B(breg_18_bF$buf5),
    .Y(_7797_)
);

NAND2X1 _18030_ (
    .A(_7796_),
    .B(_7797_),
    .Y(_7798_)
);

OAI22X1 _18031_ (
    .A(_549__bF$buf3),
    .B(_3253__bF$buf1),
    .C(_2287__bF$buf3),
    .D(_3529__bF$buf1),
    .Y(_7800_)
);

NAND3X1 _18032_ (
    .A(_7795_),
    .B(_7800_),
    .C(_7798_),
    .Y(_7801_)
);

NAND2X1 _18033_ (
    .A(areg_14_bF$buf2),
    .B(breg_19_bF$buf5),
    .Y(_7802_)
);

NOR2X1 _18034_ (
    .A(_7355_),
    .B(_7802_),
    .Y(_7803_)
);

NOR2X1 _18035_ (
    .A(_7796_),
    .B(_7797_),
    .Y(_7804_)
);

OAI21X1 _18036_ (
    .A(_7804_),
    .B(_7803_),
    .C(_7794_),
    .Y(_7805_)
);

NAND3X1 _18037_ (
    .A(_7801_),
    .B(_7805_),
    .C(_7793_),
    .Y(_7806_)
);

NOR3X1 _18038_ (
    .A(_7794_),
    .B(_7803_),
    .C(_7804_),
    .Y(_7807_)
);

AOI21X1 _18039_ (
    .A(_7800_),
    .B(_7798_),
    .C(_7795_),
    .Y(_7808_)
);

OAI21X1 _18040_ (
    .A(_7807_),
    .B(_7808_),
    .C(_7792_),
    .Y(_7809_)
);

NAND3X1 _18041_ (
    .A(_7809_),
    .B(_7806_),
    .C(_7791_),
    .Y(_7811_)
);

XNOR2X1 _18042_ (
    .A(_7790_),
    .B(_7784_),
    .Y(_7812_)
);

NOR3X1 _18043_ (
    .A(_7792_),
    .B(_7808_),
    .C(_7807_),
    .Y(_7813_)
);

AOI21X1 _18044_ (
    .A(_7801_),
    .B(_7805_),
    .C(_7793_),
    .Y(_7814_)
);

OAI21X1 _18045_ (
    .A(_7813_),
    .B(_7814_),
    .C(_7812_),
    .Y(_7815_)
);

NAND2X1 _18046_ (
    .A(_7811_),
    .B(_7815_),
    .Y(_7816_)
);

OAI21X1 _18047_ (
    .A(_7405_),
    .B(_7402_),
    .C(_7395_),
    .Y(_7817_)
);

AND2X2 _18048_ (
    .A(areg_16_bF$buf5),
    .B(breg_16_bF$buf0),
    .Y(_7818_)
);

AOI21X1 _18049_ (
    .A(_6964_),
    .B(_7818_),
    .C(_7396_),
    .Y(_7819_)
);

NAND2X1 _18050_ (
    .A(areg_15_bF$buf2),
    .B(breg_17_bF$buf3),
    .Y(_7820_)
);

INVX1 _18051_ (
    .A(_7820_),
    .Y(_7822_)
);

AND2X2 _18052_ (
    .A(breg_15_bF$buf4),
    .B(areg_17_bF$buf4),
    .Y(_7823_)
);

NAND2X1 _18053_ (
    .A(_7818_),
    .B(_7823_),
    .Y(_7824_)
);

NAND2X1 _18054_ (
    .A(areg_16_bF$buf4),
    .B(breg_16_bF$buf5),
    .Y(_7825_)
);

OAI21X1 _18055_ (
    .A(_2362__bF$buf4),
    .B(_2884__bF$buf1),
    .C(_7825_),
    .Y(_7826_)
);

NAND3X1 _18056_ (
    .A(_7822_),
    .B(_7826_),
    .C(_7824_),
    .Y(_7827_)
);

OAI21X1 _18057_ (
    .A(_2669__bF$buf0),
    .B(_2560__bF$buf0),
    .C(_7823_),
    .Y(_7828_)
);

OAI21X1 _18058_ (
    .A(_2362__bF$buf3),
    .B(_2884__bF$buf0),
    .C(_7818_),
    .Y(_7829_)
);

NAND3X1 _18059_ (
    .A(_7820_),
    .B(_7828_),
    .C(_7829_),
    .Y(_7830_)
);

NOR2X1 _18060_ (
    .A(_7392_),
    .B(_7440_),
    .Y(_7831_)
);

OAI21X1 _18061_ (
    .A(_2586__bF$buf4),
    .B(_3402__bF$buf2),
    .C(_7392_),
    .Y(_7833_)
);

AOI21X1 _18062_ (
    .A(_7465_),
    .B(_7833_),
    .C(_7831_),
    .Y(_7834_)
);

NAND3X1 _18063_ (
    .A(_7834_),
    .B(_7827_),
    .C(_7830_),
    .Y(_7835_)
);

AOI21X1 _18064_ (
    .A(_7828_),
    .B(_7829_),
    .C(_7820_),
    .Y(_7836_)
);

AOI21X1 _18065_ (
    .A(_7826_),
    .B(_7824_),
    .C(_7822_),
    .Y(_7837_)
);

NAND2X1 _18066_ (
    .A(breg_13_bF$buf0),
    .B(areg_19_bF$buf0),
    .Y(_7838_)
);

AND2X2 _18067_ (
    .A(_7392_),
    .B(_7440_),
    .Y(_7839_)
);

OAI22X1 _18068_ (
    .A(_7018_),
    .B(_7838_),
    .C(_7839_),
    .D(_7439_),
    .Y(_7840_)
);

OAI21X1 _18069_ (
    .A(_7836_),
    .B(_7837_),
    .C(_7840_),
    .Y(_7841_)
);

AOI21X1 _18070_ (
    .A(_7835_),
    .B(_7841_),
    .C(_7819_),
    .Y(_7842_)
);

OAI21X1 _18071_ (
    .A(_6970_),
    .B(_7825_),
    .C(_7388_),
    .Y(_7844_)
);

NAND3X1 _18072_ (
    .A(_7827_),
    .B(_7830_),
    .C(_7840_),
    .Y(_7845_)
);

OAI21X1 _18073_ (
    .A(_7836_),
    .B(_7837_),
    .C(_7834_),
    .Y(_7846_)
);

AOI21X1 _18074_ (
    .A(_7845_),
    .B(_7846_),
    .C(_7844_),
    .Y(_7847_)
);

OAI21X1 _18075_ (
    .A(_7842_),
    .B(_7847_),
    .C(_7817_),
    .Y(_7848_)
);

AOI21X1 _18076_ (
    .A(_7380_),
    .B(_7400_),
    .C(_7403_),
    .Y(_7849_)
);

NAND3X1 _18077_ (
    .A(_7844_),
    .B(_7845_),
    .C(_7846_),
    .Y(_7850_)
);

NOR3X1 _18078_ (
    .A(_7837_),
    .B(_7834_),
    .C(_7836_),
    .Y(_7851_)
);

AOI21X1 _18079_ (
    .A(_7827_),
    .B(_7830_),
    .C(_7840_),
    .Y(_7852_)
);

OAI21X1 _18080_ (
    .A(_7851_),
    .B(_7852_),
    .C(_7819_),
    .Y(_7853_)
);

NAND3X1 _18081_ (
    .A(_7849_),
    .B(_7850_),
    .C(_7853_),
    .Y(_7855_)
);

AOI21X1 _18082_ (
    .A(_7848_),
    .B(_7855_),
    .C(_7816_),
    .Y(_7856_)
);

OAI21X1 _18083_ (
    .A(_7807_),
    .B(_7808_),
    .C(_7793_),
    .Y(_7857_)
);

NAND3X1 _18084_ (
    .A(_7792_),
    .B(_7801_),
    .C(_7805_),
    .Y(_7858_)
);

AOI21X1 _18085_ (
    .A(_7857_),
    .B(_7858_),
    .C(_7812_),
    .Y(_7859_)
);

AOI21X1 _18086_ (
    .A(_7809_),
    .B(_7806_),
    .C(_7791_),
    .Y(_7860_)
);

NOR2X1 _18087_ (
    .A(_7859_),
    .B(_7860_),
    .Y(_7861_)
);

NAND3X1 _18088_ (
    .A(_7817_),
    .B(_7850_),
    .C(_7853_),
    .Y(_7862_)
);

OAI21X1 _18089_ (
    .A(_7842_),
    .B(_7847_),
    .C(_7849_),
    .Y(_7863_)
);

AOI21X1 _18090_ (
    .A(_7863_),
    .B(_7862_),
    .C(_7861_),
    .Y(_7864_)
);

AOI21X1 _18091_ (
    .A(_7478_),
    .B(_7476_),
    .C(_7479_),
    .Y(_7866_)
);

OAI21X1 _18092_ (
    .A(_7864_),
    .B(_7856_),
    .C(_7866_),
    .Y(_7867_)
);

NAND3X1 _18093_ (
    .A(_7863_),
    .B(_7862_),
    .C(_7861_),
    .Y(_7868_)
);

NAND3X1 _18094_ (
    .A(_7848_),
    .B(_7816_),
    .C(_7855_),
    .Y(_7869_)
);

OAI21X1 _18095_ (
    .A(_7438_),
    .B(_7480_),
    .C(_7472_),
    .Y(_7870_)
);

NAND3X1 _18096_ (
    .A(_7869_),
    .B(_7868_),
    .C(_7870_),
    .Y(_7871_)
);

NAND3X1 _18097_ (
    .A(_7783_),
    .B(_7867_),
    .C(_7871_),
    .Y(_7872_)
);

AND2X2 _18098_ (
    .A(_7414_),
    .B(_7407_),
    .Y(_7873_)
);

AOI21X1 _18099_ (
    .A(_7869_),
    .B(_7868_),
    .C(_7870_),
    .Y(_7874_)
);

NOR3X1 _18100_ (
    .A(_7856_),
    .B(_7864_),
    .C(_7866_),
    .Y(_7875_)
);

OAI21X1 _18101_ (
    .A(_7875_),
    .B(_7874_),
    .C(_7873_),
    .Y(_7877_)
);

NAND2X1 _18102_ (
    .A(_7872_),
    .B(_7877_),
    .Y(_7878_)
);

AOI21X1 _18103_ (
    .A(_7559_),
    .B(_7565_),
    .C(_7485_),
    .Y(_7879_)
);

OAI21X1 _18104_ (
    .A(_7578_),
    .B(_7879_),
    .C(_7566_),
    .Y(_7880_)
);

NAND2X1 _18105_ (
    .A(_7456_),
    .B(_7464_),
    .Y(_7881_)
);

NAND2X1 _18106_ (
    .A(breg_14_bF$buf3),
    .B(areg_18_bF$buf5),
    .Y(_7882_)
);

INVX2 _18107_ (
    .A(_7882_),
    .Y(_7883_)
);

NAND2X1 _18108_ (
    .A(breg_12_bF$buf3),
    .B(areg_20_bF$buf3),
    .Y(_7884_)
);

XOR2X1 _18109_ (
    .A(_7838_),
    .B(_7884_),
    .Y(_7885_)
);

XNOR2X1 _18110_ (
    .A(_7885_),
    .B(_7883_),
    .Y(_7886_)
);

OAI21X1 _18111_ (
    .A(_7454_),
    .B(_7444_),
    .C(_7449_),
    .Y(_7888_)
);

NAND2X1 _18112_ (
    .A(breg_11_bF$buf0),
    .B(areg_21_bF$buf0),
    .Y(_7889_)
);

AND2X2 _18113_ (
    .A(breg_9_bF$buf3),
    .B(areg_23_bF$buf3),
    .Y(_7890_)
);

OAI21X1 _18114_ (
    .A(_7217__bF$buf3),
    .B(_4551__bF$buf2),
    .C(_7890_),
    .Y(_7891_)
);

AND2X2 _18115_ (
    .A(breg_10_bF$buf5),
    .B(areg_22_bF$buf0),
    .Y(_7892_)
);

OAI21X1 _18116_ (
    .A(_6044__bF$buf0),
    .B(_4541__bF$buf2),
    .C(_7892_),
    .Y(_7893_)
);

AOI21X1 _18117_ (
    .A(_7891_),
    .B(_7893_),
    .C(_7889_),
    .Y(_7894_)
);

INVX2 _18118_ (
    .A(_7889_),
    .Y(_7895_)
);

NAND2X1 _18119_ (
    .A(_7892_),
    .B(_7890_),
    .Y(_7896_)
);

OAI21X1 _18120_ (
    .A(_6044__bF$buf5),
    .B(_4541__bF$buf1),
    .C(_7452_),
    .Y(_7897_)
);

AOI21X1 _18121_ (
    .A(_7897_),
    .B(_7896_),
    .C(_7895_),
    .Y(_7899_)
);

OAI21X1 _18122_ (
    .A(_7894_),
    .B(_7899_),
    .C(_7888_),
    .Y(_7900_)
);

AOI21X1 _18123_ (
    .A(_7445_),
    .B(_7450_),
    .C(_7453_),
    .Y(_7901_)
);

NAND3X1 _18124_ (
    .A(_7895_),
    .B(_7897_),
    .C(_7896_),
    .Y(_7902_)
);

NAND2X1 _18125_ (
    .A(breg_9_bF$buf2),
    .B(areg_23_bF$buf2),
    .Y(_7903_)
);

NOR2X1 _18126_ (
    .A(_7452_),
    .B(_7903_),
    .Y(_7904_)
);

NOR2X1 _18127_ (
    .A(_7892_),
    .B(_7890_),
    .Y(_7905_)
);

OAI21X1 _18128_ (
    .A(_7905_),
    .B(_7904_),
    .C(_7889_),
    .Y(_7906_)
);

NAND3X1 _18129_ (
    .A(_7901_),
    .B(_7902_),
    .C(_7906_),
    .Y(_7907_)
);

AOI21X1 _18130_ (
    .A(_7900_),
    .B(_7907_),
    .C(_7886_),
    .Y(_7908_)
);

XNOR2X1 _18131_ (
    .A(_7885_),
    .B(_7882_),
    .Y(_7910_)
);

NAND3X1 _18132_ (
    .A(_7902_),
    .B(_7888_),
    .C(_7906_),
    .Y(_7911_)
);

OAI21X1 _18133_ (
    .A(_7894_),
    .B(_7899_),
    .C(_7901_),
    .Y(_7912_)
);

AOI21X1 _18134_ (
    .A(_7911_),
    .B(_7912_),
    .C(_7910_),
    .Y(_7913_)
);

AOI21X1 _18135_ (
    .A(_7507_),
    .B(_7505_),
    .C(_7508_),
    .Y(_7914_)
);

OAI21X1 _18136_ (
    .A(_7908_),
    .B(_7913_),
    .C(_7914_),
    .Y(_7915_)
);

NAND3X1 _18137_ (
    .A(_7911_),
    .B(_7912_),
    .C(_7910_),
    .Y(_7916_)
);

NAND3X1 _18138_ (
    .A(_7900_),
    .B(_7907_),
    .C(_7886_),
    .Y(_7917_)
);

OAI21X1 _18139_ (
    .A(_7509_),
    .B(_7487_),
    .C(_7500_),
    .Y(_7918_)
);

NAND3X1 _18140_ (
    .A(_7918_),
    .B(_7916_),
    .C(_7917_),
    .Y(_7919_)
);

NAND3X1 _18141_ (
    .A(_7881_),
    .B(_7919_),
    .C(_7915_),
    .Y(_7921_)
);

AND2X2 _18142_ (
    .A(_7464_),
    .B(_7456_),
    .Y(_7922_)
);

AOI21X1 _18143_ (
    .A(_7916_),
    .B(_7917_),
    .C(_7918_),
    .Y(_7923_)
);

NOR3X1 _18144_ (
    .A(_7913_),
    .B(_7914_),
    .C(_7908_),
    .Y(_7924_)
);

OAI21X1 _18145_ (
    .A(_7924_),
    .B(_7923_),
    .C(_7922_),
    .Y(_7925_)
);

NAND2X1 _18146_ (
    .A(_7921_),
    .B(_7925_),
    .Y(_7926_)
);

AOI21X1 _18147_ (
    .A(_7551_),
    .B(_7546_),
    .C(_7513_),
    .Y(_7927_)
);

OAI21X1 _18148_ (
    .A(_7562_),
    .B(_7927_),
    .C(_7552_),
    .Y(_7928_)
);

INVX1 _18149_ (
    .A(_7490_),
    .Y(_7929_)
);

OAI21X1 _18150_ (
    .A(_7493_),
    .B(_7929_),
    .C(_7495_),
    .Y(_7930_)
);

NAND2X1 _18151_ (
    .A(breg[8]),
    .B(areg_24_bF$buf2),
    .Y(_7932_)
);

INVX1 _18152_ (
    .A(_7932_),
    .Y(_7933_)
);

AND2X2 _18153_ (
    .A(breg_7_bF$buf1),
    .B(areg_25_bF$buf4),
    .Y(_7934_)
);

AND2X2 _18154_ (
    .A(breg_6_bF$buf1),
    .B(areg_26_bF$buf0),
    .Y(_7935_)
);

NAND2X1 _18155_ (
    .A(_7934_),
    .B(_7935_),
    .Y(_7936_)
);

OAI22X1 _18156_ (
    .A(_5453__bF$buf5),
    .B(_6686__bF$buf2),
    .C(_4116__bF$buf2),
    .D(_6300__bF$buf0),
    .Y(_7937_)
);

NAND3X1 _18157_ (
    .A(_7933_),
    .B(_7937_),
    .C(_7936_),
    .Y(_7938_)
);

OAI21X1 _18158_ (
    .A(_4116__bF$buf1),
    .B(_6300__bF$buf3),
    .C(_7935_),
    .Y(_7939_)
);

OAI21X1 _18159_ (
    .A(_5453__bF$buf4),
    .B(_6686__bF$buf1),
    .C(_7934_),
    .Y(_7940_)
);

NAND3X1 _18160_ (
    .A(_7932_),
    .B(_7939_),
    .C(_7940_),
    .Y(_7941_)
);

OAI21X1 _18161_ (
    .A(_7524_),
    .B(_7515_),
    .C(_7519_),
    .Y(_7943_)
);

NAND3X1 _18162_ (
    .A(_7938_),
    .B(_7941_),
    .C(_7943_),
    .Y(_7944_)
);

AOI21X1 _18163_ (
    .A(_7939_),
    .B(_7940_),
    .C(_7932_),
    .Y(_7945_)
);

AOI21X1 _18164_ (
    .A(_7937_),
    .B(_7936_),
    .C(_7933_),
    .Y(_7946_)
);

AOI21X1 _18165_ (
    .A(_7516_),
    .B(_7521_),
    .C(_7523_),
    .Y(_7947_)
);

OAI21X1 _18166_ (
    .A(_7945_),
    .B(_7946_),
    .C(_7947_),
    .Y(_7948_)
);

NAND3X1 _18167_ (
    .A(_7930_),
    .B(_7944_),
    .C(_7948_),
    .Y(_7949_)
);

AOI21X1 _18168_ (
    .A(_7070_),
    .B(_7934_),
    .C(_7501_),
    .Y(_7950_)
);

NAND3X1 _18169_ (
    .A(_7947_),
    .B(_7938_),
    .C(_7941_),
    .Y(_7951_)
);

OAI21X1 _18170_ (
    .A(_7945_),
    .B(_7946_),
    .C(_7943_),
    .Y(_7952_)
);

NAND3X1 _18171_ (
    .A(_7950_),
    .B(_7951_),
    .C(_7952_),
    .Y(_7954_)
);

NAND2X1 _18172_ (
    .A(_7949_),
    .B(_7954_),
    .Y(_7955_)
);

AOI21X1 _18173_ (
    .A(_7540_),
    .B(_7535_),
    .C(_7528_),
    .Y(_7956_)
);

OAI21X1 _18174_ (
    .A(_7956_),
    .B(_7548_),
    .C(_7541_),
    .Y(_7957_)
);

NAND2X1 _18175_ (
    .A(breg_5_bF$buf1),
    .B(areg_27_bF$buf1),
    .Y(_7958_)
);

INVX1 _18176_ (
    .A(_7958_),
    .Y(_7959_)
);

AND2X2 _18177_ (
    .A(breg_3_bF$buf2),
    .B(areg_28_bF$buf2),
    .Y(_7960_)
);

AND2X2 _18178_ (
    .A(breg_4_bF$buf0),
    .B(areg_29_bF$buf3),
    .Y(_7961_)
);

AOI22X1 _18179_ (
    .A(breg_3_bF$buf1),
    .B(areg_29_bF$buf2),
    .C(breg_4_bF$buf5),
    .D(areg_28_bF$buf1),
    .Y(_7962_)
);

AOI21X1 _18180_ (
    .A(_7960_),
    .B(_7961_),
    .C(_7962_),
    .Y(_7963_)
);

XNOR2X1 _18181_ (
    .A(_7963_),
    .B(_7959_),
    .Y(_7965_)
);

OAI21X1 _18182_ (
    .A(_7529_),
    .B(_7533_),
    .C(_7532_),
    .Y(_7966_)
);

NAND2X1 _18183_ (
    .A(breg_2_bF$buf1),
    .B(areg_31_bF$buf0),
    .Y(_7967_)
);

NOR2X1 _18184_ (
    .A(_7116_),
    .B(_7967_),
    .Y(_7968_)
);

AOI22X1 _18185_ (
    .A(breg_1_bF$buf0),
    .B(areg_31_bF$buf4),
    .C(breg_2_bF$buf0),
    .D(areg_30_bF$buf5),
    .Y(_7969_)
);

NOR2X1 _18186_ (
    .A(_7969_),
    .B(_7968_),
    .Y(_7970_)
);

AND2X2 _18187_ (
    .A(_7966_),
    .B(_7970_),
    .Y(_7971_)
);

NOR2X1 _18188_ (
    .A(_7970_),
    .B(_7966_),
    .Y(_7972_)
);

NOR3X1 _18189_ (
    .A(_7965_),
    .B(_7972_),
    .C(_7971_),
    .Y(_7973_)
);

XNOR2X1 _18190_ (
    .A(_7963_),
    .B(_7958_),
    .Y(_7974_)
);

NAND2X1 _18191_ (
    .A(_7970_),
    .B(_7966_),
    .Y(_7976_)
);

OR2X2 _18192_ (
    .A(_7966_),
    .B(_7970_),
    .Y(_7977_)
);

AOI21X1 _18193_ (
    .A(_7976_),
    .B(_7977_),
    .C(_7974_),
    .Y(_7978_)
);

OAI21X1 _18194_ (
    .A(_7973_),
    .B(_7978_),
    .C(_7957_),
    .Y(_7979_)
);

NOR3X1 _18195_ (
    .A(_7543_),
    .B(_7542_),
    .C(_7544_),
    .Y(_7980_)
);

AOI21X1 _18196_ (
    .A(_7527_),
    .B(_7545_),
    .C(_7980_),
    .Y(_7981_)
);

NAND3X1 _18197_ (
    .A(_7974_),
    .B(_7976_),
    .C(_7977_),
    .Y(_7982_)
);

OAI21X1 _18198_ (
    .A(_7971_),
    .B(_7972_),
    .C(_7965_),
    .Y(_7983_)
);

NAND3X1 _18199_ (
    .A(_7982_),
    .B(_7983_),
    .C(_7981_),
    .Y(_7984_)
);

AOI21X1 _18200_ (
    .A(_7979_),
    .B(_7984_),
    .C(_7955_),
    .Y(_7985_)
);

AND2X2 _18201_ (
    .A(_7949_),
    .B(_7954_),
    .Y(_7987_)
);

NAND3X1 _18202_ (
    .A(_7982_),
    .B(_7983_),
    .C(_7957_),
    .Y(_7988_)
);

OAI21X1 _18203_ (
    .A(_7973_),
    .B(_7978_),
    .C(_7981_),
    .Y(_7989_)
);

AOI21X1 _18204_ (
    .A(_7988_),
    .B(_7989_),
    .C(_7987_),
    .Y(_7990_)
);

OAI21X1 _18205_ (
    .A(_7985_),
    .B(_7990_),
    .C(_7928_),
    .Y(_7991_)
);

NOR3X1 _18206_ (
    .A(_7555_),
    .B(_7556_),
    .C(_7554_),
    .Y(_7992_)
);

AOI21X1 _18207_ (
    .A(_7511_),
    .B(_7557_),
    .C(_7992_),
    .Y(_7993_)
);

NAND3X1 _18208_ (
    .A(_7988_),
    .B(_7989_),
    .C(_7987_),
    .Y(_7994_)
);

NAND3X1 _18209_ (
    .A(_7955_),
    .B(_7979_),
    .C(_7984_),
    .Y(_7995_)
);

NAND3X1 _18210_ (
    .A(_7994_),
    .B(_7995_),
    .C(_7993_),
    .Y(_7996_)
);

AOI21X1 _18211_ (
    .A(_7991_),
    .B(_7996_),
    .C(_7926_),
    .Y(_7998_)
);

OAI21X1 _18212_ (
    .A(_7924_),
    .B(_7923_),
    .C(_7881_),
    .Y(_7999_)
);

NAND3X1 _18213_ (
    .A(_7919_),
    .B(_7922_),
    .C(_7915_),
    .Y(_8000_)
);

NAND2X1 _18214_ (
    .A(_8000_),
    .B(_7999_),
    .Y(_8001_)
);

NAND3X1 _18215_ (
    .A(_7994_),
    .B(_7995_),
    .C(_7928_),
    .Y(_8002_)
);

OAI21X1 _18216_ (
    .A(_7985_),
    .B(_7990_),
    .C(_7993_),
    .Y(_8003_)
);

AOI21X1 _18217_ (
    .A(_8002_),
    .B(_8003_),
    .C(_8001_),
    .Y(_8004_)
);

OAI21X1 _18218_ (
    .A(_7998_),
    .B(_8004_),
    .C(_7880_),
    .Y(_8005_)
);

NOR3X1 _18219_ (
    .A(_7570_),
    .B(_7571_),
    .C(_7568_),
    .Y(_8006_)
);

AOI21X1 _18220_ (
    .A(_7483_),
    .B(_7572_),
    .C(_8006_),
    .Y(_8007_)
);

NAND3X1 _18221_ (
    .A(_8002_),
    .B(_8003_),
    .C(_8001_),
    .Y(_8009_)
);

NAND3X1 _18222_ (
    .A(_7991_),
    .B(_7996_),
    .C(_7926_),
    .Y(_8010_)
);

NAND3X1 _18223_ (
    .A(_8009_),
    .B(_8010_),
    .C(_8007_),
    .Y(_8011_)
);

AOI21X1 _18224_ (
    .A(_8005_),
    .B(_8011_),
    .C(_7878_),
    .Y(_8012_)
);

OAI21X1 _18225_ (
    .A(_7875_),
    .B(_7874_),
    .C(_7783_),
    .Y(_8013_)
);

NAND3X1 _18226_ (
    .A(_7873_),
    .B(_7867_),
    .C(_7871_),
    .Y(_8014_)
);

NAND2X1 _18227_ (
    .A(_8014_),
    .B(_8013_),
    .Y(_8015_)
);

NAND3X1 _18228_ (
    .A(_7880_),
    .B(_8009_),
    .C(_8010_),
    .Y(_8016_)
);

OAI21X1 _18229_ (
    .A(_7998_),
    .B(_8004_),
    .C(_8007_),
    .Y(_8017_)
);

AOI21X1 _18230_ (
    .A(_8016_),
    .B(_8017_),
    .C(_8015_),
    .Y(_8018_)
);

OAI21X1 _18231_ (
    .A(_8012_),
    .B(_8018_),
    .C(_7782_),
    .Y(_8019_)
);

NOR3X1 _18232_ (
    .A(_7586_),
    .B(_7587_),
    .C(_7585_),
    .Y(_8020_)
);

AOI21X1 _18233_ (
    .A(_7434_),
    .B(_7588_),
    .C(_8020_),
    .Y(_8021_)
);

NAND3X1 _18234_ (
    .A(_8016_),
    .B(_8017_),
    .C(_8015_),
    .Y(_8022_)
);

NAND3X1 _18235_ (
    .A(_8005_),
    .B(_8011_),
    .C(_7878_),
    .Y(_8023_)
);

NAND3X1 _18236_ (
    .A(_8022_),
    .B(_8023_),
    .C(_8021_),
    .Y(_8024_)
);

AOI21X1 _18237_ (
    .A(_8019_),
    .B(_8024_),
    .C(_7780_),
    .Y(_8025_)
);

NAND3X1 _18238_ (
    .A(_7768_),
    .B(_7773_),
    .C(_7775_),
    .Y(_8026_)
);

NAND3X1 _18239_ (
    .A(_7664_),
    .B(_7776_),
    .C(_7778_),
    .Y(_8027_)
);

NAND2X1 _18240_ (
    .A(_8027_),
    .B(_8026_),
    .Y(_8028_)
);

NAND3X1 _18241_ (
    .A(_8022_),
    .B(_7782_),
    .C(_8023_),
    .Y(_8030_)
);

OAI21X1 _18242_ (
    .A(_8012_),
    .B(_8018_),
    .C(_8021_),
    .Y(_8031_)
);

AOI21X1 _18243_ (
    .A(_8030_),
    .B(_8031_),
    .C(_8028_),
    .Y(_8032_)
);

OAI21X1 _18244_ (
    .A(_8025_),
    .B(_8032_),
    .C(_7663_),
    .Y(_8033_)
);

NOR3X1 _18245_ (
    .A(_7600_),
    .B(_7601_),
    .C(_7599_),
    .Y(_8034_)
);

AOI21X1 _18246_ (
    .A(_7341_),
    .B(_7603_),
    .C(_8034_),
    .Y(_8035_)
);

NAND3X1 _18247_ (
    .A(_8030_),
    .B(_8031_),
    .C(_8028_),
    .Y(_8036_)
);

NAND3X1 _18248_ (
    .A(_8019_),
    .B(_8024_),
    .C(_7780_),
    .Y(_8037_)
);

NAND3X1 _18249_ (
    .A(_8036_),
    .B(_8037_),
    .C(_8035_),
    .Y(_8038_)
);

AOI21X1 _18250_ (
    .A(_8033_),
    .B(_8038_),
    .C(_7661_),
    .Y(_8039_)
);

NAND3X1 _18251_ (
    .A(_8036_),
    .B(_8037_),
    .C(_7663_),
    .Y(_8042_)
);

OAI21X1 _18252_ (
    .A(_8025_),
    .B(_8032_),
    .C(_8035_),
    .Y(_8043_)
);

AOI21X1 _18253_ (
    .A(_8042_),
    .B(_8043_),
    .C(_7660_),
    .Y(_8044_)
);

OAI21X1 _18254_ (
    .A(_8039_),
    .B(_8044_),
    .C(_7659_),
    .Y(_8045_)
);

NOR3X1 _18255_ (
    .A(_7614_),
    .B(_7615_),
    .C(_7613_),
    .Y(_8046_)
);

AOI21X1 _18256_ (
    .A(_7221_),
    .B(_7616_),
    .C(_8046_),
    .Y(_8047_)
);

NAND3X1 _18257_ (
    .A(_7660_),
    .B(_8042_),
    .C(_8043_),
    .Y(_8048_)
);

NOR3X1 _18258_ (
    .A(_8025_),
    .B(_8032_),
    .C(_8035_),
    .Y(_8049_)
);

AOI21X1 _18259_ (
    .A(_8036_),
    .B(_8037_),
    .C(_7663_),
    .Y(_8050_)
);

OAI21X1 _18260_ (
    .A(_8049_),
    .B(_8050_),
    .C(_7661_),
    .Y(_8051_)
);

NAND3X1 _18261_ (
    .A(_8047_),
    .B(_8048_),
    .C(_8051_),
    .Y(_8053_)
);

AOI21X1 _18262_ (
    .A(_8045_),
    .B(_8053_),
    .C(_7657_),
    .Y(_8054_)
);

NAND3X1 _18263_ (
    .A(_7659_),
    .B(_8048_),
    .C(_8051_),
    .Y(_8055_)
);

OAI21X1 _18264_ (
    .A(_8039_),
    .B(_8044_),
    .C(_8047_),
    .Y(_8056_)
);

AOI21X1 _18265_ (
    .A(_8056_),
    .B(_8055_),
    .C(_7655_),
    .Y(_8057_)
);

OAI21X1 _18266_ (
    .A(_8054_),
    .B(_8057_),
    .C(_7654_),
    .Y(_8058_)
);

NOR3X1 _18267_ (
    .A(_7626_),
    .B(_7627_),
    .C(_7625_),
    .Y(_8059_)
);

AOI21X1 _18268_ (
    .A(_7219_),
    .B(_7628_),
    .C(_8059_),
    .Y(_8060_)
);

NAND3X1 _18269_ (
    .A(_7655_),
    .B(_8056_),
    .C(_8055_),
    .Y(_8061_)
);

NOR3X1 _18270_ (
    .A(_8039_),
    .B(_8044_),
    .C(_8047_),
    .Y(_8062_)
);

AOI21X1 _18271_ (
    .A(_8048_),
    .B(_8051_),
    .C(_7659_),
    .Y(_8064_)
);

OAI21X1 _18272_ (
    .A(_8062_),
    .B(_8064_),
    .C(_7657_),
    .Y(_8065_)
);

NAND3X1 _18273_ (
    .A(_8060_),
    .B(_8061_),
    .C(_8065_),
    .Y(_8066_)
);

NAND2X1 _18274_ (
    .A(_8058_),
    .B(_8066_),
    .Y(_8067_)
);

XOR2X1 _18275_ (
    .A(_7652_),
    .B(_8067_),
    .Y(_0_[32])
);

NOR3X1 _18276_ (
    .A(_8054_),
    .B(_8057_),
    .C(_8060_),
    .Y(_8068_)
);

AOI21X1 _18277_ (
    .A(_8067_),
    .B(_7652_),
    .C(_8068_),
    .Y(_8069_)
);

OAI21X1 _18278_ (
    .A(_8064_),
    .B(_7657_),
    .C(_8055_),
    .Y(_8070_)
);

OAI21X1 _18279_ (
    .A(_7696_),
    .B(_7666_),
    .C(_7704_),
    .Y(_8071_)
);

INVX2 _18280_ (
    .A(_8071_),
    .Y(_8072_)
);

OAI21X1 _18281_ (
    .A(_8050_),
    .B(_7661_),
    .C(_8042_),
    .Y(_8074_)
);

NAND2X1 _18282_ (
    .A(_7768_),
    .B(_7774_),
    .Y(_8075_)
);

INVX2 _18283_ (
    .A(_8075_),
    .Y(_8076_)
);

AOI21X1 _18284_ (
    .A(_8022_),
    .B(_8023_),
    .C(_7782_),
    .Y(_8077_)
);

OAI21X1 _18285_ (
    .A(_7780_),
    .B(_8077_),
    .C(_8030_),
    .Y(_8078_)
);

NAND2X1 _18286_ (
    .A(_7750_),
    .B(_7760_),
    .Y(_8079_)
);

NOR2X1 _18287_ (
    .A(_2519__bF$buf0),
    .B(_7225__bF$buf2),
    .Y(_8080_)
);

INVX1 _18288_ (
    .A(_8080_),
    .Y(_8081_)
);

OAI21X1 _18289_ (
    .A(_7684_),
    .B(_7670_),
    .C(_7694_),
    .Y(_8082_)
);

NOR2X1 _18290_ (
    .A(_2792_),
    .B(_6815__bF$buf1),
    .Y(_8083_)
);

INVX2 _18291_ (
    .A(_8083_),
    .Y(_8085_)
);

OAI21X1 _18292_ (
    .A(_7682_),
    .B(_7672_),
    .C(_7676_),
    .Y(_8086_)
);

NAND2X1 _18293_ (
    .A(areg_4_bF$buf4),
    .B(breg_29_bF$buf0),
    .Y(_8087_)
);

INVX2 _18294_ (
    .A(_8087_),
    .Y(_8088_)
);

AND2X2 _18295_ (
    .A(areg_5_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_8089_)
);

AND2X2 _18296_ (
    .A(areg_6_bF$buf4),
    .B(breg_27_bF$buf4),
    .Y(_8090_)
);

NAND2X1 _18297_ (
    .A(_8089_),
    .B(_8090_),
    .Y(_8091_)
);

OAI22X1 _18298_ (
    .A(_2825__bF$buf3),
    .B(_6050__bF$buf3),
    .C(_3646__bF$buf0),
    .D(_5668__bF$buf4),
    .Y(_8092_)
);

NAND3X1 _18299_ (
    .A(_8088_),
    .B(_8092_),
    .C(_8091_),
    .Y(_8093_)
);

NAND2X1 _18300_ (
    .A(areg_6_bF$buf3),
    .B(breg_28_bF$buf3),
    .Y(_8094_)
);

NOR2X1 _18301_ (
    .A(_7680_),
    .B(_8094_),
    .Y(_8096_)
);

NOR2X1 _18302_ (
    .A(_8089_),
    .B(_8090_),
    .Y(_8097_)
);

OAI21X1 _18303_ (
    .A(_8097_),
    .B(_8096_),
    .C(_8087_),
    .Y(_8098_)
);

AOI21X1 _18304_ (
    .A(_8093_),
    .B(_8098_),
    .C(_8086_),
    .Y(_8099_)
);

AOI21X1 _18305_ (
    .A(_7673_),
    .B(_7677_),
    .C(_7681_),
    .Y(_8100_)
);

OAI21X1 _18306_ (
    .A(_2825__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_8090_),
    .Y(_8101_)
);

OAI21X1 _18307_ (
    .A(_3646__bF$buf3),
    .B(_5668__bF$buf3),
    .C(_8089_),
    .Y(_8102_)
);

AOI21X1 _18308_ (
    .A(_8101_),
    .B(_8102_),
    .C(_8087_),
    .Y(_8103_)
);

AOI21X1 _18309_ (
    .A(_8092_),
    .B(_8091_),
    .C(_8088_),
    .Y(_8104_)
);

NOR3X1 _18310_ (
    .A(_8104_),
    .B(_8100_),
    .C(_8103_),
    .Y(_8105_)
);

OAI21X1 _18311_ (
    .A(_8105_),
    .B(_8099_),
    .C(_8085_),
    .Y(_8107_)
);

OAI21X1 _18312_ (
    .A(_8103_),
    .B(_8104_),
    .C(_8100_),
    .Y(_8108_)
);

NAND3X1 _18313_ (
    .A(_8093_),
    .B(_8086_),
    .C(_8098_),
    .Y(_8109_)
);

NAND3X1 _18314_ (
    .A(_8083_),
    .B(_8108_),
    .C(_8109_),
    .Y(_8110_)
);

AOI21X1 _18315_ (
    .A(_8110_),
    .B(_8107_),
    .C(_8082_),
    .Y(_8111_)
);

AOI21X1 _18316_ (
    .A(_7669_),
    .B(_7693_),
    .C(_7691_),
    .Y(_8112_)
);

AOI21X1 _18317_ (
    .A(_8108_),
    .B(_8109_),
    .C(_8083_),
    .Y(_8113_)
);

NOR3X1 _18318_ (
    .A(_8099_),
    .B(_8085_),
    .C(_8105_),
    .Y(_8114_)
);

NOR3X1 _18319_ (
    .A(_8112_),
    .B(_8113_),
    .C(_8114_),
    .Y(_8115_)
);

OAI21X1 _18320_ (
    .A(_8115_),
    .B(_8111_),
    .C(_8081_),
    .Y(_8116_)
);

OAI21X1 _18321_ (
    .A(_8114_),
    .B(_8113_),
    .C(_8112_),
    .Y(_8118_)
);

NAND3X1 _18322_ (
    .A(_8082_),
    .B(_8110_),
    .C(_8107_),
    .Y(_8119_)
);

NAND3X1 _18323_ (
    .A(_8080_),
    .B(_8119_),
    .C(_8118_),
    .Y(_8120_)
);

AND2X2 _18324_ (
    .A(_8116_),
    .B(_8120_),
    .Y(_8121_)
);

OAI21X1 _18325_ (
    .A(_7746_),
    .B(_7748_),
    .C(_7738_),
    .Y(_8122_)
);

NAND2X1 _18326_ (
    .A(_7724_),
    .B(_7730_),
    .Y(_8123_)
);

OAI21X1 _18327_ (
    .A(_7715_),
    .B(_7712_),
    .C(_7718_),
    .Y(_8124_)
);

NAND2X1 _18328_ (
    .A(areg_7_bF$buf0),
    .B(breg_26_bF$buf2),
    .Y(_8125_)
);

NAND2X1 _18329_ (
    .A(areg_8_bF$buf0),
    .B(breg_25_bF$buf4),
    .Y(_8126_)
);

NAND2X1 _18330_ (
    .A(areg_9_bF$buf0),
    .B(breg_24_bF$buf5),
    .Y(_8127_)
);

NOR2X1 _18331_ (
    .A(_8126_),
    .B(_8127_),
    .Y(_8129_)
);

AND2X2 _18332_ (
    .A(_8126_),
    .B(_8127_),
    .Y(_8130_)
);

OAI21X1 _18333_ (
    .A(_8130_),
    .B(_8129_),
    .C(_8125_),
    .Y(_8131_)
);

INVX1 _18334_ (
    .A(_8125_),
    .Y(_8132_)
);

OR2X2 _18335_ (
    .A(_8126_),
    .B(_8127_),
    .Y(_8133_)
);

OAI21X1 _18336_ (
    .A(_6582__bF$buf0),
    .B(_5315__bF$buf0),
    .C(_8126_),
    .Y(_8134_)
);

NAND3X1 _18337_ (
    .A(_8132_),
    .B(_8134_),
    .C(_8133_),
    .Y(_8135_)
);

OAI21X1 _18338_ (
    .A(_9104__bF$buf3),
    .B(_3781__bF$buf2),
    .C(_7721_),
    .Y(_8136_)
);

AOI21X1 _18339_ (
    .A(_7784_),
    .B(_8136_),
    .C(_7787_),
    .Y(_8137_)
);

INVX1 _18340_ (
    .A(_8137_),
    .Y(_8138_)
);

NAND3X1 _18341_ (
    .A(_8131_),
    .B(_8135_),
    .C(_8138_),
    .Y(_8140_)
);

AOI21X1 _18342_ (
    .A(_8134_),
    .B(_8133_),
    .C(_8132_),
    .Y(_8141_)
);

NOR3X1 _18343_ (
    .A(_8125_),
    .B(_8129_),
    .C(_8130_),
    .Y(_8142_)
);

OAI21X1 _18344_ (
    .A(_8142_),
    .B(_8141_),
    .C(_8137_),
    .Y(_8143_)
);

NAND3X1 _18345_ (
    .A(_8124_),
    .B(_8143_),
    .C(_8140_),
    .Y(_8144_)
);

INVX1 _18346_ (
    .A(_8124_),
    .Y(_8145_)
);

NAND3X1 _18347_ (
    .A(_8137_),
    .B(_8131_),
    .C(_8135_),
    .Y(_8146_)
);

OAI21X1 _18348_ (
    .A(_8142_),
    .B(_8141_),
    .C(_8138_),
    .Y(_8147_)
);

NAND3X1 _18349_ (
    .A(_8145_),
    .B(_8146_),
    .C(_8147_),
    .Y(_8148_)
);

OAI21X1 _18350_ (
    .A(_7812_),
    .B(_7814_),
    .C(_7806_),
    .Y(_8149_)
);

NAND3X1 _18351_ (
    .A(_8144_),
    .B(_8148_),
    .C(_8149_),
    .Y(_8151_)
);

AOI21X1 _18352_ (
    .A(_8146_),
    .B(_8147_),
    .C(_8145_),
    .Y(_8152_)
);

AOI21X1 _18353_ (
    .A(_8143_),
    .B(_8140_),
    .C(_8124_),
    .Y(_8153_)
);

AOI21X1 _18354_ (
    .A(_7809_),
    .B(_7791_),
    .C(_7813_),
    .Y(_8154_)
);

OAI21X1 _18355_ (
    .A(_8153_),
    .B(_8152_),
    .C(_8154_),
    .Y(_8155_)
);

NAND3X1 _18356_ (
    .A(_8123_),
    .B(_8151_),
    .C(_8155_),
    .Y(_8156_)
);

AND2X2 _18357_ (
    .A(_7730_),
    .B(_7724_),
    .Y(_8157_)
);

NAND3X1 _18358_ (
    .A(_8144_),
    .B(_8148_),
    .C(_8154_),
    .Y(_8158_)
);

OAI21X1 _18359_ (
    .A(_8153_),
    .B(_8152_),
    .C(_8149_),
    .Y(_8159_)
);

NAND3X1 _18360_ (
    .A(_8157_),
    .B(_8158_),
    .C(_8159_),
    .Y(_8160_)
);

NAND3X1 _18361_ (
    .A(_8156_),
    .B(_8160_),
    .C(_8122_),
    .Y(_8162_)
);

AOI21X1 _18362_ (
    .A(_7709_),
    .B(_7743_),
    .C(_7747_),
    .Y(_8163_)
);

AOI21X1 _18363_ (
    .A(_8158_),
    .B(_8159_),
    .C(_8157_),
    .Y(_8164_)
);

AOI21X1 _18364_ (
    .A(_8151_),
    .B(_8155_),
    .C(_8123_),
    .Y(_8165_)
);

OAI21X1 _18365_ (
    .A(_8164_),
    .B(_8165_),
    .C(_8163_),
    .Y(_8166_)
);

NAND3X1 _18366_ (
    .A(_8162_),
    .B(_8166_),
    .C(_8121_),
    .Y(_8167_)
);

NAND2X1 _18367_ (
    .A(_8120_),
    .B(_8116_),
    .Y(_8168_)
);

OAI21X1 _18368_ (
    .A(_8164_),
    .B(_8165_),
    .C(_8122_),
    .Y(_8169_)
);

NAND3X1 _18369_ (
    .A(_8156_),
    .B(_8160_),
    .C(_8163_),
    .Y(_8170_)
);

NAND3X1 _18370_ (
    .A(_8168_),
    .B(_8170_),
    .C(_8169_),
    .Y(_8171_)
);

OAI21X1 _18371_ (
    .A(_7874_),
    .B(_7873_),
    .C(_7871_),
    .Y(_8173_)
);

NAND3X1 _18372_ (
    .A(_8173_),
    .B(_8171_),
    .C(_8167_),
    .Y(_8174_)
);

AOI21X1 _18373_ (
    .A(_8170_),
    .B(_8169_),
    .C(_8168_),
    .Y(_8175_)
);

AOI21X1 _18374_ (
    .A(_8162_),
    .B(_8166_),
    .C(_8121_),
    .Y(_8176_)
);

AOI21X1 _18375_ (
    .A(_7783_),
    .B(_7867_),
    .C(_7875_),
    .Y(_8177_)
);

OAI21X1 _18376_ (
    .A(_8176_),
    .B(_8175_),
    .C(_8177_),
    .Y(_8178_)
);

NAND3X1 _18377_ (
    .A(_8079_),
    .B(_8174_),
    .C(_8178_),
    .Y(_8179_)
);

AND2X2 _18378_ (
    .A(_7760_),
    .B(_7750_),
    .Y(_8180_)
);

NAND3X1 _18379_ (
    .A(_8177_),
    .B(_8171_),
    .C(_8167_),
    .Y(_8181_)
);

OAI21X1 _18380_ (
    .A(_8176_),
    .B(_8175_),
    .C(_8173_),
    .Y(_8182_)
);

NAND3X1 _18381_ (
    .A(_8181_),
    .B(_8180_),
    .C(_8182_),
    .Y(_8184_)
);

NAND2X1 _18382_ (
    .A(_8179_),
    .B(_8184_),
    .Y(_8185_)
);

AOI21X1 _18383_ (
    .A(_8009_),
    .B(_8010_),
    .C(_7880_),
    .Y(_8186_)
);

OAI21X1 _18384_ (
    .A(_7878_),
    .B(_8186_),
    .C(_8016_),
    .Y(_8187_)
);

NAND2X1 _18385_ (
    .A(_7862_),
    .B(_7868_),
    .Y(_8188_)
);

NAND2X1 _18386_ (
    .A(areg_10_bF$buf4),
    .B(breg_23_bF$buf3),
    .Y(_8189_)
);

INVX2 _18387_ (
    .A(_8189_),
    .Y(_8190_)
);

NAND2X1 _18388_ (
    .A(areg_11_bF$buf4),
    .B(breg_22_bF$buf3),
    .Y(_8191_)
);

NAND2X1 _18389_ (
    .A(areg_12_bF$buf4),
    .B(breg_21_bF$buf3),
    .Y(_8192_)
);

XOR2X1 _18390_ (
    .A(_8191_),
    .B(_8192_),
    .Y(_8193_)
);

XNOR2X1 _18391_ (
    .A(_8193_),
    .B(_8190_),
    .Y(_8195_)
);

OAI21X1 _18392_ (
    .A(_7804_),
    .B(_7794_),
    .C(_7798_),
    .Y(_8196_)
);

NAND2X1 _18393_ (
    .A(areg_13_bF$buf2),
    .B(breg_20_bF$buf3),
    .Y(_8197_)
);

AND2X2 _18394_ (
    .A(areg_15_bF$buf1),
    .B(breg_18_bF$buf4),
    .Y(_8198_)
);

OAI21X1 _18395_ (
    .A(_2287__bF$buf2),
    .B(_3253__bF$buf0),
    .C(_8198_),
    .Y(_8199_)
);

AND2X2 _18396_ (
    .A(areg_14_bF$buf1),
    .B(breg_19_bF$buf4),
    .Y(_8200_)
);

OAI21X1 _18397_ (
    .A(_2465__bF$buf4),
    .B(_3529__bF$buf0),
    .C(_8200_),
    .Y(_8201_)
);

AOI21X1 _18398_ (
    .A(_8199_),
    .B(_8201_),
    .C(_8197_),
    .Y(_8202_)
);

INVX2 _18399_ (
    .A(_8197_),
    .Y(_8203_)
);

NAND2X1 _18400_ (
    .A(_8200_),
    .B(_8198_),
    .Y(_8204_)
);

OAI21X1 _18401_ (
    .A(_2465__bF$buf3),
    .B(_3529__bF$buf4),
    .C(_7802_),
    .Y(_8206_)
);

AOI21X1 _18402_ (
    .A(_8206_),
    .B(_8204_),
    .C(_8203_),
    .Y(_8207_)
);

OAI21X1 _18403_ (
    .A(_8202_),
    .B(_8207_),
    .C(_8196_),
    .Y(_8208_)
);

AOI21X1 _18404_ (
    .A(_7795_),
    .B(_7800_),
    .C(_7803_),
    .Y(_8209_)
);

NAND3X1 _18405_ (
    .A(_8203_),
    .B(_8206_),
    .C(_8204_),
    .Y(_8210_)
);

NAND2X1 _18406_ (
    .A(areg_15_bF$buf0),
    .B(breg_18_bF$buf3),
    .Y(_8211_)
);

NOR2X1 _18407_ (
    .A(_7802_),
    .B(_8211_),
    .Y(_8212_)
);

NOR2X1 _18408_ (
    .A(_8200_),
    .B(_8198_),
    .Y(_8213_)
);

OAI21X1 _18409_ (
    .A(_8213_),
    .B(_8212_),
    .C(_8197_),
    .Y(_8214_)
);

NAND3X1 _18410_ (
    .A(_8209_),
    .B(_8210_),
    .C(_8214_),
    .Y(_8215_)
);

AOI21X1 _18411_ (
    .A(_8208_),
    .B(_8215_),
    .C(_8195_),
    .Y(_8217_)
);

XNOR2X1 _18412_ (
    .A(_8193_),
    .B(_8189_),
    .Y(_8218_)
);

NAND3X1 _18413_ (
    .A(_8210_),
    .B(_8196_),
    .C(_8214_),
    .Y(_8219_)
);

OAI21X1 _18414_ (
    .A(_8202_),
    .B(_8207_),
    .C(_8209_),
    .Y(_8220_)
);

AOI21X1 _18415_ (
    .A(_8219_),
    .B(_8220_),
    .C(_8218_),
    .Y(_8221_)
);

OR2X2 _18416_ (
    .A(_8217_),
    .B(_8221_),
    .Y(_8222_)
);

OAI21X1 _18417_ (
    .A(_7852_),
    .B(_7819_),
    .C(_7845_),
    .Y(_8223_)
);

AND2X2 _18418_ (
    .A(breg_16_bF$buf4),
    .B(areg_17_bF$buf3),
    .Y(_8224_)
);

AOI21X1 _18419_ (
    .A(_7385_),
    .B(_8224_),
    .C(_7836_),
    .Y(_8225_)
);

NAND2X1 _18420_ (
    .A(areg_16_bF$buf3),
    .B(breg_17_bF$buf2),
    .Y(_8226_)
);

INVX1 _18421_ (
    .A(_8226_),
    .Y(_8228_)
);

AND2X2 _18422_ (
    .A(breg_15_bF$buf3),
    .B(areg_18_bF$buf4),
    .Y(_8229_)
);

NAND2X1 _18423_ (
    .A(_8224_),
    .B(_8229_),
    .Y(_8230_)
);

OAI22X1 _18424_ (
    .A(_2362__bF$buf2),
    .B(_3146__bF$buf0),
    .C(_2560__bF$buf4),
    .D(_2884__bF$buf3),
    .Y(_8231_)
);

NAND3X1 _18425_ (
    .A(_8228_),
    .B(_8231_),
    .C(_8230_),
    .Y(_8232_)
);

OAI21X1 _18426_ (
    .A(_2560__bF$buf3),
    .B(_2884__bF$buf2),
    .C(_8229_),
    .Y(_8233_)
);

OAI21X1 _18427_ (
    .A(_2362__bF$buf1),
    .B(_3146__bF$buf3),
    .C(_8224_),
    .Y(_8234_)
);

NAND3X1 _18428_ (
    .A(_8226_),
    .B(_8233_),
    .C(_8234_),
    .Y(_8235_)
);

NOR2X1 _18429_ (
    .A(_7838_),
    .B(_7884_),
    .Y(_8236_)
);

OAI21X1 _18430_ (
    .A(_2586__bF$buf3),
    .B(_3958__bF$buf3),
    .C(_7838_),
    .Y(_8237_)
);

AOI21X1 _18431_ (
    .A(_7883_),
    .B(_8237_),
    .C(_8236_),
    .Y(_8239_)
);

NAND3X1 _18432_ (
    .A(_8239_),
    .B(_8232_),
    .C(_8235_),
    .Y(_8240_)
);

AOI21X1 _18433_ (
    .A(_8233_),
    .B(_8234_),
    .C(_8226_),
    .Y(_8241_)
);

AOI21X1 _18434_ (
    .A(_8231_),
    .B(_8230_),
    .C(_8228_),
    .Y(_8242_)
);

NAND2X1 _18435_ (
    .A(breg_13_bF$buf4),
    .B(areg_20_bF$buf2),
    .Y(_8243_)
);

AND2X2 _18436_ (
    .A(_7838_),
    .B(_7884_),
    .Y(_8244_)
);

OAI22X1 _18437_ (
    .A(_7440_),
    .B(_8243_),
    .C(_8244_),
    .D(_7882_),
    .Y(_8245_)
);

OAI21X1 _18438_ (
    .A(_8241_),
    .B(_8242_),
    .C(_8245_),
    .Y(_8246_)
);

AOI21X1 _18439_ (
    .A(_8240_),
    .B(_8246_),
    .C(_8225_),
    .Y(_8247_)
);

INVX1 _18440_ (
    .A(_7823_),
    .Y(_8248_)
);

OAI21X1 _18441_ (
    .A(_7825_),
    .B(_8248_),
    .C(_7827_),
    .Y(_8250_)
);

NAND3X1 _18442_ (
    .A(_8232_),
    .B(_8235_),
    .C(_8245_),
    .Y(_8251_)
);

OAI21X1 _18443_ (
    .A(_8241_),
    .B(_8242_),
    .C(_8239_),
    .Y(_8252_)
);

AOI21X1 _18444_ (
    .A(_8251_),
    .B(_8252_),
    .C(_8250_),
    .Y(_8253_)
);

OAI21X1 _18445_ (
    .A(_8247_),
    .B(_8253_),
    .C(_8223_),
    .Y(_8254_)
);

AOI21X1 _18446_ (
    .A(_7844_),
    .B(_7846_),
    .C(_7851_),
    .Y(_8255_)
);

NAND3X1 _18447_ (
    .A(_8250_),
    .B(_8251_),
    .C(_8252_),
    .Y(_8256_)
);

NOR3X1 _18448_ (
    .A(_8242_),
    .B(_8239_),
    .C(_8241_),
    .Y(_8257_)
);

AOI21X1 _18449_ (
    .A(_8232_),
    .B(_8235_),
    .C(_8245_),
    .Y(_8258_)
);

OAI21X1 _18450_ (
    .A(_8257_),
    .B(_8258_),
    .C(_8225_),
    .Y(_8259_)
);

NAND3X1 _18451_ (
    .A(_8255_),
    .B(_8256_),
    .C(_8259_),
    .Y(_8261_)
);

AOI21X1 _18452_ (
    .A(_8254_),
    .B(_8261_),
    .C(_8222_),
    .Y(_8262_)
);

NOR2X1 _18453_ (
    .A(_8221_),
    .B(_8217_),
    .Y(_8263_)
);

NAND3X1 _18454_ (
    .A(_8223_),
    .B(_8256_),
    .C(_8259_),
    .Y(_8264_)
);

OAI21X1 _18455_ (
    .A(_8247_),
    .B(_8253_),
    .C(_8255_),
    .Y(_8265_)
);

AOI21X1 _18456_ (
    .A(_8265_),
    .B(_8264_),
    .C(_8263_),
    .Y(_8266_)
);

AOI21X1 _18457_ (
    .A(_7881_),
    .B(_7915_),
    .C(_7924_),
    .Y(_8267_)
);

OAI21X1 _18458_ (
    .A(_8262_),
    .B(_8266_),
    .C(_8267_),
    .Y(_8268_)
);

NAND3X1 _18459_ (
    .A(_8263_),
    .B(_8265_),
    .C(_8264_),
    .Y(_8269_)
);

NAND3X1 _18460_ (
    .A(_8254_),
    .B(_8261_),
    .C(_8222_),
    .Y(_8270_)
);

OAI21X1 _18461_ (
    .A(_7923_),
    .B(_7922_),
    .C(_7919_),
    .Y(_8272_)
);

NAND3X1 _18462_ (
    .A(_8269_),
    .B(_8270_),
    .C(_8272_),
    .Y(_8273_)
);

NAND3X1 _18463_ (
    .A(_8188_),
    .B(_8273_),
    .C(_8268_),
    .Y(_8274_)
);

AND2X2 _18464_ (
    .A(_7868_),
    .B(_7862_),
    .Y(_8275_)
);

AOI21X1 _18465_ (
    .A(_8269_),
    .B(_8270_),
    .C(_8272_),
    .Y(_8276_)
);

NOR3X1 _18466_ (
    .A(_8262_),
    .B(_8266_),
    .C(_8267_),
    .Y(_8277_)
);

OAI21X1 _18467_ (
    .A(_8277_),
    .B(_8276_),
    .C(_8275_),
    .Y(_8278_)
);

NAND2X1 _18468_ (
    .A(_8274_),
    .B(_8278_),
    .Y(_8279_)
);

AOI21X1 _18469_ (
    .A(_7994_),
    .B(_7995_),
    .C(_7928_),
    .Y(_8280_)
);

OAI21X1 _18470_ (
    .A(_7926_),
    .B(_8280_),
    .C(_8002_),
    .Y(_8281_)
);

NAND2X1 _18471_ (
    .A(_7911_),
    .B(_7916_),
    .Y(_8283_)
);

NAND2X1 _18472_ (
    .A(breg_14_bF$buf2),
    .B(areg_19_bF$buf5),
    .Y(_8284_)
);

INVX2 _18473_ (
    .A(_8284_),
    .Y(_8285_)
);

NAND2X1 _18474_ (
    .A(breg_12_bF$buf2),
    .B(areg_21_bF$buf4),
    .Y(_8286_)
);

XOR2X1 _18475_ (
    .A(_8243_),
    .B(_8286_),
    .Y(_8287_)
);

XNOR2X1 _18476_ (
    .A(_8287_),
    .B(_8285_),
    .Y(_8288_)
);

OAI21X1 _18477_ (
    .A(_7905_),
    .B(_7889_),
    .C(_7896_),
    .Y(_8289_)
);

NAND2X1 _18478_ (
    .A(breg_11_bF$buf4),
    .B(areg_22_bF$buf4),
    .Y(_8290_)
);

AND2X2 _18479_ (
    .A(breg_9_bF$buf1),
    .B(areg_24_bF$buf1),
    .Y(_8291_)
);

OAI21X1 _18480_ (
    .A(_7217__bF$buf2),
    .B(_4541__bF$buf0),
    .C(_8291_),
    .Y(_8292_)
);

AND2X2 _18481_ (
    .A(breg_10_bF$buf4),
    .B(areg_23_bF$buf1),
    .Y(_8294_)
);

OAI21X1 _18482_ (
    .A(_6044__bF$buf4),
    .B(_5921__bF$buf3),
    .C(_8294_),
    .Y(_8295_)
);

AOI21X1 _18483_ (
    .A(_8292_),
    .B(_8295_),
    .C(_8290_),
    .Y(_8296_)
);

INVX2 _18484_ (
    .A(_8290_),
    .Y(_8297_)
);

NAND2X1 _18485_ (
    .A(_8294_),
    .B(_8291_),
    .Y(_8298_)
);

OAI22X1 _18486_ (
    .A(_6044__bF$buf3),
    .B(_5921__bF$buf2),
    .C(_7217__bF$buf1),
    .D(_4541__bF$buf4),
    .Y(_8299_)
);

AOI21X1 _18487_ (
    .A(_8299_),
    .B(_8298_),
    .C(_8297_),
    .Y(_8300_)
);

OAI21X1 _18488_ (
    .A(_8296_),
    .B(_8300_),
    .C(_8289_),
    .Y(_8301_)
);

AOI21X1 _18489_ (
    .A(_7895_),
    .B(_7897_),
    .C(_7904_),
    .Y(_8302_)
);

NAND3X1 _18490_ (
    .A(_8297_),
    .B(_8299_),
    .C(_8298_),
    .Y(_8303_)
);

NAND2X1 _18491_ (
    .A(breg_10_bF$buf3),
    .B(areg_24_bF$buf0),
    .Y(_8305_)
);

NOR2X1 _18492_ (
    .A(_7903_),
    .B(_8305_),
    .Y(_8306_)
);

NOR2X1 _18493_ (
    .A(_8294_),
    .B(_8291_),
    .Y(_8307_)
);

OAI21X1 _18494_ (
    .A(_8307_),
    .B(_8306_),
    .C(_8290_),
    .Y(_8308_)
);

NAND3X1 _18495_ (
    .A(_8302_),
    .B(_8303_),
    .C(_8308_),
    .Y(_8309_)
);

AOI21X1 _18496_ (
    .A(_8301_),
    .B(_8309_),
    .C(_8288_),
    .Y(_8310_)
);

XNOR2X1 _18497_ (
    .A(_8287_),
    .B(_8284_),
    .Y(_8311_)
);

NAND3X1 _18498_ (
    .A(_8303_),
    .B(_8289_),
    .C(_8308_),
    .Y(_8312_)
);

OAI21X1 _18499_ (
    .A(_8296_),
    .B(_8300_),
    .C(_8302_),
    .Y(_8313_)
);

AOI21X1 _18500_ (
    .A(_8312_),
    .B(_8313_),
    .C(_8311_),
    .Y(_8314_)
);

NOR3X1 _18501_ (
    .A(_7946_),
    .B(_7947_),
    .C(_7945_),
    .Y(_8316_)
);

AOI21X1 _18502_ (
    .A(_7930_),
    .B(_7948_),
    .C(_8316_),
    .Y(_8317_)
);

OAI21X1 _18503_ (
    .A(_8310_),
    .B(_8314_),
    .C(_8317_),
    .Y(_8318_)
);

NAND3X1 _18504_ (
    .A(_8312_),
    .B(_8313_),
    .C(_8311_),
    .Y(_8319_)
);

NAND3X1 _18505_ (
    .A(_8301_),
    .B(_8309_),
    .C(_8288_),
    .Y(_8320_)
);

AOI21X1 _18506_ (
    .A(_7938_),
    .B(_7941_),
    .C(_7943_),
    .Y(_8321_)
);

OAI21X1 _18507_ (
    .A(_8321_),
    .B(_7950_),
    .C(_7944_),
    .Y(_8322_)
);

NAND3X1 _18508_ (
    .A(_8322_),
    .B(_8319_),
    .C(_8320_),
    .Y(_8323_)
);

NAND3X1 _18509_ (
    .A(_8283_),
    .B(_8323_),
    .C(_8318_),
    .Y(_8324_)
);

AND2X2 _18510_ (
    .A(_7916_),
    .B(_7911_),
    .Y(_8325_)
);

AOI21X1 _18511_ (
    .A(_8319_),
    .B(_8320_),
    .C(_8322_),
    .Y(_8327_)
);

NOR3X1 _18512_ (
    .A(_8314_),
    .B(_8317_),
    .C(_8310_),
    .Y(_8328_)
);

OAI21X1 _18513_ (
    .A(_8328_),
    .B(_8327_),
    .C(_8325_),
    .Y(_8329_)
);

NAND2X1 _18514_ (
    .A(_8324_),
    .B(_8329_),
    .Y(_8330_)
);

AOI21X1 _18515_ (
    .A(_7983_),
    .B(_7982_),
    .C(_7957_),
    .Y(_8331_)
);

OAI21X1 _18516_ (
    .A(_8331_),
    .B(_7955_),
    .C(_7988_),
    .Y(_8332_)
);

NAND2X1 _18517_ (
    .A(breg_7_bF$buf0),
    .B(areg_26_bF$buf4),
    .Y(_8333_)
);

OAI21X1 _18518_ (
    .A(_7929_),
    .B(_8333_),
    .C(_7938_),
    .Y(_8334_)
);

NAND2X1 _18519_ (
    .A(breg[8]),
    .B(areg_25_bF$buf3),
    .Y(_8335_)
);

INVX1 _18520_ (
    .A(_8335_),
    .Y(_8336_)
);

AND2X2 _18521_ (
    .A(breg_7_bF$buf5),
    .B(areg_26_bF$buf3),
    .Y(_8338_)
);

AND2X2 _18522_ (
    .A(breg_6_bF$buf0),
    .B(areg_27_bF$buf0),
    .Y(_8339_)
);

NAND2X1 _18523_ (
    .A(_8338_),
    .B(_8339_),
    .Y(_8340_)
);

OAI21X1 _18524_ (
    .A(_5453__bF$buf3),
    .B(_7100__bF$buf2),
    .C(_8333_),
    .Y(_8341_)
);

NAND3X1 _18525_ (
    .A(_8336_),
    .B(_8341_),
    .C(_8340_),
    .Y(_8342_)
);

OAI21X1 _18526_ (
    .A(_4116__bF$buf0),
    .B(_6686__bF$buf0),
    .C(_8339_),
    .Y(_8343_)
);

OAI21X1 _18527_ (
    .A(_5453__bF$buf2),
    .B(_7100__bF$buf1),
    .C(_8338_),
    .Y(_8344_)
);

NAND3X1 _18528_ (
    .A(_8335_),
    .B(_8343_),
    .C(_8344_),
    .Y(_8345_)
);

NAND2X1 _18529_ (
    .A(breg_4_bF$buf4),
    .B(areg_29_bF$buf1),
    .Y(_8346_)
);

OAI22X1 _18530_ (
    .A(_7518_),
    .B(_8346_),
    .C(_7962_),
    .D(_7958_),
    .Y(_8347_)
);

NAND3X1 _18531_ (
    .A(_8347_),
    .B(_8342_),
    .C(_8345_),
    .Y(_8349_)
);

AOI21X1 _18532_ (
    .A(_8343_),
    .B(_8344_),
    .C(_8335_),
    .Y(_8350_)
);

AOI21X1 _18533_ (
    .A(_8341_),
    .B(_8340_),
    .C(_8336_),
    .Y(_8351_)
);

INVX1 _18534_ (
    .A(_8347_),
    .Y(_8352_)
);

OAI21X1 _18535_ (
    .A(_8350_),
    .B(_8351_),
    .C(_8352_),
    .Y(_8353_)
);

NAND3X1 _18536_ (
    .A(_8334_),
    .B(_8349_),
    .C(_8353_),
    .Y(_8354_)
);

AOI21X1 _18537_ (
    .A(_7490_),
    .B(_8338_),
    .C(_7945_),
    .Y(_8355_)
);

NOR3X1 _18538_ (
    .A(_8351_),
    .B(_8352_),
    .C(_8350_),
    .Y(_8356_)
);

AOI21X1 _18539_ (
    .A(_8342_),
    .B(_8345_),
    .C(_8347_),
    .Y(_8357_)
);

OAI21X1 _18540_ (
    .A(_8356_),
    .B(_8357_),
    .C(_8355_),
    .Y(_8358_)
);

NAND2X1 _18541_ (
    .A(_8354_),
    .B(_8358_),
    .Y(_8360_)
);

NOR2X1 _18542_ (
    .A(_7967_),
    .B(_7111_),
    .Y(_8361_)
);

NAND2X1 _18543_ (
    .A(breg_5_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_8362_)
);

INVX2 _18544_ (
    .A(_8362_),
    .Y(_8363_)
);

NAND2X1 _18545_ (
    .A(breg_3_bF$buf0),
    .B(areg_30_bF$buf4),
    .Y(_8364_)
);

NOR2X1 _18546_ (
    .A(_8364_),
    .B(_7961_),
    .Y(_8365_)
);

AOI21X1 _18547_ (
    .A(breg_3_bF$buf5),
    .B(areg_30_bF$buf3),
    .C(_8346_),
    .Y(_8366_)
);

OAI21X1 _18548_ (
    .A(_8365_),
    .B(_8366_),
    .C(_8363_),
    .Y(_8367_)
);

NAND2X1 _18549_ (
    .A(breg_3_bF$buf4),
    .B(areg_29_bF$buf0),
    .Y(_8368_)
);

NAND2X1 _18550_ (
    .A(breg_4_bF$buf3),
    .B(areg_30_bF$buf2),
    .Y(_8369_)
);

NOR2X1 _18551_ (
    .A(_8368_),
    .B(_8369_),
    .Y(_8371_)
);

AND2X2 _18552_ (
    .A(_8346_),
    .B(_8364_),
    .Y(_8372_)
);

OAI21X1 _18553_ (
    .A(_8372_),
    .B(_8371_),
    .C(_8362_),
    .Y(_8373_)
);

NAND3X1 _18554_ (
    .A(_8361_),
    .B(_8373_),
    .C(_8367_),
    .Y(_8374_)
);

INVX1 _18555_ (
    .A(_8361_),
    .Y(_8375_)
);

OAI21X1 _18556_ (
    .A(_8365_),
    .B(_8366_),
    .C(_8362_),
    .Y(_8376_)
);

OAI21X1 _18557_ (
    .A(_8372_),
    .B(_8371_),
    .C(_8363_),
    .Y(_8377_)
);

NAND3X1 _18558_ (
    .A(_8375_),
    .B(_8377_),
    .C(_8376_),
    .Y(_8378_)
);

NAND2X1 _18559_ (
    .A(_8374_),
    .B(_8378_),
    .Y(_8379_)
);

OAI21X1 _18560_ (
    .A(_7973_),
    .B(_7971_),
    .C(_8379_),
    .Y(_8380_)
);

AOI21X1 _18561_ (
    .A(_7974_),
    .B(_7977_),
    .C(_7971_),
    .Y(_8381_)
);

AND2X2 _18562_ (
    .A(_8374_),
    .B(_8378_),
    .Y(_8382_)
);

NAND2X1 _18563_ (
    .A(_8381_),
    .B(_8382_),
    .Y(_8383_)
);

AOI21X1 _18564_ (
    .A(_8383_),
    .B(_8380_),
    .C(_8360_),
    .Y(_8384_)
);

NAND3X1 _18565_ (
    .A(_8355_),
    .B(_8349_),
    .C(_8353_),
    .Y(_8385_)
);

OAI21X1 _18566_ (
    .A(_8356_),
    .B(_8357_),
    .C(_8334_),
    .Y(_8386_)
);

NAND2X1 _18567_ (
    .A(_8385_),
    .B(_8386_),
    .Y(_8387_)
);

OAI21X1 _18568_ (
    .A(_7973_),
    .B(_7971_),
    .C(_8382_),
    .Y(_8388_)
);

NAND2X1 _18569_ (
    .A(_8379_),
    .B(_8381_),
    .Y(_8389_)
);

AOI21X1 _18570_ (
    .A(_8389_),
    .B(_8388_),
    .C(_8387_),
    .Y(_8390_)
);

OAI21X1 _18571_ (
    .A(_8384_),
    .B(_8390_),
    .C(_8332_),
    .Y(_8392_)
);

NOR3X1 _18572_ (
    .A(_7973_),
    .B(_7978_),
    .C(_7981_),
    .Y(_8393_)
);

AOI21X1 _18573_ (
    .A(_7987_),
    .B(_7989_),
    .C(_8393_),
    .Y(_8394_)
);

NAND3X1 _18574_ (
    .A(_8389_),
    .B(_8388_),
    .C(_8387_),
    .Y(_8395_)
);

NOR2X1 _18575_ (
    .A(_8379_),
    .B(_8381_),
    .Y(_8396_)
);

AND2X2 _18576_ (
    .A(_8381_),
    .B(_8379_),
    .Y(_8397_)
);

OAI21X1 _18577_ (
    .A(_8397_),
    .B(_8396_),
    .C(_8360_),
    .Y(_8398_)
);

NAND3X1 _18578_ (
    .A(_8395_),
    .B(_8398_),
    .C(_8394_),
    .Y(_8399_)
);

AOI21X1 _18579_ (
    .A(_8392_),
    .B(_8399_),
    .C(_8330_),
    .Y(_8400_)
);

OAI21X1 _18580_ (
    .A(_8328_),
    .B(_8327_),
    .C(_8283_),
    .Y(_8401_)
);

NAND3X1 _18581_ (
    .A(_8323_),
    .B(_8325_),
    .C(_8318_),
    .Y(_8403_)
);

NAND2X1 _18582_ (
    .A(_8403_),
    .B(_8401_),
    .Y(_8404_)
);

NAND3X1 _18583_ (
    .A(_8332_),
    .B(_8398_),
    .C(_8395_),
    .Y(_8405_)
);

OAI21X1 _18584_ (
    .A(_8384_),
    .B(_8390_),
    .C(_8394_),
    .Y(_8406_)
);

AOI21X1 _18585_ (
    .A(_8405_),
    .B(_8406_),
    .C(_8404_),
    .Y(_8407_)
);

OAI21X1 _18586_ (
    .A(_8400_),
    .B(_8407_),
    .C(_8281_),
    .Y(_8408_)
);

NOR3X1 _18587_ (
    .A(_7985_),
    .B(_7990_),
    .C(_7993_),
    .Y(_8409_)
);

AOI21X1 _18588_ (
    .A(_8001_),
    .B(_8003_),
    .C(_8409_),
    .Y(_8410_)
);

NAND3X1 _18589_ (
    .A(_8405_),
    .B(_8406_),
    .C(_8404_),
    .Y(_8411_)
);

NAND3X1 _18590_ (
    .A(_8392_),
    .B(_8399_),
    .C(_8330_),
    .Y(_8412_)
);

NAND3X1 _18591_ (
    .A(_8411_),
    .B(_8412_),
    .C(_8410_),
    .Y(_8414_)
);

AOI21X1 _18592_ (
    .A(_8408_),
    .B(_8414_),
    .C(_8279_),
    .Y(_8415_)
);

OAI21X1 _18593_ (
    .A(_8277_),
    .B(_8276_),
    .C(_8188_),
    .Y(_8416_)
);

NAND3X1 _18594_ (
    .A(_8273_),
    .B(_8275_),
    .C(_8268_),
    .Y(_8417_)
);

NAND2X1 _18595_ (
    .A(_8417_),
    .B(_8416_),
    .Y(_8418_)
);

NAND3X1 _18596_ (
    .A(_8411_),
    .B(_8412_),
    .C(_8281_),
    .Y(_8419_)
);

OAI21X1 _18597_ (
    .A(_8400_),
    .B(_8407_),
    .C(_8410_),
    .Y(_8420_)
);

AOI21X1 _18598_ (
    .A(_8419_),
    .B(_8420_),
    .C(_8418_),
    .Y(_8421_)
);

OAI21X1 _18599_ (
    .A(_8415_),
    .B(_8421_),
    .C(_8187_),
    .Y(_8422_)
);

NOR3X1 _18600_ (
    .A(_7998_),
    .B(_8004_),
    .C(_8007_),
    .Y(_8423_)
);

AOI21X1 _18601_ (
    .A(_8015_),
    .B(_8017_),
    .C(_8423_),
    .Y(_8425_)
);

NAND3X1 _18602_ (
    .A(_8419_),
    .B(_8420_),
    .C(_8418_),
    .Y(_8426_)
);

NAND3X1 _18603_ (
    .A(_8408_),
    .B(_8414_),
    .C(_8279_),
    .Y(_8427_)
);

NAND3X1 _18604_ (
    .A(_8426_),
    .B(_8427_),
    .C(_8425_),
    .Y(_8428_)
);

AOI21X1 _18605_ (
    .A(_8422_),
    .B(_8428_),
    .C(_8185_),
    .Y(_8429_)
);

NAND3X1 _18606_ (
    .A(_8174_),
    .B(_8180_),
    .C(_8178_),
    .Y(_8430_)
);

NAND3X1 _18607_ (
    .A(_8079_),
    .B(_8181_),
    .C(_8182_),
    .Y(_8431_)
);

NAND2X1 _18608_ (
    .A(_8431_),
    .B(_8430_),
    .Y(_8432_)
);

NAND3X1 _18609_ (
    .A(_8426_),
    .B(_8427_),
    .C(_8187_),
    .Y(_8433_)
);

OAI21X1 _18610_ (
    .A(_8415_),
    .B(_8421_),
    .C(_8425_),
    .Y(_8434_)
);

AOI21X1 _18611_ (
    .A(_8433_),
    .B(_8434_),
    .C(_8432_),
    .Y(_8436_)
);

OAI21X1 _18612_ (
    .A(_8429_),
    .B(_8436_),
    .C(_8078_),
    .Y(_8437_)
);

NOR3X1 _18613_ (
    .A(_8012_),
    .B(_8018_),
    .C(_8021_),
    .Y(_8438_)
);

AOI21X1 _18614_ (
    .A(_8028_),
    .B(_8031_),
    .C(_8438_),
    .Y(_8439_)
);

NAND3X1 _18615_ (
    .A(_8433_),
    .B(_8434_),
    .C(_8432_),
    .Y(_8440_)
);

NAND3X1 _18616_ (
    .A(_8422_),
    .B(_8428_),
    .C(_8185_),
    .Y(_8441_)
);

NAND3X1 _18617_ (
    .A(_8440_),
    .B(_8441_),
    .C(_8439_),
    .Y(_8442_)
);

AOI21X1 _18618_ (
    .A(_8437_),
    .B(_8442_),
    .C(_8076_),
    .Y(_8443_)
);

NAND3X1 _18619_ (
    .A(_8440_),
    .B(_8441_),
    .C(_8078_),
    .Y(_8444_)
);

OAI21X1 _18620_ (
    .A(_8429_),
    .B(_8436_),
    .C(_8439_),
    .Y(_8445_)
);

AOI21X1 _18621_ (
    .A(_8444_),
    .B(_8445_),
    .C(_8075_),
    .Y(_8447_)
);

OAI21X1 _18622_ (
    .A(_8443_),
    .B(_8447_),
    .C(_8074_),
    .Y(_8448_)
);

AOI21X1 _18623_ (
    .A(_7660_),
    .B(_8043_),
    .C(_8049_),
    .Y(_8449_)
);

NAND3X1 _18624_ (
    .A(_8075_),
    .B(_8444_),
    .C(_8445_),
    .Y(_8450_)
);

NAND3X1 _18625_ (
    .A(_8076_),
    .B(_8437_),
    .C(_8442_),
    .Y(_8451_)
);

NAND3X1 _18626_ (
    .A(_8450_),
    .B(_8451_),
    .C(_8449_),
    .Y(_8452_)
);

AOI21X1 _18627_ (
    .A(_8448_),
    .B(_8452_),
    .C(_8072_),
    .Y(_8453_)
);

NAND3X1 _18628_ (
    .A(_8450_),
    .B(_8451_),
    .C(_8074_),
    .Y(_8454_)
);

OAI21X1 _18629_ (
    .A(_8443_),
    .B(_8447_),
    .C(_8449_),
    .Y(_8455_)
);

AOI21X1 _18630_ (
    .A(_8454_),
    .B(_8455_),
    .C(_8071_),
    .Y(_8456_)
);

OAI21X1 _18631_ (
    .A(_8453_),
    .B(_8456_),
    .C(_8070_),
    .Y(_8458_)
);

AOI21X1 _18632_ (
    .A(_7655_),
    .B(_8056_),
    .C(_8062_),
    .Y(_8459_)
);

NAND3X1 _18633_ (
    .A(_8071_),
    .B(_8454_),
    .C(_8455_),
    .Y(_8460_)
);

NAND3X1 _18634_ (
    .A(_8072_),
    .B(_8448_),
    .C(_8452_),
    .Y(_8461_)
);

NAND3X1 _18635_ (
    .A(_8460_),
    .B(_8461_),
    .C(_8459_),
    .Y(_8462_)
);

NAND2X1 _18636_ (
    .A(_8458_),
    .B(_8462_),
    .Y(_8463_)
);

XNOR2X1 _18637_ (
    .A(_8069_),
    .B(_8463_),
    .Y(_0_[33])
);

NAND3X1 _18638_ (
    .A(_7654_),
    .B(_8061_),
    .C(_8065_),
    .Y(_8464_)
);

NAND3X1 _18639_ (
    .A(_8460_),
    .B(_8461_),
    .C(_8070_),
    .Y(_8465_)
);

OAI21X1 _18640_ (
    .A(_8453_),
    .B(_8456_),
    .C(_8459_),
    .Y(_8466_)
);

INVX1 _18641_ (
    .A(_8466_),
    .Y(_8468_)
);

AOI21X1 _18642_ (
    .A(_8464_),
    .B(_8465_),
    .C(_8468_),
    .Y(_8469_)
);

AOI22X1 _18643_ (
    .A(_8458_),
    .B(_8462_),
    .C(_8058_),
    .D(_8066_),
    .Y(_8470_)
);

AOI21X1 _18644_ (
    .A(_8470_),
    .B(_7652_),
    .C(_8469_),
    .Y(_8471_)
);

AOI21X1 _18645_ (
    .A(_8450_),
    .B(_8451_),
    .C(_8074_),
    .Y(_8472_)
);

OAI21X1 _18646_ (
    .A(_8472_),
    .B(_8072_),
    .C(_8454_),
    .Y(_8473_)
);

OAI21X1 _18647_ (
    .A(_8111_),
    .B(_8081_),
    .C(_8119_),
    .Y(_8474_)
);

INVX2 _18648_ (
    .A(_8474_),
    .Y(_8475_)
);

AOI21X1 _18649_ (
    .A(_8440_),
    .B(_8441_),
    .C(_8078_),
    .Y(_8476_)
);

OAI21X1 _18650_ (
    .A(_8476_),
    .B(_8076_),
    .C(_8444_),
    .Y(_8477_)
);

NAND2X1 _18651_ (
    .A(_8174_),
    .B(_8179_),
    .Y(_8479_)
);

INVX2 _18652_ (
    .A(_8479_),
    .Y(_8480_)
);

AOI21X1 _18653_ (
    .A(_8426_),
    .B(_8427_),
    .C(_8187_),
    .Y(_8481_)
);

OAI21X1 _18654_ (
    .A(_8185_),
    .B(_8481_),
    .C(_8433_),
    .Y(_8482_)
);

NAND2X1 _18655_ (
    .A(_8162_),
    .B(_8167_),
    .Y(_8483_)
);

NOR2X1 _18656_ (
    .A(_2792_),
    .B(_7225__bF$buf1),
    .Y(_8484_)
);

INVX1 _18657_ (
    .A(_8484_),
    .Y(_8485_)
);

OAI21X1 _18658_ (
    .A(_8099_),
    .B(_8085_),
    .C(_8109_),
    .Y(_8486_)
);

NOR2X1 _18659_ (
    .A(_2562__bF$buf0),
    .B(_6815__bF$buf0),
    .Y(_8487_)
);

INVX2 _18660_ (
    .A(_8487_),
    .Y(_8488_)
);

OAI21X1 _18661_ (
    .A(_8097_),
    .B(_8087_),
    .C(_8091_),
    .Y(_8490_)
);

NAND2X1 _18662_ (
    .A(areg_5_bF$buf1),
    .B(breg_29_bF$buf4),
    .Y(_8491_)
);

INVX2 _18663_ (
    .A(_8491_),
    .Y(_8492_)
);

AND2X2 _18664_ (
    .A(areg_6_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_8493_)
);

AND2X2 _18665_ (
    .A(areg_7_bF$buf4),
    .B(breg_27_bF$buf3),
    .Y(_8494_)
);

NAND2X1 _18666_ (
    .A(_8493_),
    .B(_8494_),
    .Y(_8495_)
);

OAI21X1 _18667_ (
    .A(_4434__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_8094_),
    .Y(_8496_)
);

NAND3X1 _18668_ (
    .A(_8492_),
    .B(_8496_),
    .C(_8495_),
    .Y(_8497_)
);

NAND2X1 _18669_ (
    .A(areg_7_bF$buf3),
    .B(breg_27_bF$buf2),
    .Y(_8498_)
);

NOR2X1 _18670_ (
    .A(_8094_),
    .B(_8498_),
    .Y(_8499_)
);

NOR2X1 _18671_ (
    .A(_8493_),
    .B(_8494_),
    .Y(_8501_)
);

OAI21X1 _18672_ (
    .A(_8501_),
    .B(_8499_),
    .C(_8491_),
    .Y(_8502_)
);

AOI21X1 _18673_ (
    .A(_8497_),
    .B(_8502_),
    .C(_8490_),
    .Y(_8503_)
);

AOI21X1 _18674_ (
    .A(_8088_),
    .B(_8092_),
    .C(_8096_),
    .Y(_8504_)
);

OAI21X1 _18675_ (
    .A(_3646__bF$buf2),
    .B(_6050__bF$buf1),
    .C(_8494_),
    .Y(_8505_)
);

OAI21X1 _18676_ (
    .A(_4434__bF$buf1),
    .B(_5668__bF$buf1),
    .C(_8493_),
    .Y(_8506_)
);

AOI21X1 _18677_ (
    .A(_8505_),
    .B(_8506_),
    .C(_8491_),
    .Y(_8507_)
);

AOI21X1 _18678_ (
    .A(_8496_),
    .B(_8495_),
    .C(_8492_),
    .Y(_8508_)
);

NOR3X1 _18679_ (
    .A(_8508_),
    .B(_8504_),
    .C(_8507_),
    .Y(_8509_)
);

OAI21X1 _18680_ (
    .A(_8509_),
    .B(_8503_),
    .C(_8488_),
    .Y(_8510_)
);

OAI21X1 _18681_ (
    .A(_8507_),
    .B(_8508_),
    .C(_8504_),
    .Y(_8512_)
);

NAND3X1 _18682_ (
    .A(_8497_),
    .B(_8490_),
    .C(_8502_),
    .Y(_8513_)
);

NAND3X1 _18683_ (
    .A(_8487_),
    .B(_8512_),
    .C(_8513_),
    .Y(_8514_)
);

AOI21X1 _18684_ (
    .A(_8514_),
    .B(_8510_),
    .C(_8486_),
    .Y(_8515_)
);

AOI21X1 _18685_ (
    .A(_8083_),
    .B(_8108_),
    .C(_8105_),
    .Y(_8516_)
);

AOI21X1 _18686_ (
    .A(_8512_),
    .B(_8513_),
    .C(_8487_),
    .Y(_8517_)
);

NOR3X1 _18687_ (
    .A(_8503_),
    .B(_8488_),
    .C(_8509_),
    .Y(_8518_)
);

NOR3X1 _18688_ (
    .A(_8516_),
    .B(_8517_),
    .C(_8518_),
    .Y(_8519_)
);

OAI21X1 _18689_ (
    .A(_8519_),
    .B(_8515_),
    .C(_8485_),
    .Y(_8520_)
);

OAI21X1 _18690_ (
    .A(_8518_),
    .B(_8517_),
    .C(_8516_),
    .Y(_8521_)
);

NAND3X1 _18691_ (
    .A(_8486_),
    .B(_8514_),
    .C(_8510_),
    .Y(_8523_)
);

NAND3X1 _18692_ (
    .A(_8484_),
    .B(_8523_),
    .C(_8521_),
    .Y(_8524_)
);

AND2X2 _18693_ (
    .A(_8520_),
    .B(_8524_),
    .Y(_8525_)
);

AOI21X1 _18694_ (
    .A(_8148_),
    .B(_8144_),
    .C(_8149_),
    .Y(_8526_)
);

OAI21X1 _18695_ (
    .A(_8526_),
    .B(_8157_),
    .C(_8151_),
    .Y(_8527_)
);

NAND2X1 _18696_ (
    .A(_8140_),
    .B(_8144_),
    .Y(_8528_)
);

OAI21X1 _18697_ (
    .A(_8130_),
    .B(_8125_),
    .C(_8133_),
    .Y(_8529_)
);

NAND2X1 _18698_ (
    .A(areg_8_bF$buf4),
    .B(breg_26_bF$buf1),
    .Y(_8530_)
);

NAND2X1 _18699_ (
    .A(areg_9_bF$buf4),
    .B(breg_25_bF$buf3),
    .Y(_8531_)
);

NAND2X1 _18700_ (
    .A(areg_10_bF$buf3),
    .B(breg_24_bF$buf4),
    .Y(_8532_)
);

NOR2X1 _18701_ (
    .A(_8531_),
    .B(_8532_),
    .Y(_8534_)
);

AND2X2 _18702_ (
    .A(_8531_),
    .B(_8532_),
    .Y(_8535_)
);

OAI21X1 _18703_ (
    .A(_8535_),
    .B(_8534_),
    .C(_8530_),
    .Y(_8536_)
);

INVX1 _18704_ (
    .A(_8530_),
    .Y(_8537_)
);

OR2X2 _18705_ (
    .A(_8531_),
    .B(_8532_),
    .Y(_8538_)
);

OAI21X1 _18706_ (
    .A(_7711__bF$buf0),
    .B(_5315__bF$buf4),
    .C(_8531_),
    .Y(_8539_)
);

NAND3X1 _18707_ (
    .A(_8537_),
    .B(_8539_),
    .C(_8538_),
    .Y(_8540_)
);

NAND2X1 _18708_ (
    .A(areg_12_bF$buf3),
    .B(breg_22_bF$buf2),
    .Y(_8541_)
);

AND2X2 _18709_ (
    .A(_8191_),
    .B(_8192_),
    .Y(_8542_)
);

OAI22X1 _18710_ (
    .A(_7786_),
    .B(_8541_),
    .C(_8542_),
    .D(_8189_),
    .Y(_8543_)
);

NAND3X1 _18711_ (
    .A(_8536_),
    .B(_8540_),
    .C(_8543_),
    .Y(_8545_)
);

AOI21X1 _18712_ (
    .A(_8539_),
    .B(_8538_),
    .C(_8537_),
    .Y(_8546_)
);

NOR3X1 _18713_ (
    .A(_8530_),
    .B(_8534_),
    .C(_8535_),
    .Y(_8547_)
);

NOR2X1 _18714_ (
    .A(_8191_),
    .B(_8192_),
    .Y(_8548_)
);

OAI21X1 _18715_ (
    .A(_10869__bF$buf0),
    .B(_3781__bF$buf1),
    .C(_8191_),
    .Y(_8549_)
);

AOI21X1 _18716_ (
    .A(_8190_),
    .B(_8549_),
    .C(_8548_),
    .Y(_8550_)
);

OAI21X1 _18717_ (
    .A(_8547_),
    .B(_8546_),
    .C(_8550_),
    .Y(_8551_)
);

NAND3X1 _18718_ (
    .A(_8529_),
    .B(_8545_),
    .C(_8551_),
    .Y(_8552_)
);

INVX1 _18719_ (
    .A(_8529_),
    .Y(_8553_)
);

NAND3X1 _18720_ (
    .A(_8550_),
    .B(_8536_),
    .C(_8540_),
    .Y(_8554_)
);

OAI21X1 _18721_ (
    .A(_8547_),
    .B(_8546_),
    .C(_8543_),
    .Y(_8556_)
);

NAND3X1 _18722_ (
    .A(_8553_),
    .B(_8554_),
    .C(_8556_),
    .Y(_8557_)
);

AOI21X1 _18723_ (
    .A(_8210_),
    .B(_8214_),
    .C(_8196_),
    .Y(_8558_)
);

OAI21X1 _18724_ (
    .A(_8195_),
    .B(_8558_),
    .C(_8219_),
    .Y(_8559_)
);

NAND3X1 _18725_ (
    .A(_8552_),
    .B(_8557_),
    .C(_8559_),
    .Y(_8560_)
);

AOI21X1 _18726_ (
    .A(_8554_),
    .B(_8556_),
    .C(_8553_),
    .Y(_8561_)
);

AOI21X1 _18727_ (
    .A(_8545_),
    .B(_8551_),
    .C(_8529_),
    .Y(_8562_)
);

NOR3X1 _18728_ (
    .A(_8207_),
    .B(_8209_),
    .C(_8202_),
    .Y(_8563_)
);

AOI21X1 _18729_ (
    .A(_8220_),
    .B(_8218_),
    .C(_8563_),
    .Y(_8564_)
);

OAI21X1 _18730_ (
    .A(_8562_),
    .B(_8561_),
    .C(_8564_),
    .Y(_8565_)
);

NAND3X1 _18731_ (
    .A(_8528_),
    .B(_8565_),
    .C(_8560_),
    .Y(_8567_)
);

AND2X2 _18732_ (
    .A(_8144_),
    .B(_8140_),
    .Y(_8568_)
);

NOR3X1 _18733_ (
    .A(_8562_),
    .B(_8561_),
    .C(_8564_),
    .Y(_8569_)
);

AOI21X1 _18734_ (
    .A(_8552_),
    .B(_8557_),
    .C(_8559_),
    .Y(_8570_)
);

OAI21X1 _18735_ (
    .A(_8569_),
    .B(_8570_),
    .C(_8568_),
    .Y(_8571_)
);

NAND3X1 _18736_ (
    .A(_8527_),
    .B(_8567_),
    .C(_8571_),
    .Y(_8572_)
);

NOR3X1 _18737_ (
    .A(_8153_),
    .B(_8152_),
    .C(_8154_),
    .Y(_8573_)
);

AOI21X1 _18738_ (
    .A(_8123_),
    .B(_8155_),
    .C(_8573_),
    .Y(_8574_)
);

NAND3X1 _18739_ (
    .A(_8552_),
    .B(_8557_),
    .C(_8564_),
    .Y(_8575_)
);

OAI21X1 _18740_ (
    .A(_8562_),
    .B(_8561_),
    .C(_8559_),
    .Y(_8576_)
);

AOI21X1 _18741_ (
    .A(_8576_),
    .B(_8575_),
    .C(_8568_),
    .Y(_8578_)
);

AOI21X1 _18742_ (
    .A(_8565_),
    .B(_8560_),
    .C(_8528_),
    .Y(_8579_)
);

OAI21X1 _18743_ (
    .A(_8578_),
    .B(_8579_),
    .C(_8574_),
    .Y(_8580_)
);

NAND3X1 _18744_ (
    .A(_8572_),
    .B(_8580_),
    .C(_8525_),
    .Y(_8581_)
);

NAND2X1 _18745_ (
    .A(_8524_),
    .B(_8520_),
    .Y(_8582_)
);

OAI21X1 _18746_ (
    .A(_8578_),
    .B(_8579_),
    .C(_8527_),
    .Y(_8583_)
);

NAND3X1 _18747_ (
    .A(_8567_),
    .B(_8571_),
    .C(_8574_),
    .Y(_8584_)
);

NAND3X1 _18748_ (
    .A(_8582_),
    .B(_8583_),
    .C(_8584_),
    .Y(_8585_)
);

OAI21X1 _18749_ (
    .A(_8276_),
    .B(_8275_),
    .C(_8273_),
    .Y(_8586_)
);

NAND3X1 _18750_ (
    .A(_8586_),
    .B(_8585_),
    .C(_8581_),
    .Y(_8587_)
);

AOI21X1 _18751_ (
    .A(_8583_),
    .B(_8584_),
    .C(_8582_),
    .Y(_8589_)
);

AOI21X1 _18752_ (
    .A(_8572_),
    .B(_8580_),
    .C(_8525_),
    .Y(_8590_)
);

AOI21X1 _18753_ (
    .A(_8188_),
    .B(_8268_),
    .C(_8277_),
    .Y(_8591_)
);

OAI21X1 _18754_ (
    .A(_8589_),
    .B(_8590_),
    .C(_8591_),
    .Y(_8592_)
);

NAND3X1 _18755_ (
    .A(_8483_),
    .B(_8587_),
    .C(_8592_),
    .Y(_8593_)
);

AND2X2 _18756_ (
    .A(_8167_),
    .B(_8162_),
    .Y(_8594_)
);

NAND3X1 _18757_ (
    .A(_8591_),
    .B(_8585_),
    .C(_8581_),
    .Y(_8595_)
);

OAI21X1 _18758_ (
    .A(_8589_),
    .B(_8590_),
    .C(_8586_),
    .Y(_8596_)
);

NAND3X1 _18759_ (
    .A(_8595_),
    .B(_8594_),
    .C(_8596_),
    .Y(_8597_)
);

NAND2X1 _18760_ (
    .A(_8593_),
    .B(_8597_),
    .Y(_8598_)
);

AOI21X1 _18761_ (
    .A(_8411_),
    .B(_8412_),
    .C(_8281_),
    .Y(_8600_)
);

OAI21X1 _18762_ (
    .A(_8279_),
    .B(_8600_),
    .C(_8419_),
    .Y(_8601_)
);

NAND2X1 _18763_ (
    .A(_8264_),
    .B(_8269_),
    .Y(_8602_)
);

NAND2X1 _18764_ (
    .A(areg_11_bF$buf3),
    .B(breg_23_bF$buf2),
    .Y(_8603_)
);

INVX2 _18765_ (
    .A(_8603_),
    .Y(_8604_)
);

NAND2X1 _18766_ (
    .A(areg_13_bF$buf1),
    .B(breg_21_bF$buf2),
    .Y(_8605_)
);

XOR2X1 _18767_ (
    .A(_8541_),
    .B(_8605_),
    .Y(_8606_)
);

XNOR2X1 _18768_ (
    .A(_8606_),
    .B(_8604_),
    .Y(_8607_)
);

OAI21X1 _18769_ (
    .A(_8213_),
    .B(_8197_),
    .C(_8204_),
    .Y(_8608_)
);

NOR2X1 _18770_ (
    .A(_2287__bF$buf1),
    .B(_3526_),
    .Y(_8609_)
);

INVX2 _18771_ (
    .A(_8609_),
    .Y(_8611_)
);

AND2X2 _18772_ (
    .A(areg_16_bF$buf2),
    .B(breg_18_bF$buf2),
    .Y(_8612_)
);

OAI21X1 _18773_ (
    .A(_2465__bF$buf2),
    .B(_3253__bF$buf3),
    .C(_8612_),
    .Y(_8613_)
);

AND2X2 _18774_ (
    .A(areg_15_bF$buf4),
    .B(breg_19_bF$buf3),
    .Y(_8614_)
);

OAI21X1 _18775_ (
    .A(_2669__bF$buf3),
    .B(_3529__bF$buf3),
    .C(_8614_),
    .Y(_8615_)
);

AOI21X1 _18776_ (
    .A(_8613_),
    .B(_8615_),
    .C(_8611_),
    .Y(_8616_)
);

NAND2X1 _18777_ (
    .A(_8614_),
    .B(_8612_),
    .Y(_8617_)
);

OAI22X1 _18778_ (
    .A(_2465__bF$buf1),
    .B(_3253__bF$buf2),
    .C(_2669__bF$buf2),
    .D(_3529__bF$buf2),
    .Y(_8618_)
);

AOI21X1 _18779_ (
    .A(_8618_),
    .B(_8617_),
    .C(_8609_),
    .Y(_8619_)
);

OAI21X1 _18780_ (
    .A(_8616_),
    .B(_8619_),
    .C(_8608_),
    .Y(_8620_)
);

AOI21X1 _18781_ (
    .A(_8203_),
    .B(_8206_),
    .C(_8212_),
    .Y(_8622_)
);

NAND3X1 _18782_ (
    .A(_8609_),
    .B(_8618_),
    .C(_8617_),
    .Y(_8623_)
);

NAND2X1 _18783_ (
    .A(areg_16_bF$buf1),
    .B(breg_19_bF$buf2),
    .Y(_8624_)
);

NOR2X1 _18784_ (
    .A(_8211_),
    .B(_8624_),
    .Y(_8625_)
);

NOR2X1 _18785_ (
    .A(_8614_),
    .B(_8612_),
    .Y(_8626_)
);

OAI21X1 _18786_ (
    .A(_8626_),
    .B(_8625_),
    .C(_8611_),
    .Y(_8627_)
);

NAND3X1 _18787_ (
    .A(_8622_),
    .B(_8623_),
    .C(_8627_),
    .Y(_8628_)
);

AOI21X1 _18788_ (
    .A(_8628_),
    .B(_8620_),
    .C(_8607_),
    .Y(_8629_)
);

XNOR2X1 _18789_ (
    .A(_8606_),
    .B(_8603_),
    .Y(_8630_)
);

NAND3X1 _18790_ (
    .A(_8623_),
    .B(_8608_),
    .C(_8627_),
    .Y(_8631_)
);

OAI21X1 _18791_ (
    .A(_8616_),
    .B(_8619_),
    .C(_8622_),
    .Y(_8633_)
);

AOI21X1 _18792_ (
    .A(_8631_),
    .B(_8633_),
    .C(_8630_),
    .Y(_8634_)
);

OR2X2 _18793_ (
    .A(_8629_),
    .B(_8634_),
    .Y(_8635_)
);

OAI21X1 _18794_ (
    .A(_8258_),
    .B(_8225_),
    .C(_8251_),
    .Y(_8636_)
);

AND2X2 _18795_ (
    .A(breg_16_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_8637_)
);

AOI21X1 _18796_ (
    .A(_7823_),
    .B(_8637_),
    .C(_8241_),
    .Y(_8638_)
);

NAND2X1 _18797_ (
    .A(areg_17_bF$buf2),
    .B(breg_17_bF$buf1),
    .Y(_8639_)
);

INVX1 _18798_ (
    .A(_8639_),
    .Y(_8640_)
);

AND2X2 _18799_ (
    .A(breg_15_bF$buf2),
    .B(areg_19_bF$buf4),
    .Y(_8641_)
);

NAND2X1 _18800_ (
    .A(_8637_),
    .B(_8641_),
    .Y(_8642_)
);

NAND2X1 _18801_ (
    .A(breg_16_bF$buf2),
    .B(areg_18_bF$buf2),
    .Y(_8644_)
);

OAI21X1 _18802_ (
    .A(_2362__bF$buf0),
    .B(_3402__bF$buf1),
    .C(_8644_),
    .Y(_8645_)
);

NAND3X1 _18803_ (
    .A(_8640_),
    .B(_8645_),
    .C(_8642_),
    .Y(_8646_)
);

OAI21X1 _18804_ (
    .A(_2560__bF$buf2),
    .B(_3146__bF$buf2),
    .C(_8641_),
    .Y(_8647_)
);

OAI21X1 _18805_ (
    .A(_2362__bF$buf5),
    .B(_3402__bF$buf0),
    .C(_8637_),
    .Y(_8648_)
);

NAND3X1 _18806_ (
    .A(_8639_),
    .B(_8647_),
    .C(_8648_),
    .Y(_8649_)
);

NOR2X1 _18807_ (
    .A(_8243_),
    .B(_8286_),
    .Y(_8650_)
);

OAI21X1 _18808_ (
    .A(_2586__bF$buf2),
    .B(_3961__bF$buf4),
    .C(_8243_),
    .Y(_8651_)
);

AOI21X1 _18809_ (
    .A(_8285_),
    .B(_8651_),
    .C(_8650_),
    .Y(_8652_)
);

NAND3X1 _18810_ (
    .A(_8652_),
    .B(_8646_),
    .C(_8649_),
    .Y(_8653_)
);

AOI21X1 _18811_ (
    .A(_8647_),
    .B(_8648_),
    .C(_8639_),
    .Y(_8655_)
);

AOI21X1 _18812_ (
    .A(_8645_),
    .B(_8642_),
    .C(_8640_),
    .Y(_8656_)
);

NAND2X1 _18813_ (
    .A(breg_13_bF$buf3),
    .B(areg_21_bF$buf3),
    .Y(_8657_)
);

AND2X2 _18814_ (
    .A(_8243_),
    .B(_8286_),
    .Y(_8658_)
);

OAI22X1 _18815_ (
    .A(_7884_),
    .B(_8657_),
    .C(_8658_),
    .D(_8284_),
    .Y(_8659_)
);

OAI21X1 _18816_ (
    .A(_8655_),
    .B(_8656_),
    .C(_8659_),
    .Y(_8660_)
);

AOI21X1 _18817_ (
    .A(_8653_),
    .B(_8660_),
    .C(_8638_),
    .Y(_8661_)
);

OAI21X1 _18818_ (
    .A(_8248_),
    .B(_8644_),
    .C(_8232_),
    .Y(_8662_)
);

NAND3X1 _18819_ (
    .A(_8646_),
    .B(_8649_),
    .C(_8659_),
    .Y(_8663_)
);

OAI21X1 _18820_ (
    .A(_8655_),
    .B(_8656_),
    .C(_8652_),
    .Y(_8664_)
);

AOI21X1 _18821_ (
    .A(_8663_),
    .B(_8664_),
    .C(_8662_),
    .Y(_8666_)
);

OAI21X1 _18822_ (
    .A(_8661_),
    .B(_8666_),
    .C(_8636_),
    .Y(_8667_)
);

AOI21X1 _18823_ (
    .A(_8250_),
    .B(_8252_),
    .C(_8257_),
    .Y(_8668_)
);

NAND3X1 _18824_ (
    .A(_8662_),
    .B(_8663_),
    .C(_8664_),
    .Y(_8669_)
);

NOR3X1 _18825_ (
    .A(_8656_),
    .B(_8652_),
    .C(_8655_),
    .Y(_8670_)
);

AOI21X1 _18826_ (
    .A(_8646_),
    .B(_8649_),
    .C(_8659_),
    .Y(_8671_)
);

OAI21X1 _18827_ (
    .A(_8670_),
    .B(_8671_),
    .C(_8638_),
    .Y(_8672_)
);

NAND3X1 _18828_ (
    .A(_8668_),
    .B(_8669_),
    .C(_8672_),
    .Y(_8673_)
);

AOI21X1 _18829_ (
    .A(_8667_),
    .B(_8673_),
    .C(_8635_),
    .Y(_8674_)
);

NOR2X1 _18830_ (
    .A(_8634_),
    .B(_8629_),
    .Y(_8675_)
);

NAND3X1 _18831_ (
    .A(_8636_),
    .B(_8669_),
    .C(_8672_),
    .Y(_8677_)
);

OAI21X1 _18832_ (
    .A(_8661_),
    .B(_8666_),
    .C(_8668_),
    .Y(_8678_)
);

AOI21X1 _18833_ (
    .A(_8678_),
    .B(_8677_),
    .C(_8675_),
    .Y(_8679_)
);

AOI21X1 _18834_ (
    .A(_8283_),
    .B(_8318_),
    .C(_8328_),
    .Y(_8680_)
);

OAI21X1 _18835_ (
    .A(_8674_),
    .B(_8679_),
    .C(_8680_),
    .Y(_8681_)
);

NAND3X1 _18836_ (
    .A(_8678_),
    .B(_8675_),
    .C(_8677_),
    .Y(_8682_)
);

NAND3X1 _18837_ (
    .A(_8667_),
    .B(_8673_),
    .C(_8635_),
    .Y(_8683_)
);

OAI21X1 _18838_ (
    .A(_8327_),
    .B(_8325_),
    .C(_8323_),
    .Y(_8684_)
);

NAND3X1 _18839_ (
    .A(_8682_),
    .B(_8684_),
    .C(_8683_),
    .Y(_8685_)
);

NAND3X1 _18840_ (
    .A(_8602_),
    .B(_8685_),
    .C(_8681_),
    .Y(_8686_)
);

AND2X2 _18841_ (
    .A(_8269_),
    .B(_8264_),
    .Y(_8688_)
);

AOI21X1 _18842_ (
    .A(_8682_),
    .B(_8683_),
    .C(_8684_),
    .Y(_8689_)
);

NOR3X1 _18843_ (
    .A(_8674_),
    .B(_8679_),
    .C(_8680_),
    .Y(_8690_)
);

OAI21X1 _18844_ (
    .A(_8690_),
    .B(_8689_),
    .C(_8688_),
    .Y(_8691_)
);

NAND2X1 _18845_ (
    .A(_8686_),
    .B(_8691_),
    .Y(_8692_)
);

AOI21X1 _18846_ (
    .A(_8398_),
    .B(_8395_),
    .C(_8332_),
    .Y(_8693_)
);

OAI21X1 _18847_ (
    .A(_8330_),
    .B(_8693_),
    .C(_8405_),
    .Y(_8694_)
);

NAND2X1 _18848_ (
    .A(_8312_),
    .B(_8319_),
    .Y(_8695_)
);

NAND2X1 _18849_ (
    .A(breg_14_bF$buf1),
    .B(areg_20_bF$buf1),
    .Y(_8696_)
);

INVX2 _18850_ (
    .A(_8696_),
    .Y(_8697_)
);

NAND2X1 _18851_ (
    .A(breg_12_bF$buf1),
    .B(areg_22_bF$buf3),
    .Y(_8699_)
);

XOR2X1 _18852_ (
    .A(_8657_),
    .B(_8699_),
    .Y(_8700_)
);

XNOR2X1 _18853_ (
    .A(_8700_),
    .B(_8697_),
    .Y(_8701_)
);

OAI21X1 _18854_ (
    .A(_8307_),
    .B(_8290_),
    .C(_8298_),
    .Y(_8702_)
);

NAND2X1 _18855_ (
    .A(breg_11_bF$buf3),
    .B(areg_23_bF$buf0),
    .Y(_8703_)
);

AND2X2 _18856_ (
    .A(breg_9_bF$buf0),
    .B(areg_25_bF$buf2),
    .Y(_8704_)
);

OAI21X1 _18857_ (
    .A(_7217__bF$buf0),
    .B(_5921__bF$buf1),
    .C(_8704_),
    .Y(_8705_)
);

AND2X2 _18858_ (
    .A(breg_10_bF$buf2),
    .B(areg_24_bF$buf4),
    .Y(_8706_)
);

OAI21X1 _18859_ (
    .A(_6044__bF$buf2),
    .B(_6300__bF$buf2),
    .C(_8706_),
    .Y(_8707_)
);

AOI21X1 _18860_ (
    .A(_8705_),
    .B(_8707_),
    .C(_8703_),
    .Y(_8708_)
);

INVX2 _18861_ (
    .A(_8703_),
    .Y(_8710_)
);

NAND2X1 _18862_ (
    .A(_8706_),
    .B(_8704_),
    .Y(_8711_)
);

OAI21X1 _18863_ (
    .A(_6044__bF$buf1),
    .B(_6300__bF$buf1),
    .C(_8305_),
    .Y(_8712_)
);

AOI21X1 _18864_ (
    .A(_8712_),
    .B(_8711_),
    .C(_8710_),
    .Y(_8713_)
);

OAI21X1 _18865_ (
    .A(_8708_),
    .B(_8713_),
    .C(_8702_),
    .Y(_8714_)
);

AOI21X1 _18866_ (
    .A(_8297_),
    .B(_8299_),
    .C(_8306_),
    .Y(_8715_)
);

NAND3X1 _18867_ (
    .A(_8710_),
    .B(_8712_),
    .C(_8711_),
    .Y(_8716_)
);

NAND2X1 _18868_ (
    .A(breg_9_bF$buf5),
    .B(areg_25_bF$buf1),
    .Y(_8717_)
);

NOR2X1 _18869_ (
    .A(_8305_),
    .B(_8717_),
    .Y(_8718_)
);

NOR2X1 _18870_ (
    .A(_8706_),
    .B(_8704_),
    .Y(_8719_)
);

OAI21X1 _18871_ (
    .A(_8719_),
    .B(_8718_),
    .C(_8703_),
    .Y(_8721_)
);

NAND3X1 _18872_ (
    .A(_8715_),
    .B(_8716_),
    .C(_8721_),
    .Y(_8722_)
);

AOI21X1 _18873_ (
    .A(_8714_),
    .B(_8722_),
    .C(_8701_),
    .Y(_8723_)
);

XNOR2X1 _18874_ (
    .A(_8700_),
    .B(_8696_),
    .Y(_8724_)
);

NAND3X1 _18875_ (
    .A(_8716_),
    .B(_8702_),
    .C(_8721_),
    .Y(_8725_)
);

OAI21X1 _18876_ (
    .A(_8708_),
    .B(_8713_),
    .C(_8715_),
    .Y(_8726_)
);

AOI21X1 _18877_ (
    .A(_8725_),
    .B(_8726_),
    .C(_8724_),
    .Y(_8727_)
);

AOI21X1 _18878_ (
    .A(_8334_),
    .B(_8353_),
    .C(_8356_),
    .Y(_8728_)
);

OAI21X1 _18879_ (
    .A(_8723_),
    .B(_8727_),
    .C(_8728_),
    .Y(_8729_)
);

NAND3X1 _18880_ (
    .A(_8725_),
    .B(_8726_),
    .C(_8724_),
    .Y(_8730_)
);

NAND3X1 _18881_ (
    .A(_8714_),
    .B(_8722_),
    .C(_8701_),
    .Y(_8732_)
);

OAI21X1 _18882_ (
    .A(_8357_),
    .B(_8355_),
    .C(_8349_),
    .Y(_8733_)
);

NAND3X1 _18883_ (
    .A(_8733_),
    .B(_8730_),
    .C(_8732_),
    .Y(_8734_)
);

NAND3X1 _18884_ (
    .A(_8695_),
    .B(_8734_),
    .C(_8729_),
    .Y(_8735_)
);

AND2X2 _18885_ (
    .A(_8319_),
    .B(_8312_),
    .Y(_8736_)
);

AOI21X1 _18886_ (
    .A(_8730_),
    .B(_8732_),
    .C(_8733_),
    .Y(_8737_)
);

NOR3X1 _18887_ (
    .A(_8727_),
    .B(_8728_),
    .C(_8723_),
    .Y(_8738_)
);

OAI21X1 _18888_ (
    .A(_8738_),
    .B(_8737_),
    .C(_8736_),
    .Y(_8739_)
);

NAND2X1 _18889_ (
    .A(_8735_),
    .B(_8739_),
    .Y(_8740_)
);

OAI21X1 _18890_ (
    .A(_8360_),
    .B(_8397_),
    .C(_8388_),
    .Y(_8741_)
);

AND2X2 _18891_ (
    .A(breg_7_bF$buf4),
    .B(areg_27_bF$buf5),
    .Y(_8743_)
);

AOI21X1 _18892_ (
    .A(_7935_),
    .B(_8743_),
    .C(_8350_),
    .Y(_8744_)
);

NAND2X1 _18893_ (
    .A(breg[8]),
    .B(areg_26_bF$buf2),
    .Y(_8745_)
);

INVX1 _18894_ (
    .A(_8745_),
    .Y(_8746_)
);

AND2X2 _18895_ (
    .A(breg_6_bF$buf5),
    .B(areg_28_bF$buf5),
    .Y(_8747_)
);

NAND2X1 _18896_ (
    .A(_8743_),
    .B(_8747_),
    .Y(_8748_)
);

OAI22X1 _18897_ (
    .A(_5453__bF$buf1),
    .B(_7520__bF$buf2),
    .C(_4116__bF$buf4),
    .D(_7100__bF$buf0),
    .Y(_8749_)
);

NAND3X1 _18898_ (
    .A(_8746_),
    .B(_8749_),
    .C(_8748_),
    .Y(_8750_)
);

OAI21X1 _18899_ (
    .A(_4116__bF$buf3),
    .B(_7100__bF$buf3),
    .C(_8747_),
    .Y(_8751_)
);

OAI21X1 _18900_ (
    .A(_5453__bF$buf0),
    .B(_7520__bF$buf1),
    .C(_8743_),
    .Y(_8752_)
);

NAND3X1 _18901_ (
    .A(_8745_),
    .B(_8751_),
    .C(_8752_),
    .Y(_8754_)
);

OAI22X1 _18902_ (
    .A(_8368_),
    .B(_8369_),
    .C(_8372_),
    .D(_8362_),
    .Y(_8755_)
);

NAND3X1 _18903_ (
    .A(_8750_),
    .B(_8754_),
    .C(_8755_),
    .Y(_8756_)
);

AOI21X1 _18904_ (
    .A(_8751_),
    .B(_8752_),
    .C(_8745_),
    .Y(_8757_)
);

AOI21X1 _18905_ (
    .A(_8749_),
    .B(_8748_),
    .C(_8746_),
    .Y(_8758_)
);

INVX4 _18906_ (
    .A(areg_30_bF$buf1),
    .Y(_8759_)
);

OAI21X1 _18907_ (
    .A(_2365_),
    .B(_8759_),
    .C(_8346_),
    .Y(_8760_)
);

AOI21X1 _18908_ (
    .A(_8363_),
    .B(_8760_),
    .C(_8371_),
    .Y(_8761_)
);

OAI21X1 _18909_ (
    .A(_8757_),
    .B(_8758_),
    .C(_8761_),
    .Y(_8762_)
);

NAND3X1 _18910_ (
    .A(_8744_),
    .B(_8756_),
    .C(_8762_),
    .Y(_8763_)
);

INVX1 _18911_ (
    .A(_8339_),
    .Y(_8765_)
);

OAI21X1 _18912_ (
    .A(_8333_),
    .B(_8765_),
    .C(_8342_),
    .Y(_8766_)
);

NOR3X1 _18913_ (
    .A(_8758_),
    .B(_8761_),
    .C(_8757_),
    .Y(_8767_)
);

AOI21X1 _18914_ (
    .A(_8750_),
    .B(_8754_),
    .C(_8755_),
    .Y(_8768_)
);

OAI21X1 _18915_ (
    .A(_8767_),
    .B(_8768_),
    .C(_8766_),
    .Y(_8769_)
);

AOI21X1 _18916_ (
    .A(_8377_),
    .B(_8376_),
    .C(_8375_),
    .Y(_8770_)
);

NAND2X1 _18917_ (
    .A(breg_5_bF$buf3),
    .B(areg_29_bF$buf5),
    .Y(_8771_)
);

NAND2X1 _18918_ (
    .A(breg_4_bF$buf2),
    .B(areg_31_bF$buf3),
    .Y(_8772_)
);

INVX8 _18919_ (
    .A(areg_31_bF$buf2),
    .Y(_8773_)
);

OAI21X1 _18920_ (
    .A(_2365_),
    .B(_8773_),
    .C(_8369_),
    .Y(_8774_)
);

OAI21X1 _18921_ (
    .A(_8364_),
    .B(_8772_),
    .C(_8774_),
    .Y(_8776_)
);

XNOR2X1 _18922_ (
    .A(_8776_),
    .B(_8771_),
    .Y(_8777_)
);

OAI21X1 _18923_ (
    .A(_8770_),
    .B(_7968_),
    .C(_8777_),
    .Y(_8778_)
);

INVX2 _18924_ (
    .A(_7968_),
    .Y(_8779_)
);

INVX2 _18925_ (
    .A(_8771_),
    .Y(_8780_)
);

XNOR2X1 _18926_ (
    .A(_8776_),
    .B(_8780_),
    .Y(_8781_)
);

NAND3X1 _18927_ (
    .A(_8779_),
    .B(_8374_),
    .C(_8781_),
    .Y(_8782_)
);

AOI22X1 _18928_ (
    .A(_8778_),
    .B(_8782_),
    .C(_8769_),
    .D(_8763_),
    .Y(_8783_)
);

NAND3X1 _18929_ (
    .A(_8766_),
    .B(_8756_),
    .C(_8762_),
    .Y(_8784_)
);

OAI21X1 _18930_ (
    .A(_8767_),
    .B(_8768_),
    .C(_8744_),
    .Y(_8785_)
);

OAI21X1 _18931_ (
    .A(_8770_),
    .B(_7968_),
    .C(_8781_),
    .Y(_8787_)
);

NAND3X1 _18932_ (
    .A(_8779_),
    .B(_8374_),
    .C(_8777_),
    .Y(_8788_)
);

AOI22X1 _18933_ (
    .A(_8787_),
    .B(_8788_),
    .C(_8785_),
    .D(_8784_),
    .Y(_8789_)
);

OAI21X1 _18934_ (
    .A(_8783_),
    .B(_8789_),
    .C(_8741_),
    .Y(_8790_)
);

AOI21X1 _18935_ (
    .A(_8389_),
    .B(_8387_),
    .C(_8396_),
    .Y(_8791_)
);

NOR2X1 _18936_ (
    .A(_8783_),
    .B(_8789_),
    .Y(_8792_)
);

NAND2X1 _18937_ (
    .A(_8791_),
    .B(_8792_),
    .Y(_8793_)
);

AOI21X1 _18938_ (
    .A(_8790_),
    .B(_8793_),
    .C(_8740_),
    .Y(_8794_)
);

OAI21X1 _18939_ (
    .A(_8738_),
    .B(_8737_),
    .C(_8695_),
    .Y(_8795_)
);

NAND3X1 _18940_ (
    .A(_8734_),
    .B(_8736_),
    .C(_8729_),
    .Y(_8796_)
);

NAND2X1 _18941_ (
    .A(_8796_),
    .B(_8795_),
    .Y(_8798_)
);

OAI21X1 _18942_ (
    .A(_8384_),
    .B(_8396_),
    .C(_8792_),
    .Y(_8799_)
);

OAI21X1 _18943_ (
    .A(_8783_),
    .B(_8789_),
    .C(_8791_),
    .Y(_8800_)
);

AOI21X1 _18944_ (
    .A(_8799_),
    .B(_8800_),
    .C(_8798_),
    .Y(_8801_)
);

OAI21X1 _18945_ (
    .A(_8794_),
    .B(_8801_),
    .C(_8694_),
    .Y(_8802_)
);

NOR3X1 _18946_ (
    .A(_8384_),
    .B(_8390_),
    .C(_8394_),
    .Y(_8803_)
);

AOI21X1 _18947_ (
    .A(_8406_),
    .B(_8404_),
    .C(_8803_),
    .Y(_8804_)
);

NAND3X1 _18948_ (
    .A(_8799_),
    .B(_8800_),
    .C(_8798_),
    .Y(_8805_)
);

NAND3X1 _18949_ (
    .A(_8761_),
    .B(_8750_),
    .C(_8754_),
    .Y(_8806_)
);

OAI21X1 _18950_ (
    .A(_8757_),
    .B(_8758_),
    .C(_8755_),
    .Y(_8807_)
);

AOI21X1 _18951_ (
    .A(_8806_),
    .B(_8807_),
    .C(_8766_),
    .Y(_8809_)
);

AOI21X1 _18952_ (
    .A(_8756_),
    .B(_8762_),
    .C(_8744_),
    .Y(_8810_)
);

AOI21X1 _18953_ (
    .A(_8779_),
    .B(_8374_),
    .C(_8781_),
    .Y(_8811_)
);

NOR3X1 _18954_ (
    .A(_8770_),
    .B(_7968_),
    .C(_8777_),
    .Y(_8812_)
);

OAI22X1 _18955_ (
    .A(_8809_),
    .B(_8810_),
    .C(_8812_),
    .D(_8811_),
    .Y(_8813_)
);

AOI21X1 _18956_ (
    .A(_8806_),
    .B(_8807_),
    .C(_8744_),
    .Y(_8814_)
);

AOI21X1 _18957_ (
    .A(_8756_),
    .B(_8762_),
    .C(_8766_),
    .Y(_8815_)
);

AOI21X1 _18958_ (
    .A(_8779_),
    .B(_8374_),
    .C(_8777_),
    .Y(_8816_)
);

NOR3X1 _18959_ (
    .A(_8770_),
    .B(_7968_),
    .C(_8781_),
    .Y(_8817_)
);

OAI22X1 _18960_ (
    .A(_8814_),
    .B(_8815_),
    .C(_8817_),
    .D(_8816_),
    .Y(_8818_)
);

NAND2X1 _18961_ (
    .A(_8813_),
    .B(_8818_),
    .Y(_8820_)
);

NOR2X1 _18962_ (
    .A(_8791_),
    .B(_8820_),
    .Y(_8821_)
);

NOR2X1 _18963_ (
    .A(_8741_),
    .B(_8792_),
    .Y(_8822_)
);

OAI21X1 _18964_ (
    .A(_8822_),
    .B(_8821_),
    .C(_8740_),
    .Y(_8823_)
);

NAND3X1 _18965_ (
    .A(_8805_),
    .B(_8823_),
    .C(_8804_),
    .Y(_8824_)
);

AOI21X1 _18966_ (
    .A(_8824_),
    .B(_8802_),
    .C(_8692_),
    .Y(_8825_)
);

OAI21X1 _18967_ (
    .A(_8690_),
    .B(_8689_),
    .C(_8602_),
    .Y(_8826_)
);

NAND3X1 _18968_ (
    .A(_8688_),
    .B(_8685_),
    .C(_8681_),
    .Y(_8827_)
);

NAND2X1 _18969_ (
    .A(_8827_),
    .B(_8826_),
    .Y(_8828_)
);

NAND3X1 _18970_ (
    .A(_8805_),
    .B(_8823_),
    .C(_8694_),
    .Y(_8829_)
);

OAI21X1 _18971_ (
    .A(_8794_),
    .B(_8801_),
    .C(_8804_),
    .Y(_8831_)
);

AOI21X1 _18972_ (
    .A(_8829_),
    .B(_8831_),
    .C(_8828_),
    .Y(_8832_)
);

OAI21X1 _18973_ (
    .A(_8825_),
    .B(_8832_),
    .C(_8601_),
    .Y(_8833_)
);

NOR3X1 _18974_ (
    .A(_8400_),
    .B(_8407_),
    .C(_8410_),
    .Y(_8834_)
);

AOI21X1 _18975_ (
    .A(_8418_),
    .B(_8420_),
    .C(_8834_),
    .Y(_8835_)
);

NAND3X1 _18976_ (
    .A(_8829_),
    .B(_8831_),
    .C(_8828_),
    .Y(_8836_)
);

NAND3X1 _18977_ (
    .A(_8802_),
    .B(_8824_),
    .C(_8692_),
    .Y(_8837_)
);

NAND3X1 _18978_ (
    .A(_8836_),
    .B(_8837_),
    .C(_8835_),
    .Y(_8838_)
);

AOI21X1 _18979_ (
    .A(_8838_),
    .B(_8833_),
    .C(_8598_),
    .Y(_8839_)
);

NAND3X1 _18980_ (
    .A(_8587_),
    .B(_8594_),
    .C(_8592_),
    .Y(_8840_)
);

NAND3X1 _18981_ (
    .A(_8483_),
    .B(_8595_),
    .C(_8596_),
    .Y(_8841_)
);

NAND2X1 _18982_ (
    .A(_8841_),
    .B(_8840_),
    .Y(_8842_)
);

NAND3X1 _18983_ (
    .A(_8836_),
    .B(_8837_),
    .C(_8601_),
    .Y(_8843_)
);

OAI21X1 _18984_ (
    .A(_8825_),
    .B(_8832_),
    .C(_8835_),
    .Y(_8844_)
);

AOI21X1 _18985_ (
    .A(_8843_),
    .B(_8844_),
    .C(_8842_),
    .Y(_8845_)
);

OAI21X1 _18986_ (
    .A(_8839_),
    .B(_8845_),
    .C(_8482_),
    .Y(_8846_)
);

NOR3X1 _18987_ (
    .A(_8415_),
    .B(_8421_),
    .C(_8425_),
    .Y(_8847_)
);

AOI21X1 _18988_ (
    .A(_8432_),
    .B(_8434_),
    .C(_8847_),
    .Y(_8848_)
);

NAND3X1 _18989_ (
    .A(_8843_),
    .B(_8844_),
    .C(_8842_),
    .Y(_8849_)
);

NAND3X1 _18990_ (
    .A(_8838_),
    .B(_8598_),
    .C(_8833_),
    .Y(_8850_)
);

NAND3X1 _18991_ (
    .A(_8849_),
    .B(_8850_),
    .C(_8848_),
    .Y(_8853_)
);

AOI21X1 _18992_ (
    .A(_8853_),
    .B(_8846_),
    .C(_8480_),
    .Y(_8854_)
);

NAND3X1 _18993_ (
    .A(_8849_),
    .B(_8850_),
    .C(_8482_),
    .Y(_8855_)
);

OAI21X1 _18994_ (
    .A(_8839_),
    .B(_8845_),
    .C(_8848_),
    .Y(_8856_)
);

AOI21X1 _18995_ (
    .A(_8855_),
    .B(_8856_),
    .C(_8479_),
    .Y(_8857_)
);

OAI21X1 _18996_ (
    .A(_8854_),
    .B(_8857_),
    .C(_8477_),
    .Y(_8858_)
);

NOR3X1 _18997_ (
    .A(_8429_),
    .B(_8436_),
    .C(_8439_),
    .Y(_8859_)
);

AOI21X1 _18998_ (
    .A(_8075_),
    .B(_8445_),
    .C(_8859_),
    .Y(_8860_)
);

NAND3X1 _18999_ (
    .A(_8479_),
    .B(_8855_),
    .C(_8856_),
    .Y(_8861_)
);

NAND3X1 _19000_ (
    .A(_8480_),
    .B(_8853_),
    .C(_8846_),
    .Y(_8862_)
);

NAND3X1 _19001_ (
    .A(_8861_),
    .B(_8862_),
    .C(_8860_),
    .Y(_8864_)
);

AOI21X1 _19002_ (
    .A(_8864_),
    .B(_8858_),
    .C(_8475_),
    .Y(_8865_)
);

NAND3X1 _19003_ (
    .A(_8861_),
    .B(_8477_),
    .C(_8862_),
    .Y(_8866_)
);

OAI21X1 _19004_ (
    .A(_8854_),
    .B(_8857_),
    .C(_8860_),
    .Y(_8867_)
);

AOI21X1 _19005_ (
    .A(_8866_),
    .B(_8867_),
    .C(_8474_),
    .Y(_8868_)
);

OAI21X1 _19006_ (
    .A(_8865_),
    .B(_8868_),
    .C(_8473_),
    .Y(_8869_)
);

NOR3X1 _19007_ (
    .A(_8443_),
    .B(_8447_),
    .C(_8449_),
    .Y(_8870_)
);

AOI21X1 _19008_ (
    .A(_8071_),
    .B(_8455_),
    .C(_8870_),
    .Y(_8871_)
);

NAND3X1 _19009_ (
    .A(_8474_),
    .B(_8866_),
    .C(_8867_),
    .Y(_8872_)
);

NAND3X1 _19010_ (
    .A(_8475_),
    .B(_8864_),
    .C(_8858_),
    .Y(_8873_)
);

NAND3X1 _19011_ (
    .A(_8872_),
    .B(_8873_),
    .C(_8871_),
    .Y(_8875_)
);

NAND2X1 _19012_ (
    .A(_8875_),
    .B(_8869_),
    .Y(_8876_)
);

XNOR2X1 _19013_ (
    .A(_8471_),
    .B(_8876_),
    .Y(_0_[34])
);

INVX1 _19014_ (
    .A(_8471_),
    .Y(_8877_)
);

NOR3X1 _19015_ (
    .A(_8865_),
    .B(_8868_),
    .C(_8871_),
    .Y(_8878_)
);

AOI21X1 _19016_ (
    .A(_8876_),
    .B(_8877_),
    .C(_8878_),
    .Y(_8879_)
);

AOI21X1 _19017_ (
    .A(_8861_),
    .B(_8862_),
    .C(_8477_),
    .Y(_8880_)
);

OAI21X1 _19018_ (
    .A(_8880_),
    .B(_8475_),
    .C(_8866_),
    .Y(_8881_)
);

OAI21X1 _19019_ (
    .A(_8515_),
    .B(_8485_),
    .C(_8523_),
    .Y(_8882_)
);

INVX2 _19020_ (
    .A(_8882_),
    .Y(_8883_)
);

AOI21X1 _19021_ (
    .A(_8849_),
    .B(_8850_),
    .C(_8482_),
    .Y(_8885_)
);

OAI21X1 _19022_ (
    .A(_8885_),
    .B(_8480_),
    .C(_8855_),
    .Y(_8886_)
);

NAND2X1 _19023_ (
    .A(_8587_),
    .B(_8593_),
    .Y(_8887_)
);

INVX2 _19024_ (
    .A(_8887_),
    .Y(_8888_)
);

AOI21X1 _19025_ (
    .A(_8836_),
    .B(_8837_),
    .C(_8601_),
    .Y(_8889_)
);

OAI21X1 _19026_ (
    .A(_8889_),
    .B(_8598_),
    .C(_8843_),
    .Y(_8890_)
);

NAND2X1 _19027_ (
    .A(_8572_),
    .B(_8581_),
    .Y(_8891_)
);

NOR2X1 _19028_ (
    .A(_2562__bF$buf4),
    .B(_7225__bF$buf0),
    .Y(_8892_)
);

INVX1 _19029_ (
    .A(_8892_),
    .Y(_8893_)
);

OAI21X1 _19030_ (
    .A(_8503_),
    .B(_8488_),
    .C(_8513_),
    .Y(_8894_)
);

NOR2X1 _19031_ (
    .A(_2825__bF$buf1),
    .B(_6815__bF$buf4),
    .Y(_8896_)
);

INVX2 _19032_ (
    .A(_8896_),
    .Y(_8897_)
);

OAI21X1 _19033_ (
    .A(_8501_),
    .B(_8491_),
    .C(_8495_),
    .Y(_8898_)
);

NAND2X1 _19034_ (
    .A(areg_6_bF$buf1),
    .B(breg_29_bF$buf3),
    .Y(_8899_)
);

INVX2 _19035_ (
    .A(_8899_),
    .Y(_8900_)
);

AND2X2 _19036_ (
    .A(areg_7_bF$buf2),
    .B(breg_28_bF$buf1),
    .Y(_8901_)
);

AND2X2 _19037_ (
    .A(areg_8_bF$buf3),
    .B(breg_27_bF$buf1),
    .Y(_8902_)
);

NAND2X1 _19038_ (
    .A(_8901_),
    .B(_8902_),
    .Y(_8903_)
);

OAI22X1 _19039_ (
    .A(_4434__bF$buf0),
    .B(_6050__bF$buf0),
    .C(_5190__bF$buf3),
    .D(_5668__bF$buf0),
    .Y(_8904_)
);

NAND3X1 _19040_ (
    .A(_8900_),
    .B(_8904_),
    .C(_8903_),
    .Y(_8905_)
);

NAND2X1 _19041_ (
    .A(areg_8_bF$buf2),
    .B(breg_28_bF$buf0),
    .Y(_8907_)
);

NOR2X1 _19042_ (
    .A(_8498_),
    .B(_8907_),
    .Y(_8908_)
);

NOR2X1 _19043_ (
    .A(_8901_),
    .B(_8902_),
    .Y(_8909_)
);

OAI21X1 _19044_ (
    .A(_8909_),
    .B(_8908_),
    .C(_8899_),
    .Y(_8910_)
);

AOI21X1 _19045_ (
    .A(_8905_),
    .B(_8910_),
    .C(_8898_),
    .Y(_8911_)
);

AOI21X1 _19046_ (
    .A(_8492_),
    .B(_8496_),
    .C(_8499_),
    .Y(_8912_)
);

OAI21X1 _19047_ (
    .A(_4434__bF$buf3),
    .B(_6050__bF$buf3),
    .C(_8902_),
    .Y(_8913_)
);

OAI21X1 _19048_ (
    .A(_5190__bF$buf2),
    .B(_5668__bF$buf5),
    .C(_8901_),
    .Y(_8914_)
);

AOI21X1 _19049_ (
    .A(_8913_),
    .B(_8914_),
    .C(_8899_),
    .Y(_8915_)
);

AOI21X1 _19050_ (
    .A(_8904_),
    .B(_8903_),
    .C(_8900_),
    .Y(_8916_)
);

NOR3X1 _19051_ (
    .A(_8916_),
    .B(_8912_),
    .C(_8915_),
    .Y(_8918_)
);

OAI21X1 _19052_ (
    .A(_8918_),
    .B(_8911_),
    .C(_8897_),
    .Y(_8919_)
);

OAI21X1 _19053_ (
    .A(_8915_),
    .B(_8916_),
    .C(_8912_),
    .Y(_8920_)
);

NAND3X1 _19054_ (
    .A(_8905_),
    .B(_8898_),
    .C(_8910_),
    .Y(_8921_)
);

NAND3X1 _19055_ (
    .A(_8896_),
    .B(_8920_),
    .C(_8921_),
    .Y(_8922_)
);

AOI21X1 _19056_ (
    .A(_8922_),
    .B(_8919_),
    .C(_8894_),
    .Y(_8923_)
);

AOI21X1 _19057_ (
    .A(_8487_),
    .B(_8512_),
    .C(_8509_),
    .Y(_8924_)
);

AOI21X1 _19058_ (
    .A(_8920_),
    .B(_8921_),
    .C(_8896_),
    .Y(_8925_)
);

NOR3X1 _19059_ (
    .A(_8911_),
    .B(_8897_),
    .C(_8918_),
    .Y(_8926_)
);

NOR3X1 _19060_ (
    .A(_8924_),
    .B(_8925_),
    .C(_8926_),
    .Y(_8927_)
);

OAI21X1 _19061_ (
    .A(_8927_),
    .B(_8923_),
    .C(_8893_),
    .Y(_8929_)
);

OAI21X1 _19062_ (
    .A(_8926_),
    .B(_8925_),
    .C(_8924_),
    .Y(_8930_)
);

NAND3X1 _19063_ (
    .A(_8894_),
    .B(_8922_),
    .C(_8919_),
    .Y(_8931_)
);

NAND3X1 _19064_ (
    .A(_8892_),
    .B(_8931_),
    .C(_8930_),
    .Y(_8932_)
);

AND2X2 _19065_ (
    .A(_8929_),
    .B(_8932_),
    .Y(_8933_)
);

OAI21X1 _19066_ (
    .A(_8568_),
    .B(_8570_),
    .C(_8560_),
    .Y(_8934_)
);

NAND2X1 _19067_ (
    .A(_8545_),
    .B(_8552_),
    .Y(_8935_)
);

OAI21X1 _19068_ (
    .A(_8535_),
    .B(_8530_),
    .C(_8538_),
    .Y(_8936_)
);

NAND2X1 _19069_ (
    .A(areg_9_bF$buf3),
    .B(breg_26_bF$buf0),
    .Y(_8937_)
);

NAND2X1 _19070_ (
    .A(areg_10_bF$buf2),
    .B(breg_25_bF$buf2),
    .Y(_8938_)
);

NAND2X1 _19071_ (
    .A(areg_11_bF$buf2),
    .B(breg_24_bF$buf3),
    .Y(_8940_)
);

NOR2X1 _19072_ (
    .A(_8938_),
    .B(_8940_),
    .Y(_8941_)
);

AND2X2 _19073_ (
    .A(_8938_),
    .B(_8940_),
    .Y(_8942_)
);

OAI21X1 _19074_ (
    .A(_8942_),
    .B(_8941_),
    .C(_8937_),
    .Y(_8943_)
);

INVX1 _19075_ (
    .A(_8937_),
    .Y(_8944_)
);

OR2X2 _19076_ (
    .A(_8938_),
    .B(_8940_),
    .Y(_8945_)
);

OAI21X1 _19077_ (
    .A(_9104__bF$buf2),
    .B(_5315__bF$buf3),
    .C(_8938_),
    .Y(_8946_)
);

NAND3X1 _19078_ (
    .A(_8944_),
    .B(_8946_),
    .C(_8945_),
    .Y(_8947_)
);

NAND2X1 _19079_ (
    .A(areg_13_bF$buf0),
    .B(breg_22_bF$buf1),
    .Y(_8948_)
);

AND2X2 _19080_ (
    .A(_8541_),
    .B(_8605_),
    .Y(_8949_)
);

OAI22X1 _19081_ (
    .A(_8192_),
    .B(_8948_),
    .C(_8949_),
    .D(_8603_),
    .Y(_8951_)
);

NAND3X1 _19082_ (
    .A(_8943_),
    .B(_8947_),
    .C(_8951_),
    .Y(_8952_)
);

AOI21X1 _19083_ (
    .A(_8946_),
    .B(_8945_),
    .C(_8944_),
    .Y(_8953_)
);

NOR3X1 _19084_ (
    .A(_8937_),
    .B(_8941_),
    .C(_8942_),
    .Y(_8954_)
);

NOR2X1 _19085_ (
    .A(_8541_),
    .B(_8605_),
    .Y(_8955_)
);

OAI21X1 _19086_ (
    .A(_549__bF$buf2),
    .B(_3781__bF$buf0),
    .C(_8541_),
    .Y(_8956_)
);

AOI21X1 _19087_ (
    .A(_8604_),
    .B(_8956_),
    .C(_8955_),
    .Y(_8957_)
);

OAI21X1 _19088_ (
    .A(_8954_),
    .B(_8953_),
    .C(_8957_),
    .Y(_8958_)
);

NAND3X1 _19089_ (
    .A(_8936_),
    .B(_8952_),
    .C(_8958_),
    .Y(_8959_)
);

INVX1 _19090_ (
    .A(_8936_),
    .Y(_8960_)
);

NAND3X1 _19091_ (
    .A(_8957_),
    .B(_8943_),
    .C(_8947_),
    .Y(_8962_)
);

OAI21X1 _19092_ (
    .A(_8954_),
    .B(_8953_),
    .C(_8951_),
    .Y(_8963_)
);

NAND3X1 _19093_ (
    .A(_8960_),
    .B(_8962_),
    .C(_8963_),
    .Y(_8964_)
);

AOI21X1 _19094_ (
    .A(_8623_),
    .B(_8627_),
    .C(_8608_),
    .Y(_8965_)
);

OAI21X1 _19095_ (
    .A(_8607_),
    .B(_8965_),
    .C(_8631_),
    .Y(_8966_)
);

NAND3X1 _19096_ (
    .A(_8959_),
    .B(_8964_),
    .C(_8966_),
    .Y(_8967_)
);

AOI21X1 _19097_ (
    .A(_8962_),
    .B(_8963_),
    .C(_8960_),
    .Y(_8968_)
);

AOI21X1 _19098_ (
    .A(_8952_),
    .B(_8958_),
    .C(_8936_),
    .Y(_8969_)
);

NOR3X1 _19099_ (
    .A(_8619_),
    .B(_8622_),
    .C(_8616_),
    .Y(_8970_)
);

AOI21X1 _19100_ (
    .A(_8633_),
    .B(_8630_),
    .C(_8970_),
    .Y(_8971_)
);

OAI21X1 _19101_ (
    .A(_8969_),
    .B(_8968_),
    .C(_8971_),
    .Y(_8973_)
);

NAND3X1 _19102_ (
    .A(_8935_),
    .B(_8973_),
    .C(_8967_),
    .Y(_8974_)
);

AND2X2 _19103_ (
    .A(_8552_),
    .B(_8545_),
    .Y(_8975_)
);

NAND3X1 _19104_ (
    .A(_8959_),
    .B(_8964_),
    .C(_8971_),
    .Y(_8976_)
);

OAI21X1 _19105_ (
    .A(_8969_),
    .B(_8968_),
    .C(_8966_),
    .Y(_8977_)
);

NAND3X1 _19106_ (
    .A(_8975_),
    .B(_8977_),
    .C(_8976_),
    .Y(_8978_)
);

NAND3X1 _19107_ (
    .A(_8974_),
    .B(_8978_),
    .C(_8934_),
    .Y(_8979_)
);

AOI21X1 _19108_ (
    .A(_8528_),
    .B(_8565_),
    .C(_8569_),
    .Y(_8980_)
);

AOI21X1 _19109_ (
    .A(_8977_),
    .B(_8976_),
    .C(_8975_),
    .Y(_8981_)
);

AOI21X1 _19110_ (
    .A(_8973_),
    .B(_8967_),
    .C(_8935_),
    .Y(_8982_)
);

OAI21X1 _19111_ (
    .A(_8981_),
    .B(_8982_),
    .C(_8980_),
    .Y(_8984_)
);

NAND3X1 _19112_ (
    .A(_8979_),
    .B(_8984_),
    .C(_8933_),
    .Y(_8985_)
);

NAND2X1 _19113_ (
    .A(_8932_),
    .B(_8929_),
    .Y(_8986_)
);

OAI21X1 _19114_ (
    .A(_8981_),
    .B(_8982_),
    .C(_8934_),
    .Y(_8987_)
);

NAND3X1 _19115_ (
    .A(_8974_),
    .B(_8978_),
    .C(_8980_),
    .Y(_8988_)
);

NAND3X1 _19116_ (
    .A(_8988_),
    .B(_8986_),
    .C(_8987_),
    .Y(_8989_)
);

OAI21X1 _19117_ (
    .A(_8689_),
    .B(_8688_),
    .C(_8685_),
    .Y(_8990_)
);

NAND3X1 _19118_ (
    .A(_8989_),
    .B(_8990_),
    .C(_8985_),
    .Y(_8991_)
);

AOI21X1 _19119_ (
    .A(_8988_),
    .B(_8987_),
    .C(_8986_),
    .Y(_8992_)
);

AOI21X1 _19120_ (
    .A(_8979_),
    .B(_8984_),
    .C(_8933_),
    .Y(_8993_)
);

AOI21X1 _19121_ (
    .A(_8602_),
    .B(_8681_),
    .C(_8690_),
    .Y(_8995_)
);

OAI21X1 _19122_ (
    .A(_8993_),
    .B(_8992_),
    .C(_8995_),
    .Y(_8996_)
);

NAND3X1 _19123_ (
    .A(_8891_),
    .B(_8991_),
    .C(_8996_),
    .Y(_8997_)
);

AND2X2 _19124_ (
    .A(_8581_),
    .B(_8572_),
    .Y(_8998_)
);

NAND3X1 _19125_ (
    .A(_8989_),
    .B(_8995_),
    .C(_8985_),
    .Y(_8999_)
);

OAI21X1 _19126_ (
    .A(_8993_),
    .B(_8992_),
    .C(_8990_),
    .Y(_9000_)
);

NAND3X1 _19127_ (
    .A(_8999_),
    .B(_9000_),
    .C(_8998_),
    .Y(_9001_)
);

NAND2X1 _19128_ (
    .A(_8997_),
    .B(_9001_),
    .Y(_9002_)
);

AOI21X1 _19129_ (
    .A(_8805_),
    .B(_8823_),
    .C(_8694_),
    .Y(_9003_)
);

OAI21X1 _19130_ (
    .A(_8692_),
    .B(_9003_),
    .C(_8829_),
    .Y(_9004_)
);

NAND2X1 _19131_ (
    .A(_8677_),
    .B(_8682_),
    .Y(_9006_)
);

NOR2X1 _19132_ (
    .A(_10869__bF$buf3),
    .B(_5369_),
    .Y(_9007_)
);

INVX2 _19133_ (
    .A(_9007_),
    .Y(_9008_)
);

NAND2X1 _19134_ (
    .A(areg_14_bF$buf0),
    .B(breg_21_bF$buf1),
    .Y(_9009_)
);

NOR2X1 _19135_ (
    .A(_8948_),
    .B(_9009_),
    .Y(_9010_)
);

AND2X2 _19136_ (
    .A(_8948_),
    .B(_9009_),
    .Y(_9011_)
);

NOR2X1 _19137_ (
    .A(_9010_),
    .B(_9011_),
    .Y(_9012_)
);

XNOR2X1 _19138_ (
    .A(_9012_),
    .B(_9008_),
    .Y(_9013_)
);

OAI21X1 _19139_ (
    .A(_8611_),
    .B(_8626_),
    .C(_8617_),
    .Y(_9014_)
);

NAND2X1 _19140_ (
    .A(areg_15_bF$buf3),
    .B(breg_20_bF$buf2),
    .Y(_9015_)
);

INVX2 _19141_ (
    .A(_9015_),
    .Y(_9017_)
);

AND2X2 _19142_ (
    .A(areg_16_bF$buf0),
    .B(breg_19_bF$buf1),
    .Y(_9018_)
);

AND2X2 _19143_ (
    .A(areg_17_bF$buf1),
    .B(breg_18_bF$buf1),
    .Y(_9019_)
);

NAND2X1 _19144_ (
    .A(_9018_),
    .B(_9019_),
    .Y(_9020_)
);

OAI21X1 _19145_ (
    .A(_2884__bF$buf1),
    .B(_3529__bF$buf1),
    .C(_8624_),
    .Y(_9021_)
);

NAND3X1 _19146_ (
    .A(_9017_),
    .B(_9021_),
    .C(_9020_),
    .Y(_9022_)
);

NAND2X1 _19147_ (
    .A(areg_17_bF$buf0),
    .B(breg_18_bF$buf0),
    .Y(_9023_)
);

NOR2X1 _19148_ (
    .A(_8624_),
    .B(_9023_),
    .Y(_9024_)
);

NOR2X1 _19149_ (
    .A(_9018_),
    .B(_9019_),
    .Y(_9025_)
);

OAI21X1 _19150_ (
    .A(_9025_),
    .B(_9024_),
    .C(_9015_),
    .Y(_9026_)
);

NAND3X1 _19151_ (
    .A(_9022_),
    .B(_9026_),
    .C(_9014_),
    .Y(_9028_)
);

AOI21X1 _19152_ (
    .A(_8609_),
    .B(_8618_),
    .C(_8625_),
    .Y(_9029_)
);

NOR3X1 _19153_ (
    .A(_9015_),
    .B(_9024_),
    .C(_9025_),
    .Y(_9030_)
);

AOI21X1 _19154_ (
    .A(_9021_),
    .B(_9020_),
    .C(_9017_),
    .Y(_9031_)
);

OAI21X1 _19155_ (
    .A(_9030_),
    .B(_9031_),
    .C(_9029_),
    .Y(_9032_)
);

NAND3X1 _19156_ (
    .A(_9028_),
    .B(_9032_),
    .C(_9013_),
    .Y(_9033_)
);

XNOR2X1 _19157_ (
    .A(_9012_),
    .B(_9007_),
    .Y(_9034_)
);

NOR3X1 _19158_ (
    .A(_9029_),
    .B(_9031_),
    .C(_9030_),
    .Y(_9035_)
);

AOI21X1 _19159_ (
    .A(_9022_),
    .B(_9026_),
    .C(_9014_),
    .Y(_9036_)
);

OAI21X1 _19160_ (
    .A(_9035_),
    .B(_9036_),
    .C(_9034_),
    .Y(_9037_)
);

NAND2X1 _19161_ (
    .A(_9033_),
    .B(_9037_),
    .Y(_9039_)
);

OAI21X1 _19162_ (
    .A(_8671_),
    .B(_8638_),
    .C(_8663_),
    .Y(_9040_)
);

AND2X2 _19163_ (
    .A(breg_16_bF$buf1),
    .B(areg_19_bF$buf3),
    .Y(_9041_)
);

AOI21X1 _19164_ (
    .A(_8229_),
    .B(_9041_),
    .C(_8655_),
    .Y(_9042_)
);

NAND2X1 _19165_ (
    .A(breg_17_bF$buf0),
    .B(areg_18_bF$buf1),
    .Y(_9043_)
);

INVX1 _19166_ (
    .A(_9043_),
    .Y(_9044_)
);

AND2X2 _19167_ (
    .A(breg_15_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_9045_)
);

NAND2X1 _19168_ (
    .A(_9041_),
    .B(_9045_),
    .Y(_9046_)
);

OAI22X1 _19169_ (
    .A(_2362__bF$buf4),
    .B(_3958__bF$buf2),
    .C(_2560__bF$buf1),
    .D(_3402__bF$buf3),
    .Y(_9047_)
);

NAND3X1 _19170_ (
    .A(_9044_),
    .B(_9047_),
    .C(_9046_),
    .Y(_9048_)
);

OAI21X1 _19171_ (
    .A(_2560__bF$buf0),
    .B(_3402__bF$buf2),
    .C(_9045_),
    .Y(_9050_)
);

OAI21X1 _19172_ (
    .A(_2362__bF$buf3),
    .B(_3958__bF$buf1),
    .C(_9041_),
    .Y(_9051_)
);

NAND3X1 _19173_ (
    .A(_9043_),
    .B(_9050_),
    .C(_9051_),
    .Y(_9052_)
);

NOR2X1 _19174_ (
    .A(_8657_),
    .B(_8699_),
    .Y(_9053_)
);

OAI21X1 _19175_ (
    .A(_2586__bF$buf1),
    .B(_4551__bF$buf1),
    .C(_8657_),
    .Y(_9054_)
);

AOI21X1 _19176_ (
    .A(_8697_),
    .B(_9054_),
    .C(_9053_),
    .Y(_9055_)
);

NAND3X1 _19177_ (
    .A(_9055_),
    .B(_9048_),
    .C(_9052_),
    .Y(_9056_)
);

AOI21X1 _19178_ (
    .A(_9050_),
    .B(_9051_),
    .C(_9043_),
    .Y(_9057_)
);

AOI21X1 _19179_ (
    .A(_9047_),
    .B(_9046_),
    .C(_9044_),
    .Y(_9058_)
);

NAND2X1 _19180_ (
    .A(breg_13_bF$buf2),
    .B(areg_22_bF$buf2),
    .Y(_9059_)
);

AND2X2 _19181_ (
    .A(_8657_),
    .B(_8699_),
    .Y(_9061_)
);

OAI22X1 _19182_ (
    .A(_8286_),
    .B(_9059_),
    .C(_9061_),
    .D(_8696_),
    .Y(_9062_)
);

OAI21X1 _19183_ (
    .A(_9057_),
    .B(_9058_),
    .C(_9062_),
    .Y(_9063_)
);

AOI21X1 _19184_ (
    .A(_9056_),
    .B(_9063_),
    .C(_9042_),
    .Y(_9064_)
);

INVX1 _19185_ (
    .A(_8641_),
    .Y(_9065_)
);

OAI21X1 _19186_ (
    .A(_8644_),
    .B(_9065_),
    .C(_8646_),
    .Y(_9066_)
);

NAND3X1 _19187_ (
    .A(_9048_),
    .B(_9052_),
    .C(_9062_),
    .Y(_9067_)
);

OAI21X1 _19188_ (
    .A(_9057_),
    .B(_9058_),
    .C(_9055_),
    .Y(_9068_)
);

AOI21X1 _19189_ (
    .A(_9067_),
    .B(_9068_),
    .C(_9066_),
    .Y(_9069_)
);

OAI21X1 _19190_ (
    .A(_9064_),
    .B(_9069_),
    .C(_9040_),
    .Y(_9070_)
);

AOI21X1 _19191_ (
    .A(_8662_),
    .B(_8664_),
    .C(_8670_),
    .Y(_9072_)
);

NAND3X1 _19192_ (
    .A(_9066_),
    .B(_9067_),
    .C(_9068_),
    .Y(_9073_)
);

NOR3X1 _19193_ (
    .A(_9058_),
    .B(_9055_),
    .C(_9057_),
    .Y(_9074_)
);

AOI21X1 _19194_ (
    .A(_9048_),
    .B(_9052_),
    .C(_9062_),
    .Y(_9075_)
);

OAI21X1 _19195_ (
    .A(_9074_),
    .B(_9075_),
    .C(_9042_),
    .Y(_9076_)
);

NAND3X1 _19196_ (
    .A(_9072_),
    .B(_9073_),
    .C(_9076_),
    .Y(_9077_)
);

AOI21X1 _19197_ (
    .A(_9070_),
    .B(_9077_),
    .C(_9039_),
    .Y(_9078_)
);

AND2X2 _19198_ (
    .A(_9037_),
    .B(_9033_),
    .Y(_9079_)
);

NAND3X1 _19199_ (
    .A(_9040_),
    .B(_9073_),
    .C(_9076_),
    .Y(_9080_)
);

OAI21X1 _19200_ (
    .A(_9064_),
    .B(_9069_),
    .C(_9072_),
    .Y(_9081_)
);

AOI21X1 _19201_ (
    .A(_9080_),
    .B(_9081_),
    .C(_9079_),
    .Y(_9082_)
);

AOI21X1 _19202_ (
    .A(_8695_),
    .B(_8729_),
    .C(_8738_),
    .Y(_9083_)
);

OAI21X1 _19203_ (
    .A(_9082_),
    .B(_9078_),
    .C(_9083_),
    .Y(_9084_)
);

NAND3X1 _19204_ (
    .A(_9080_),
    .B(_9081_),
    .C(_9079_),
    .Y(_9085_)
);

NAND3X1 _19205_ (
    .A(_9070_),
    .B(_9039_),
    .C(_9077_),
    .Y(_9086_)
);

OAI21X1 _19206_ (
    .A(_8737_),
    .B(_8736_),
    .C(_8734_),
    .Y(_9087_)
);

NAND3X1 _19207_ (
    .A(_9086_),
    .B(_9087_),
    .C(_9085_),
    .Y(_9088_)
);

NAND3X1 _19208_ (
    .A(_9006_),
    .B(_9088_),
    .C(_9084_),
    .Y(_9089_)
);

INVX2 _19209_ (
    .A(_9006_),
    .Y(_9090_)
);

AOI21X1 _19210_ (
    .A(_9086_),
    .B(_9085_),
    .C(_9087_),
    .Y(_9091_)
);

NOR3X1 _19211_ (
    .A(_9082_),
    .B(_9078_),
    .C(_9083_),
    .Y(_9093_)
);

OAI21X1 _19212_ (
    .A(_9093_),
    .B(_9091_),
    .C(_9090_),
    .Y(_9094_)
);

NAND2X1 _19213_ (
    .A(_9089_),
    .B(_9094_),
    .Y(_9095_)
);

OAI21X1 _19214_ (
    .A(_8740_),
    .B(_8822_),
    .C(_8799_),
    .Y(_9096_)
);

NAND2X1 _19215_ (
    .A(_8725_),
    .B(_8730_),
    .Y(_9097_)
);

NAND2X1 _19216_ (
    .A(breg_14_bF$buf0),
    .B(areg_21_bF$buf2),
    .Y(_9098_)
);

INVX2 _19217_ (
    .A(_9098_),
    .Y(_9099_)
);

NAND2X1 _19218_ (
    .A(breg_12_bF$buf0),
    .B(areg_23_bF$buf4),
    .Y(_9100_)
);

XOR2X1 _19219_ (
    .A(_9059_),
    .B(_9100_),
    .Y(_9101_)
);

XNOR2X1 _19220_ (
    .A(_9101_),
    .B(_9099_),
    .Y(_9102_)
);

OAI21X1 _19221_ (
    .A(_8719_),
    .B(_8703_),
    .C(_8711_),
    .Y(_9105_)
);

NAND2X1 _19222_ (
    .A(breg_11_bF$buf2),
    .B(areg_24_bF$buf3),
    .Y(_9106_)
);

NAND2X1 _19223_ (
    .A(breg_10_bF$buf1),
    .B(areg_26_bF$buf1),
    .Y(_9107_)
);

NOR2X1 _19224_ (
    .A(_8717_),
    .B(_9107_),
    .Y(_9108_)
);

AND2X2 _19225_ (
    .A(breg_10_bF$buf0),
    .B(areg_25_bF$buf0),
    .Y(_9109_)
);

AND2X2 _19226_ (
    .A(breg_9_bF$buf4),
    .B(areg_26_bF$buf0),
    .Y(_9110_)
);

NOR2X1 _19227_ (
    .A(_9109_),
    .B(_9110_),
    .Y(_9111_)
);

NOR3X1 _19228_ (
    .A(_9106_),
    .B(_9108_),
    .C(_9111_),
    .Y(_9112_)
);

INVX2 _19229_ (
    .A(_9106_),
    .Y(_9113_)
);

NAND2X1 _19230_ (
    .A(_9109_),
    .B(_9110_),
    .Y(_9114_)
);

OAI22X1 _19231_ (
    .A(_6044__bF$buf0),
    .B(_6686__bF$buf3),
    .C(_7217__bF$buf4),
    .D(_6300__bF$buf0),
    .Y(_9116_)
);

AOI21X1 _19232_ (
    .A(_9116_),
    .B(_9114_),
    .C(_9113_),
    .Y(_9117_)
);

OAI21X1 _19233_ (
    .A(_9112_),
    .B(_9117_),
    .C(_9105_),
    .Y(_9118_)
);

AOI21X1 _19234_ (
    .A(_8710_),
    .B(_8712_),
    .C(_8718_),
    .Y(_9119_)
);

NAND3X1 _19235_ (
    .A(_9113_),
    .B(_9116_),
    .C(_9114_),
    .Y(_9120_)
);

OAI21X1 _19236_ (
    .A(_9111_),
    .B(_9108_),
    .C(_9106_),
    .Y(_9121_)
);

NAND3X1 _19237_ (
    .A(_9119_),
    .B(_9120_),
    .C(_9121_),
    .Y(_9122_)
);

AOI21X1 _19238_ (
    .A(_9122_),
    .B(_9118_),
    .C(_9102_),
    .Y(_9123_)
);

XNOR2X1 _19239_ (
    .A(_9101_),
    .B(_9098_),
    .Y(_9124_)
);

NAND3X1 _19240_ (
    .A(_9120_),
    .B(_9105_),
    .C(_9121_),
    .Y(_9125_)
);

OAI21X1 _19241_ (
    .A(_9112_),
    .B(_9117_),
    .C(_9119_),
    .Y(_9127_)
);

AOI21X1 _19242_ (
    .A(_9125_),
    .B(_9127_),
    .C(_9124_),
    .Y(_9128_)
);

AOI21X1 _19243_ (
    .A(_8766_),
    .B(_8762_),
    .C(_8767_),
    .Y(_9129_)
);

OAI21X1 _19244_ (
    .A(_9123_),
    .B(_9128_),
    .C(_9129_),
    .Y(_9130_)
);

NAND3X1 _19245_ (
    .A(_9125_),
    .B(_9127_),
    .C(_9124_),
    .Y(_9131_)
);

NAND3X1 _19246_ (
    .A(_9122_),
    .B(_9118_),
    .C(_9102_),
    .Y(_9132_)
);

OAI21X1 _19247_ (
    .A(_8768_),
    .B(_8744_),
    .C(_8756_),
    .Y(_9133_)
);

NAND3X1 _19248_ (
    .A(_9133_),
    .B(_9131_),
    .C(_9132_),
    .Y(_9134_)
);

NAND3X1 _19249_ (
    .A(_9097_),
    .B(_9134_),
    .C(_9130_),
    .Y(_9135_)
);

AND2X2 _19250_ (
    .A(_8730_),
    .B(_8725_),
    .Y(_9136_)
);

AOI21X1 _19251_ (
    .A(_9131_),
    .B(_9132_),
    .C(_9133_),
    .Y(_9138_)
);

NOR3X1 _19252_ (
    .A(_9128_),
    .B(_9129_),
    .C(_9123_),
    .Y(_9139_)
);

OAI21X1 _19253_ (
    .A(_9139_),
    .B(_9138_),
    .C(_9136_),
    .Y(_9140_)
);

NAND2X1 _19254_ (
    .A(_9135_),
    .B(_9140_),
    .Y(_9141_)
);

AND2X2 _19255_ (
    .A(breg_7_bF$buf3),
    .B(areg_28_bF$buf4),
    .Y(_9142_)
);

AOI21X1 _19256_ (
    .A(_8339_),
    .B(_9142_),
    .C(_8757_),
    .Y(_9143_)
);

NAND2X1 _19257_ (
    .A(breg[8]),
    .B(areg_27_bF$buf4),
    .Y(_9144_)
);

INVX1 _19258_ (
    .A(_9144_),
    .Y(_9145_)
);

AND2X2 _19259_ (
    .A(breg_6_bF$buf4),
    .B(areg_29_bF$buf4),
    .Y(_9146_)
);

NAND2X1 _19260_ (
    .A(_9142_),
    .B(_9146_),
    .Y(_9147_)
);

NAND2X1 _19261_ (
    .A(breg_6_bF$buf3),
    .B(areg_29_bF$buf3),
    .Y(_9149_)
);

OAI21X1 _19262_ (
    .A(_4116__bF$buf2),
    .B(_7520__bF$buf0),
    .C(_9149_),
    .Y(_9150_)
);

NAND3X1 _19263_ (
    .A(_9145_),
    .B(_9150_),
    .C(_9147_),
    .Y(_9151_)
);

OAI21X1 _19264_ (
    .A(_4116__bF$buf1),
    .B(_7520__bF$buf3),
    .C(_9146_),
    .Y(_9152_)
);

INVX4 _19265_ (
    .A(areg_29_bF$buf2),
    .Y(_9153_)
);

OAI21X1 _19266_ (
    .A(_5453__bF$buf5),
    .B(_9153_),
    .C(_9142_),
    .Y(_9154_)
);

NAND3X1 _19267_ (
    .A(_9144_),
    .B(_9152_),
    .C(_9154_),
    .Y(_9155_)
);

NAND2X1 _19268_ (
    .A(breg_3_bF$buf3),
    .B(areg_31_bF$buf1),
    .Y(_9156_)
);

NOR2X1 _19269_ (
    .A(_8369_),
    .B(_9156_),
    .Y(_9157_)
);

AOI21X1 _19270_ (
    .A(_8780_),
    .B(_8774_),
    .C(_9157_),
    .Y(_9158_)
);

NAND3X1 _19271_ (
    .A(_9158_),
    .B(_9151_),
    .C(_9155_),
    .Y(_9160_)
);

AOI21X1 _19272_ (
    .A(_9152_),
    .B(_9154_),
    .C(_9144_),
    .Y(_9161_)
);

AOI21X1 _19273_ (
    .A(_9150_),
    .B(_9147_),
    .C(_9145_),
    .Y(_9162_)
);

AND2X2 _19274_ (
    .A(_8369_),
    .B(_9156_),
    .Y(_9163_)
);

OAI22X1 _19275_ (
    .A(_8364_),
    .B(_8772_),
    .C(_9163_),
    .D(_8771_),
    .Y(_9164_)
);

OAI21X1 _19276_ (
    .A(_9161_),
    .B(_9162_),
    .C(_9164_),
    .Y(_9165_)
);

AOI21X1 _19277_ (
    .A(_9160_),
    .B(_9165_),
    .C(_9143_),
    .Y(_9166_)
);

INVX1 _19278_ (
    .A(_9142_),
    .Y(_9167_)
);

OAI21X1 _19279_ (
    .A(_8765_),
    .B(_9167_),
    .C(_8750_),
    .Y(_9168_)
);

NAND3X1 _19280_ (
    .A(_9151_),
    .B(_9155_),
    .C(_9164_),
    .Y(_9169_)
);

OAI21X1 _19281_ (
    .A(_9161_),
    .B(_9162_),
    .C(_9158_),
    .Y(_9171_)
);

AOI21X1 _19282_ (
    .A(_9169_),
    .B(_9171_),
    .C(_9168_),
    .Y(_9172_)
);

NAND2X1 _19283_ (
    .A(breg_5_bF$buf2),
    .B(areg_31_bF$buf0),
    .Y(_9173_)
);

OAI21X1 _19284_ (
    .A(_4258__bF$buf3),
    .B(_8759_),
    .C(_8772_),
    .Y(_9174_)
);

OAI21X1 _19285_ (
    .A(_8369_),
    .B(_9173_),
    .C(_9174_),
    .Y(_9175_)
);

OAI21X1 _19286_ (
    .A(_9172_),
    .B(_9166_),
    .C(_9175_),
    .Y(_9176_)
);

NAND3X1 _19287_ (
    .A(_9168_),
    .B(_9169_),
    .C(_9171_),
    .Y(_9177_)
);

NOR3X1 _19288_ (
    .A(_9162_),
    .B(_9158_),
    .C(_9161_),
    .Y(_9178_)
);

AOI21X1 _19289_ (
    .A(_9151_),
    .B(_9155_),
    .C(_9164_),
    .Y(_9179_)
);

OAI21X1 _19290_ (
    .A(_9178_),
    .B(_9179_),
    .C(_9143_),
    .Y(_9180_)
);

INVX1 _19291_ (
    .A(_9175_),
    .Y(_9182_)
);

NAND3X1 _19292_ (
    .A(_9177_),
    .B(_9182_),
    .C(_9180_),
    .Y(_9183_)
);

NAND2X1 _19293_ (
    .A(_9176_),
    .B(_9183_),
    .Y(_9184_)
);

OAI21X1 _19294_ (
    .A(_8816_),
    .B(_8783_),
    .C(_9184_),
    .Y(_9185_)
);

NOR2X1 _19295_ (
    .A(_8816_),
    .B(_8783_),
    .Y(_9186_)
);

NAND3X1 _19296_ (
    .A(_9176_),
    .B(_9183_),
    .C(_9186_),
    .Y(_9187_)
);

AOI21X1 _19297_ (
    .A(_9185_),
    .B(_9187_),
    .C(_9141_),
    .Y(_9188_)
);

OAI21X1 _19298_ (
    .A(_9139_),
    .B(_9138_),
    .C(_9097_),
    .Y(_9189_)
);

NAND3X1 _19299_ (
    .A(_9134_),
    .B(_9136_),
    .C(_9130_),
    .Y(_9190_)
);

NAND2X1 _19300_ (
    .A(_9190_),
    .B(_9189_),
    .Y(_9191_)
);

NAND2X1 _19301_ (
    .A(_8787_),
    .B(_8813_),
    .Y(_9193_)
);

NAND3X1 _19302_ (
    .A(_9176_),
    .B(_9183_),
    .C(_9193_),
    .Y(_9194_)
);

NAND2X1 _19303_ (
    .A(_9184_),
    .B(_9186_),
    .Y(_9195_)
);

AOI21X1 _19304_ (
    .A(_9194_),
    .B(_9195_),
    .C(_9191_),
    .Y(_9196_)
);

OAI21X1 _19305_ (
    .A(_9188_),
    .B(_9196_),
    .C(_9096_),
    .Y(_9197_)
);

AOI21X1 _19306_ (
    .A(_8800_),
    .B(_8798_),
    .C(_8821_),
    .Y(_9198_)
);

NAND3X1 _19307_ (
    .A(_9194_),
    .B(_9195_),
    .C(_9191_),
    .Y(_9199_)
);

NOR2X1 _19308_ (
    .A(_9184_),
    .B(_9186_),
    .Y(_9200_)
);

AOI21X1 _19309_ (
    .A(_9176_),
    .B(_9183_),
    .C(_9193_),
    .Y(_9201_)
);

OAI21X1 _19310_ (
    .A(_9200_),
    .B(_9201_),
    .C(_9141_),
    .Y(_9202_)
);

NAND3X1 _19311_ (
    .A(_9202_),
    .B(_9198_),
    .C(_9199_),
    .Y(_9204_)
);

AOI21X1 _19312_ (
    .A(_9204_),
    .B(_9197_),
    .C(_9095_),
    .Y(_9205_)
);

OAI21X1 _19313_ (
    .A(_9093_),
    .B(_9091_),
    .C(_9006_),
    .Y(_9206_)
);

NAND3X1 _19314_ (
    .A(_9084_),
    .B(_9088_),
    .C(_9090_),
    .Y(_9207_)
);

NAND2X1 _19315_ (
    .A(_9207_),
    .B(_9206_),
    .Y(_9208_)
);

NAND3X1 _19316_ (
    .A(_9202_),
    .B(_9096_),
    .C(_9199_),
    .Y(_9209_)
);

OAI21X1 _19317_ (
    .A(_9188_),
    .B(_9196_),
    .C(_9198_),
    .Y(_9210_)
);

AOI21X1 _19318_ (
    .A(_9209_),
    .B(_9210_),
    .C(_9208_),
    .Y(_9211_)
);

OAI21X1 _19319_ (
    .A(_9205_),
    .B(_9211_),
    .C(_9004_),
    .Y(_9212_)
);

NOR3X1 _19320_ (
    .A(_8794_),
    .B(_8801_),
    .C(_8804_),
    .Y(_9213_)
);

AOI21X1 _19321_ (
    .A(_8831_),
    .B(_8828_),
    .C(_9213_),
    .Y(_9215_)
);

NAND3X1 _19322_ (
    .A(_9209_),
    .B(_9210_),
    .C(_9208_),
    .Y(_9216_)
);

NAND3X1 _19323_ (
    .A(_9204_),
    .B(_9197_),
    .C(_9095_),
    .Y(_9217_)
);

NAND3X1 _19324_ (
    .A(_9216_),
    .B(_9217_),
    .C(_9215_),
    .Y(_9218_)
);

AOI21X1 _19325_ (
    .A(_9218_),
    .B(_9212_),
    .C(_9002_),
    .Y(_9219_)
);

AOI21X1 _19326_ (
    .A(_8999_),
    .B(_9000_),
    .C(_8998_),
    .Y(_9220_)
);

AOI21X1 _19327_ (
    .A(_8991_),
    .B(_8996_),
    .C(_8891_),
    .Y(_9221_)
);

NOR2X1 _19328_ (
    .A(_9220_),
    .B(_9221_),
    .Y(_9222_)
);

NAND3X1 _19329_ (
    .A(_9216_),
    .B(_9004_),
    .C(_9217_),
    .Y(_9223_)
);

OAI21X1 _19330_ (
    .A(_9205_),
    .B(_9211_),
    .C(_9215_),
    .Y(_9224_)
);

AOI21X1 _19331_ (
    .A(_9223_),
    .B(_9224_),
    .C(_9222_),
    .Y(_9226_)
);

OAI21X1 _19332_ (
    .A(_9219_),
    .B(_9226_),
    .C(_8890_),
    .Y(_9227_)
);

NOR3X1 _19333_ (
    .A(_8825_),
    .B(_8832_),
    .C(_8835_),
    .Y(_9228_)
);

AOI21X1 _19334_ (
    .A(_8842_),
    .B(_8844_),
    .C(_9228_),
    .Y(_9229_)
);

NAND3X1 _19335_ (
    .A(_9223_),
    .B(_9224_),
    .C(_9222_),
    .Y(_9230_)
);

NAND3X1 _19336_ (
    .A(_9002_),
    .B(_9218_),
    .C(_9212_),
    .Y(_9231_)
);

NAND3X1 _19337_ (
    .A(_9231_),
    .B(_9230_),
    .C(_9229_),
    .Y(_9232_)
);

AOI21X1 _19338_ (
    .A(_9232_),
    .B(_9227_),
    .C(_8888_),
    .Y(_9233_)
);

NAND3X1 _19339_ (
    .A(_9231_),
    .B(_8890_),
    .C(_9230_),
    .Y(_9234_)
);

OAI21X1 _19340_ (
    .A(_9219_),
    .B(_9226_),
    .C(_9229_),
    .Y(_9235_)
);

AOI21X1 _19341_ (
    .A(_9234_),
    .B(_9235_),
    .C(_8887_),
    .Y(_9237_)
);

OAI21X1 _19342_ (
    .A(_9233_),
    .B(_9237_),
    .C(_8886_),
    .Y(_9238_)
);

NOR3X1 _19343_ (
    .A(_8839_),
    .B(_8845_),
    .C(_8848_),
    .Y(_9239_)
);

AOI21X1 _19344_ (
    .A(_8479_),
    .B(_8856_),
    .C(_9239_),
    .Y(_9240_)
);

NAND3X1 _19345_ (
    .A(_8887_),
    .B(_9234_),
    .C(_9235_),
    .Y(_9241_)
);

NAND3X1 _19346_ (
    .A(_8888_),
    .B(_9232_),
    .C(_9227_),
    .Y(_9242_)
);

NAND3X1 _19347_ (
    .A(_9241_),
    .B(_9242_),
    .C(_9240_),
    .Y(_9243_)
);

AOI21X1 _19348_ (
    .A(_9243_),
    .B(_9238_),
    .C(_8883_),
    .Y(_9244_)
);

NAND3X1 _19349_ (
    .A(_8886_),
    .B(_9241_),
    .C(_9242_),
    .Y(_9245_)
);

OAI21X1 _19350_ (
    .A(_9233_),
    .B(_9237_),
    .C(_9240_),
    .Y(_9246_)
);

AOI21X1 _19351_ (
    .A(_9245_),
    .B(_9246_),
    .C(_8882_),
    .Y(_9248_)
);

OAI21X1 _19352_ (
    .A(_9244_),
    .B(_9248_),
    .C(_8881_),
    .Y(_9249_)
);

NOR3X1 _19353_ (
    .A(_8854_),
    .B(_8857_),
    .C(_8860_),
    .Y(_9250_)
);

AOI21X1 _19354_ (
    .A(_8474_),
    .B(_8867_),
    .C(_9250_),
    .Y(_9251_)
);

NAND3X1 _19355_ (
    .A(_8882_),
    .B(_9245_),
    .C(_9246_),
    .Y(_9252_)
);

NAND3X1 _19356_ (
    .A(_8883_),
    .B(_9243_),
    .C(_9238_),
    .Y(_9253_)
);

NAND3X1 _19357_ (
    .A(_9252_),
    .B(_9253_),
    .C(_9251_),
    .Y(_9254_)
);

NAND2X1 _19358_ (
    .A(_9254_),
    .B(_9249_),
    .Y(_9255_)
);

XNOR2X1 _19359_ (
    .A(_8879_),
    .B(_9255_),
    .Y(_0_[35])
);

AOI22X1 _19360_ (
    .A(_8869_),
    .B(_8875_),
    .C(_9249_),
    .D(_9254_),
    .Y(_9256_)
);

NAND2X1 _19361_ (
    .A(_9252_),
    .B(_9253_),
    .Y(_9258_)
);

OR2X2 _19362_ (
    .A(_9258_),
    .B(_9251_),
    .Y(_9259_)
);

OAI21X1 _19363_ (
    .A(_9244_),
    .B(_9248_),
    .C(_9251_),
    .Y(_9260_)
);

NAND2X1 _19364_ (
    .A(_9260_),
    .B(_8878_),
    .Y(_9261_)
);

NAND2X1 _19365_ (
    .A(_9259_),
    .B(_9261_),
    .Y(_9262_)
);

AOI21X1 _19366_ (
    .A(_9256_),
    .B(_8469_),
    .C(_9262_),
    .Y(_9263_)
);

NAND2X1 _19367_ (
    .A(_9256_),
    .B(_8470_),
    .Y(_9264_)
);

OAI21X1 _19368_ (
    .A(_7651_),
    .B(_9264_),
    .C(_9263_),
    .Y(_9265_)
);

AOI21X1 _19369_ (
    .A(_9241_),
    .B(_9242_),
    .C(_8886_),
    .Y(_9266_)
);

OAI21X1 _19370_ (
    .A(_9266_),
    .B(_8883_),
    .C(_9245_),
    .Y(_9267_)
);

OAI21X1 _19371_ (
    .A(_8923_),
    .B(_8893_),
    .C(_8931_),
    .Y(_9269_)
);

INVX2 _19372_ (
    .A(_9269_),
    .Y(_9270_)
);

AOI21X1 _19373_ (
    .A(_9231_),
    .B(_9230_),
    .C(_8890_),
    .Y(_9271_)
);

OAI21X1 _19374_ (
    .A(_9271_),
    .B(_8888_),
    .C(_9234_),
    .Y(_9272_)
);

NAND2X1 _19375_ (
    .A(_8991_),
    .B(_8997_),
    .Y(_9273_)
);

INVX2 _19376_ (
    .A(_9273_),
    .Y(_9274_)
);

AOI21X1 _19377_ (
    .A(_9216_),
    .B(_9217_),
    .C(_9004_),
    .Y(_9275_)
);

OAI21X1 _19378_ (
    .A(_9275_),
    .B(_9002_),
    .C(_9223_),
    .Y(_9276_)
);

NAND2X1 _19379_ (
    .A(_8979_),
    .B(_8985_),
    .Y(_9277_)
);

NOR2X1 _19380_ (
    .A(_2825__bF$buf0),
    .B(_7225__bF$buf4),
    .Y(_9278_)
);

INVX1 _19381_ (
    .A(_9278_),
    .Y(_9280_)
);

OAI21X1 _19382_ (
    .A(_8911_),
    .B(_8897_),
    .C(_8921_),
    .Y(_9281_)
);

NOR2X1 _19383_ (
    .A(_3646__bF$buf1),
    .B(_6815__bF$buf3),
    .Y(_9282_)
);

INVX2 _19384_ (
    .A(_9282_),
    .Y(_9283_)
);

OAI21X1 _19385_ (
    .A(_8909_),
    .B(_8899_),
    .C(_8903_),
    .Y(_9284_)
);

NAND2X1 _19386_ (
    .A(areg_7_bF$buf1),
    .B(breg_29_bF$buf2),
    .Y(_9285_)
);

INVX2 _19387_ (
    .A(_9285_),
    .Y(_9286_)
);

AND2X2 _19388_ (
    .A(areg_8_bF$buf1),
    .B(breg_28_bF$buf5),
    .Y(_9287_)
);

AND2X2 _19389_ (
    .A(areg_9_bF$buf2),
    .B(breg_27_bF$buf0),
    .Y(_9288_)
);

NAND2X1 _19390_ (
    .A(_9287_),
    .B(_9288_),
    .Y(_9289_)
);

OAI21X1 _19391_ (
    .A(_6582__bF$buf3),
    .B(_5668__bF$buf4),
    .C(_8907_),
    .Y(_9291_)
);

NAND3X1 _19392_ (
    .A(_9286_),
    .B(_9291_),
    .C(_9289_),
    .Y(_9292_)
);

NAND2X1 _19393_ (
    .A(areg_9_bF$buf1),
    .B(breg_27_bF$buf5),
    .Y(_9293_)
);

NOR2X1 _19394_ (
    .A(_8907_),
    .B(_9293_),
    .Y(_9294_)
);

NOR2X1 _19395_ (
    .A(_9287_),
    .B(_9288_),
    .Y(_9295_)
);

OAI21X1 _19396_ (
    .A(_9295_),
    .B(_9294_),
    .C(_9285_),
    .Y(_9296_)
);

AOI21X1 _19397_ (
    .A(_9292_),
    .B(_9296_),
    .C(_9284_),
    .Y(_9297_)
);

AOI21X1 _19398_ (
    .A(_8900_),
    .B(_8904_),
    .C(_8908_),
    .Y(_9298_)
);

NOR3X1 _19399_ (
    .A(_9285_),
    .B(_9294_),
    .C(_9295_),
    .Y(_9299_)
);

AOI21X1 _19400_ (
    .A(_9291_),
    .B(_9289_),
    .C(_9286_),
    .Y(_9300_)
);

NOR3X1 _19401_ (
    .A(_9300_),
    .B(_9298_),
    .C(_9299_),
    .Y(_9302_)
);

OAI21X1 _19402_ (
    .A(_9302_),
    .B(_9297_),
    .C(_9283_),
    .Y(_9303_)
);

OAI21X1 _19403_ (
    .A(_9299_),
    .B(_9300_),
    .C(_9298_),
    .Y(_9304_)
);

NAND3X1 _19404_ (
    .A(_9292_),
    .B(_9284_),
    .C(_9296_),
    .Y(_9305_)
);

NAND3X1 _19405_ (
    .A(_9282_),
    .B(_9305_),
    .C(_9304_),
    .Y(_9306_)
);

AOI21X1 _19406_ (
    .A(_9306_),
    .B(_9303_),
    .C(_9281_),
    .Y(_9307_)
);

AOI21X1 _19407_ (
    .A(_8896_),
    .B(_8920_),
    .C(_8918_),
    .Y(_9308_)
);

AOI21X1 _19408_ (
    .A(_9305_),
    .B(_9304_),
    .C(_9282_),
    .Y(_9309_)
);

NOR3X1 _19409_ (
    .A(_9297_),
    .B(_9283_),
    .C(_9302_),
    .Y(_9310_)
);

NOR3X1 _19410_ (
    .A(_9308_),
    .B(_9309_),
    .C(_9310_),
    .Y(_9311_)
);

OAI21X1 _19411_ (
    .A(_9311_),
    .B(_9307_),
    .C(_9280_),
    .Y(_9313_)
);

OAI21X1 _19412_ (
    .A(_9310_),
    .B(_9309_),
    .C(_9308_),
    .Y(_9314_)
);

NAND3X1 _19413_ (
    .A(_9281_),
    .B(_9306_),
    .C(_9303_),
    .Y(_9315_)
);

NAND3X1 _19414_ (
    .A(_9278_),
    .B(_9315_),
    .C(_9314_),
    .Y(_9316_)
);

AND2X2 _19415_ (
    .A(_9313_),
    .B(_9316_),
    .Y(_9317_)
);

AOI21X1 _19416_ (
    .A(_8959_),
    .B(_8964_),
    .C(_8966_),
    .Y(_9318_)
);

OAI21X1 _19417_ (
    .A(_9318_),
    .B(_8975_),
    .C(_8967_),
    .Y(_9319_)
);

NAND2X1 _19418_ (
    .A(_8952_),
    .B(_8959_),
    .Y(_9320_)
);

OAI21X1 _19419_ (
    .A(_8942_),
    .B(_8937_),
    .C(_8945_),
    .Y(_9321_)
);

NAND2X1 _19420_ (
    .A(areg_10_bF$buf1),
    .B(breg_26_bF$buf4),
    .Y(_9322_)
);

NAND2X1 _19421_ (
    .A(areg_11_bF$buf1),
    .B(breg_25_bF$buf1),
    .Y(_9324_)
);

NAND2X1 _19422_ (
    .A(areg_12_bF$buf2),
    .B(breg_24_bF$buf2),
    .Y(_9325_)
);

NOR2X1 _19423_ (
    .A(_9324_),
    .B(_9325_),
    .Y(_9326_)
);

AND2X2 _19424_ (
    .A(_9324_),
    .B(_9325_),
    .Y(_9327_)
);

OAI21X1 _19425_ (
    .A(_9327_),
    .B(_9326_),
    .C(_9322_),
    .Y(_9328_)
);

INVX1 _19426_ (
    .A(_9322_),
    .Y(_9329_)
);

OR2X2 _19427_ (
    .A(_9324_),
    .B(_9325_),
    .Y(_9330_)
);

OAI21X1 _19428_ (
    .A(_10869__bF$buf2),
    .B(_5315__bF$buf2),
    .C(_9324_),
    .Y(_9331_)
);

NAND3X1 _19429_ (
    .A(_9329_),
    .B(_9331_),
    .C(_9330_),
    .Y(_9332_)
);

NAND2X1 _19430_ (
    .A(areg_14_bF$buf4),
    .B(breg_22_bF$buf0),
    .Y(_9333_)
);

OAI22X1 _19431_ (
    .A(_8605_),
    .B(_9333_),
    .C(_9008_),
    .D(_9011_),
    .Y(_9335_)
);

NAND3X1 _19432_ (
    .A(_9328_),
    .B(_9332_),
    .C(_9335_),
    .Y(_9336_)
);

AOI21X1 _19433_ (
    .A(_9331_),
    .B(_9330_),
    .C(_9329_),
    .Y(_9337_)
);

NOR3X1 _19434_ (
    .A(_9322_),
    .B(_9326_),
    .C(_9327_),
    .Y(_9338_)
);

OAI21X1 _19435_ (
    .A(_2287__bF$buf0),
    .B(_3781__bF$buf3),
    .C(_8948_),
    .Y(_9339_)
);

AOI21X1 _19436_ (
    .A(_9007_),
    .B(_9339_),
    .C(_9010_),
    .Y(_9340_)
);

OAI21X1 _19437_ (
    .A(_9338_),
    .B(_9337_),
    .C(_9340_),
    .Y(_9341_)
);

NAND3X1 _19438_ (
    .A(_9321_),
    .B(_9341_),
    .C(_9336_),
    .Y(_9342_)
);

INVX1 _19439_ (
    .A(_9321_),
    .Y(_9343_)
);

NAND3X1 _19440_ (
    .A(_9340_),
    .B(_9328_),
    .C(_9332_),
    .Y(_9344_)
);

OAI21X1 _19441_ (
    .A(_9338_),
    .B(_9337_),
    .C(_9335_),
    .Y(_9346_)
);

NAND3X1 _19442_ (
    .A(_9343_),
    .B(_9344_),
    .C(_9346_),
    .Y(_9347_)
);

OAI21X1 _19443_ (
    .A(_9034_),
    .B(_9036_),
    .C(_9028_),
    .Y(_9348_)
);

NAND3X1 _19444_ (
    .A(_9342_),
    .B(_9347_),
    .C(_9348_),
    .Y(_9349_)
);

AOI21X1 _19445_ (
    .A(_9344_),
    .B(_9346_),
    .C(_9343_),
    .Y(_9350_)
);

AOI21X1 _19446_ (
    .A(_9341_),
    .B(_9336_),
    .C(_9321_),
    .Y(_9351_)
);

AOI21X1 _19447_ (
    .A(_9032_),
    .B(_9013_),
    .C(_9035_),
    .Y(_9352_)
);

OAI21X1 _19448_ (
    .A(_9351_),
    .B(_9350_),
    .C(_9352_),
    .Y(_9353_)
);

NAND3X1 _19449_ (
    .A(_9320_),
    .B(_9353_),
    .C(_9349_),
    .Y(_9354_)
);

INVX2 _19450_ (
    .A(_9320_),
    .Y(_9355_)
);

NOR3X1 _19451_ (
    .A(_9351_),
    .B(_9350_),
    .C(_9352_),
    .Y(_9357_)
);

AOI21X1 _19452_ (
    .A(_9342_),
    .B(_9347_),
    .C(_9348_),
    .Y(_9358_)
);

OAI21X1 _19453_ (
    .A(_9357_),
    .B(_9358_),
    .C(_9355_),
    .Y(_9359_)
);

NAND3X1 _19454_ (
    .A(_9319_),
    .B(_9354_),
    .C(_9359_),
    .Y(_9360_)
);

NAND2X1 _19455_ (
    .A(_8959_),
    .B(_8964_),
    .Y(_9361_)
);

NOR2X1 _19456_ (
    .A(_8971_),
    .B(_9361_),
    .Y(_9362_)
);

AOI21X1 _19457_ (
    .A(_8935_),
    .B(_8973_),
    .C(_9362_),
    .Y(_9363_)
);

NAND3X1 _19458_ (
    .A(_9342_),
    .B(_9347_),
    .C(_9352_),
    .Y(_9364_)
);

OAI21X1 _19459_ (
    .A(_9351_),
    .B(_9350_),
    .C(_9348_),
    .Y(_9365_)
);

AOI21X1 _19460_ (
    .A(_9365_),
    .B(_9364_),
    .C(_9355_),
    .Y(_9366_)
);

AOI21X1 _19461_ (
    .A(_9353_),
    .B(_9349_),
    .C(_9320_),
    .Y(_9368_)
);

OAI21X1 _19462_ (
    .A(_9366_),
    .B(_9368_),
    .C(_9363_),
    .Y(_9369_)
);

NAND3X1 _19463_ (
    .A(_9369_),
    .B(_9360_),
    .C(_9317_),
    .Y(_9370_)
);

NAND2X1 _19464_ (
    .A(_9316_),
    .B(_9313_),
    .Y(_9371_)
);

OAI21X1 _19465_ (
    .A(_9366_),
    .B(_9368_),
    .C(_9319_),
    .Y(_9372_)
);

NAND3X1 _19466_ (
    .A(_9354_),
    .B(_9359_),
    .C(_9363_),
    .Y(_9373_)
);

NAND3X1 _19467_ (
    .A(_9371_),
    .B(_9372_),
    .C(_9373_),
    .Y(_9374_)
);

OAI21X1 _19468_ (
    .A(_9090_),
    .B(_9091_),
    .C(_9088_),
    .Y(_9375_)
);

NAND3X1 _19469_ (
    .A(_9374_),
    .B(_9375_),
    .C(_9370_),
    .Y(_9376_)
);

AOI21X1 _19470_ (
    .A(_9372_),
    .B(_9373_),
    .C(_9371_),
    .Y(_9377_)
);

AOI21X1 _19471_ (
    .A(_9369_),
    .B(_9360_),
    .C(_9317_),
    .Y(_9379_)
);

AOI21X1 _19472_ (
    .A(_9006_),
    .B(_9084_),
    .C(_9093_),
    .Y(_9380_)
);

OAI21X1 _19473_ (
    .A(_9377_),
    .B(_9379_),
    .C(_9380_),
    .Y(_9381_)
);

NAND3X1 _19474_ (
    .A(_9277_),
    .B(_9376_),
    .C(_9381_),
    .Y(_9382_)
);

AND2X2 _19475_ (
    .A(_8985_),
    .B(_8979_),
    .Y(_9383_)
);

NAND3X1 _19476_ (
    .A(_9374_),
    .B(_9380_),
    .C(_9370_),
    .Y(_9384_)
);

OAI21X1 _19477_ (
    .A(_9377_),
    .B(_9379_),
    .C(_9375_),
    .Y(_9385_)
);

NAND3X1 _19478_ (
    .A(_9383_),
    .B(_9384_),
    .C(_9385_),
    .Y(_9386_)
);

NAND2X1 _19479_ (
    .A(_9382_),
    .B(_9386_),
    .Y(_9387_)
);

AOI21X1 _19480_ (
    .A(_9202_),
    .B(_9199_),
    .C(_9096_),
    .Y(_9388_)
);

OAI21X1 _19481_ (
    .A(_9095_),
    .B(_9388_),
    .C(_9209_),
    .Y(_9390_)
);

NAND2X1 _19482_ (
    .A(_9080_),
    .B(_9085_),
    .Y(_9391_)
);

NOR2X1 _19483_ (
    .A(_549__bF$buf1),
    .B(_5369_),
    .Y(_9392_)
);

INVX2 _19484_ (
    .A(_9392_),
    .Y(_9393_)
);

NAND2X1 _19485_ (
    .A(areg_15_bF$buf2),
    .B(breg_21_bF$buf0),
    .Y(_9394_)
);

NOR2X1 _19486_ (
    .A(_9333_),
    .B(_9394_),
    .Y(_9395_)
);

AND2X2 _19487_ (
    .A(_9333_),
    .B(_9394_),
    .Y(_9396_)
);

NOR2X1 _19488_ (
    .A(_9395_),
    .B(_9396_),
    .Y(_9397_)
);

XNOR2X1 _19489_ (
    .A(_9397_),
    .B(_9393_),
    .Y(_9398_)
);

OAI21X1 _19490_ (
    .A(_9025_),
    .B(_9015_),
    .C(_9020_),
    .Y(_9399_)
);

NAND2X1 _19491_ (
    .A(areg_16_bF$buf5),
    .B(breg_20_bF$buf1),
    .Y(_9401_)
);

INVX2 _19492_ (
    .A(_9401_),
    .Y(_9402_)
);

AND2X2 _19493_ (
    .A(areg_17_bF$buf5),
    .B(breg_19_bF$buf0),
    .Y(_9403_)
);

AND2X2 _19494_ (
    .A(areg_18_bF$buf0),
    .B(breg_18_bF$buf5),
    .Y(_9404_)
);

NAND2X1 _19495_ (
    .A(_9403_),
    .B(_9404_),
    .Y(_9405_)
);

OAI22X1 _19496_ (
    .A(_2884__bF$buf0),
    .B(_3253__bF$buf1),
    .C(_3146__bF$buf1),
    .D(_3529__bF$buf0),
    .Y(_9406_)
);

NAND3X1 _19497_ (
    .A(_9402_),
    .B(_9406_),
    .C(_9405_),
    .Y(_9407_)
);

NAND2X1 _19498_ (
    .A(areg_18_bF$buf5),
    .B(breg_19_bF$buf5),
    .Y(_9408_)
);

NOR2X1 _19499_ (
    .A(_9023_),
    .B(_9408_),
    .Y(_9409_)
);

NOR2X1 _19500_ (
    .A(_9403_),
    .B(_9404_),
    .Y(_9410_)
);

OAI21X1 _19501_ (
    .A(_9410_),
    .B(_9409_),
    .C(_9401_),
    .Y(_9412_)
);

NAND3X1 _19502_ (
    .A(_9407_),
    .B(_9399_),
    .C(_9412_),
    .Y(_9413_)
);

AOI21X1 _19503_ (
    .A(_9017_),
    .B(_9021_),
    .C(_9024_),
    .Y(_9414_)
);

NOR3X1 _19504_ (
    .A(_9401_),
    .B(_9409_),
    .C(_9410_),
    .Y(_9415_)
);

AOI21X1 _19505_ (
    .A(_9406_),
    .B(_9405_),
    .C(_9402_),
    .Y(_9416_)
);

OAI21X1 _19506_ (
    .A(_9415_),
    .B(_9416_),
    .C(_9414_),
    .Y(_9417_)
);

NAND3X1 _19507_ (
    .A(_9413_),
    .B(_9417_),
    .C(_9398_),
    .Y(_9418_)
);

XNOR2X1 _19508_ (
    .A(_9397_),
    .B(_9392_),
    .Y(_9419_)
);

NOR3X1 _19509_ (
    .A(_9414_),
    .B(_9416_),
    .C(_9415_),
    .Y(_9420_)
);

AOI21X1 _19510_ (
    .A(_9407_),
    .B(_9412_),
    .C(_9399_),
    .Y(_9421_)
);

OAI21X1 _19511_ (
    .A(_9420_),
    .B(_9421_),
    .C(_9419_),
    .Y(_9423_)
);

NAND2X1 _19512_ (
    .A(_9418_),
    .B(_9423_),
    .Y(_9424_)
);

OAI21X1 _19513_ (
    .A(_9075_),
    .B(_9042_),
    .C(_9067_),
    .Y(_9425_)
);

AND2X2 _19514_ (
    .A(breg_16_bF$buf0),
    .B(areg_20_bF$buf4),
    .Y(_9426_)
);

AOI21X1 _19515_ (
    .A(_8641_),
    .B(_9426_),
    .C(_9057_),
    .Y(_9427_)
);

NAND2X1 _19516_ (
    .A(breg_17_bF$buf4),
    .B(areg_19_bF$buf2),
    .Y(_9428_)
);

INVX1 _19517_ (
    .A(_9428_),
    .Y(_9429_)
);

AND2X2 _19518_ (
    .A(breg_15_bF$buf0),
    .B(areg_21_bF$buf1),
    .Y(_9430_)
);

NAND2X1 _19519_ (
    .A(_9426_),
    .B(_9430_),
    .Y(_9431_)
);

NAND2X1 _19520_ (
    .A(breg_16_bF$buf5),
    .B(areg_20_bF$buf3),
    .Y(_9432_)
);

OAI21X1 _19521_ (
    .A(_2362__bF$buf2),
    .B(_3961__bF$buf3),
    .C(_9432_),
    .Y(_9434_)
);

NAND3X1 _19522_ (
    .A(_9429_),
    .B(_9434_),
    .C(_9431_),
    .Y(_9435_)
);

OAI21X1 _19523_ (
    .A(_2560__bF$buf4),
    .B(_3958__bF$buf0),
    .C(_9430_),
    .Y(_9436_)
);

OAI21X1 _19524_ (
    .A(_2362__bF$buf1),
    .B(_3961__bF$buf2),
    .C(_9426_),
    .Y(_9437_)
);

NAND3X1 _19525_ (
    .A(_9428_),
    .B(_9436_),
    .C(_9437_),
    .Y(_9438_)
);

NOR2X1 _19526_ (
    .A(_9059_),
    .B(_9100_),
    .Y(_9439_)
);

OAI21X1 _19527_ (
    .A(_2586__bF$buf0),
    .B(_4541__bF$buf3),
    .C(_9059_),
    .Y(_9440_)
);

AOI21X1 _19528_ (
    .A(_9099_),
    .B(_9440_),
    .C(_9439_),
    .Y(_9441_)
);

NAND3X1 _19529_ (
    .A(_9441_),
    .B(_9435_),
    .C(_9438_),
    .Y(_9442_)
);

AOI21X1 _19530_ (
    .A(_9436_),
    .B(_9437_),
    .C(_9428_),
    .Y(_9443_)
);

AOI21X1 _19531_ (
    .A(_9434_),
    .B(_9431_),
    .C(_9429_),
    .Y(_9445_)
);

NAND2X1 _19532_ (
    .A(breg_13_bF$buf1),
    .B(areg_23_bF$buf3),
    .Y(_9446_)
);

AND2X2 _19533_ (
    .A(_9059_),
    .B(_9100_),
    .Y(_9447_)
);

OAI22X1 _19534_ (
    .A(_8699_),
    .B(_9446_),
    .C(_9447_),
    .D(_9098_),
    .Y(_9448_)
);

OAI21X1 _19535_ (
    .A(_9443_),
    .B(_9445_),
    .C(_9448_),
    .Y(_9449_)
);

AOI21X1 _19536_ (
    .A(_9442_),
    .B(_9449_),
    .C(_9427_),
    .Y(_9450_)
);

OAI21X1 _19537_ (
    .A(_9065_),
    .B(_9432_),
    .C(_9048_),
    .Y(_9451_)
);

NAND3X1 _19538_ (
    .A(_9435_),
    .B(_9438_),
    .C(_9448_),
    .Y(_9452_)
);

OAI21X1 _19539_ (
    .A(_9443_),
    .B(_9445_),
    .C(_9441_),
    .Y(_9453_)
);

AOI21X1 _19540_ (
    .A(_9452_),
    .B(_9453_),
    .C(_9451_),
    .Y(_9454_)
);

OAI21X1 _19541_ (
    .A(_9450_),
    .B(_9454_),
    .C(_9425_),
    .Y(_9456_)
);

AOI21X1 _19542_ (
    .A(_9066_),
    .B(_9068_),
    .C(_9074_),
    .Y(_9457_)
);

NAND3X1 _19543_ (
    .A(_9451_),
    .B(_9452_),
    .C(_9453_),
    .Y(_9458_)
);

NOR3X1 _19544_ (
    .A(_9445_),
    .B(_9441_),
    .C(_9443_),
    .Y(_9459_)
);

AOI21X1 _19545_ (
    .A(_9435_),
    .B(_9438_),
    .C(_9448_),
    .Y(_9460_)
);

OAI21X1 _19546_ (
    .A(_9459_),
    .B(_9460_),
    .C(_9427_),
    .Y(_9461_)
);

NAND3X1 _19547_ (
    .A(_9457_),
    .B(_9458_),
    .C(_9461_),
    .Y(_9462_)
);

AOI21X1 _19548_ (
    .A(_9456_),
    .B(_9462_),
    .C(_9424_),
    .Y(_9463_)
);

AND2X2 _19549_ (
    .A(_9423_),
    .B(_9418_),
    .Y(_9464_)
);

NAND3X1 _19550_ (
    .A(_9425_),
    .B(_9458_),
    .C(_9461_),
    .Y(_9465_)
);

OAI21X1 _19551_ (
    .A(_9450_),
    .B(_9454_),
    .C(_9457_),
    .Y(_9467_)
);

AOI21X1 _19552_ (
    .A(_9465_),
    .B(_9467_),
    .C(_9464_),
    .Y(_9468_)
);

AOI21X1 _19553_ (
    .A(_9097_),
    .B(_9130_),
    .C(_9139_),
    .Y(_9469_)
);

OAI21X1 _19554_ (
    .A(_9468_),
    .B(_9463_),
    .C(_9469_),
    .Y(_9470_)
);

NAND3X1 _19555_ (
    .A(_9465_),
    .B(_9467_),
    .C(_9464_),
    .Y(_9471_)
);

NAND3X1 _19556_ (
    .A(_9456_),
    .B(_9424_),
    .C(_9462_),
    .Y(_9472_)
);

OAI21X1 _19557_ (
    .A(_9138_),
    .B(_9136_),
    .C(_9134_),
    .Y(_9473_)
);

NAND3X1 _19558_ (
    .A(_9472_),
    .B(_9473_),
    .C(_9471_),
    .Y(_9474_)
);

NAND3X1 _19559_ (
    .A(_9391_),
    .B(_9474_),
    .C(_9470_),
    .Y(_9475_)
);

AND2X2 _19560_ (
    .A(_9085_),
    .B(_9080_),
    .Y(_9476_)
);

AOI21X1 _19561_ (
    .A(_9472_),
    .B(_9471_),
    .C(_9473_),
    .Y(_9478_)
);

NOR3X1 _19562_ (
    .A(_9468_),
    .B(_9463_),
    .C(_9469_),
    .Y(_9479_)
);

OAI21X1 _19563_ (
    .A(_9479_),
    .B(_9478_),
    .C(_9476_),
    .Y(_9480_)
);

NAND2X1 _19564_ (
    .A(_9475_),
    .B(_9480_),
    .Y(_9481_)
);

OAI21X1 _19565_ (
    .A(_9141_),
    .B(_9201_),
    .C(_9194_),
    .Y(_9482_)
);

NAND2X1 _19566_ (
    .A(_9125_),
    .B(_9131_),
    .Y(_9483_)
);

NAND2X1 _19567_ (
    .A(breg_14_bF$buf3),
    .B(areg_22_bF$buf1),
    .Y(_9484_)
);

NAND2X1 _19568_ (
    .A(breg_12_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_9485_)
);

XOR2X1 _19569_ (
    .A(_9446_),
    .B(_9485_),
    .Y(_9486_)
);

XNOR2X1 _19570_ (
    .A(_9486_),
    .B(_9484_),
    .Y(_9487_)
);

OAI21X1 _19571_ (
    .A(_9111_),
    .B(_9106_),
    .C(_9114_),
    .Y(_9489_)
);

NAND2X1 _19572_ (
    .A(breg_11_bF$buf1),
    .B(areg_25_bF$buf4),
    .Y(_9490_)
);

INVX2 _19573_ (
    .A(_9490_),
    .Y(_9491_)
);

AND2X2 _19574_ (
    .A(breg_10_bF$buf5),
    .B(areg_26_bF$buf4),
    .Y(_9492_)
);

AND2X2 _19575_ (
    .A(breg_9_bF$buf3),
    .B(areg_27_bF$buf3),
    .Y(_9493_)
);

NAND2X1 _19576_ (
    .A(_9492_),
    .B(_9493_),
    .Y(_9494_)
);

OAI21X1 _19577_ (
    .A(_6044__bF$buf5),
    .B(_7100__bF$buf2),
    .C(_9107_),
    .Y(_9495_)
);

NAND3X1 _19578_ (
    .A(_9491_),
    .B(_9495_),
    .C(_9494_),
    .Y(_9496_)
);

NAND2X1 _19579_ (
    .A(breg_9_bF$buf2),
    .B(areg_27_bF$buf2),
    .Y(_9497_)
);

NOR2X1 _19580_ (
    .A(_9107_),
    .B(_9497_),
    .Y(_9498_)
);

NOR2X1 _19581_ (
    .A(_9492_),
    .B(_9493_),
    .Y(_9500_)
);

OAI21X1 _19582_ (
    .A(_9500_),
    .B(_9498_),
    .C(_9490_),
    .Y(_9501_)
);

NAND3X1 _19583_ (
    .A(_9496_),
    .B(_9489_),
    .C(_9501_),
    .Y(_9502_)
);

AOI21X1 _19584_ (
    .A(_9113_),
    .B(_9116_),
    .C(_9108_),
    .Y(_9503_)
);

OAI21X1 _19585_ (
    .A(_7217__bF$buf3),
    .B(_6686__bF$buf2),
    .C(_9493_),
    .Y(_9504_)
);

OAI21X1 _19586_ (
    .A(_6044__bF$buf4),
    .B(_7100__bF$buf1),
    .C(_9492_),
    .Y(_9505_)
);

AOI21X1 _19587_ (
    .A(_9504_),
    .B(_9505_),
    .C(_9490_),
    .Y(_9506_)
);

AOI21X1 _19588_ (
    .A(_9495_),
    .B(_9494_),
    .C(_9491_),
    .Y(_9507_)
);

OAI21X1 _19589_ (
    .A(_9506_),
    .B(_9507_),
    .C(_9503_),
    .Y(_9508_)
);

NAND3X1 _19590_ (
    .A(_9502_),
    .B(_9508_),
    .C(_9487_),
    .Y(_9509_)
);

INVX2 _19591_ (
    .A(_9484_),
    .Y(_9511_)
);

XNOR2X1 _19592_ (
    .A(_9486_),
    .B(_9511_),
    .Y(_9512_)
);

OAI21X1 _19593_ (
    .A(_9506_),
    .B(_9507_),
    .C(_9489_),
    .Y(_9513_)
);

NAND3X1 _19594_ (
    .A(_9503_),
    .B(_9496_),
    .C(_9501_),
    .Y(_9514_)
);

NAND3X1 _19595_ (
    .A(_9513_),
    .B(_9514_),
    .C(_9512_),
    .Y(_9515_)
);

OAI21X1 _19596_ (
    .A(_9179_),
    .B(_9143_),
    .C(_9169_),
    .Y(_9516_)
);

NAND3X1 _19597_ (
    .A(_9516_),
    .B(_9509_),
    .C(_9515_),
    .Y(_9517_)
);

AOI21X1 _19598_ (
    .A(_9513_),
    .B(_9514_),
    .C(_9512_),
    .Y(_9518_)
);

AOI21X1 _19599_ (
    .A(_9502_),
    .B(_9508_),
    .C(_9487_),
    .Y(_9519_)
);

AOI21X1 _19600_ (
    .A(_9168_),
    .B(_9171_),
    .C(_9178_),
    .Y(_9520_)
);

OAI21X1 _19601_ (
    .A(_9518_),
    .B(_9519_),
    .C(_9520_),
    .Y(_9522_)
);

NAND3X1 _19602_ (
    .A(_9483_),
    .B(_9517_),
    .C(_9522_),
    .Y(_9523_)
);

AND2X2 _19603_ (
    .A(_9131_),
    .B(_9125_),
    .Y(_9524_)
);

NAND3X1 _19604_ (
    .A(_9520_),
    .B(_9509_),
    .C(_9515_),
    .Y(_9525_)
);

OAI21X1 _19605_ (
    .A(_9518_),
    .B(_9519_),
    .C(_9516_),
    .Y(_9526_)
);

NAND3X1 _19606_ (
    .A(_9525_),
    .B(_9526_),
    .C(_9524_),
    .Y(_9527_)
);

NAND2X1 _19607_ (
    .A(_9523_),
    .B(_9527_),
    .Y(_9528_)
);

AOI21X1 _19608_ (
    .A(_9142_),
    .B(_9146_),
    .C(_9161_),
    .Y(_9529_)
);

NOR2X1 _19609_ (
    .A(_8369_),
    .B(_9173_),
    .Y(_9530_)
);

INVX2 _19610_ (
    .A(_9530_),
    .Y(_9531_)
);

NAND2X1 _19611_ (
    .A(breg[8]),
    .B(areg_28_bF$buf3),
    .Y(_9533_)
);

INVX1 _19612_ (
    .A(_9533_),
    .Y(_9534_)
);

AND2X2 _19613_ (
    .A(breg_7_bF$buf2),
    .B(areg_30_bF$buf0),
    .Y(_9535_)
);

NAND2X1 _19614_ (
    .A(_9146_),
    .B(_9535_),
    .Y(_9536_)
);

NAND2X1 _19615_ (
    .A(breg_7_bF$buf1),
    .B(areg_29_bF$buf1),
    .Y(_9537_)
);

OAI21X1 _19616_ (
    .A(_5453__bF$buf4),
    .B(_8759_),
    .C(_9537_),
    .Y(_9538_)
);

NAND3X1 _19617_ (
    .A(_9534_),
    .B(_9538_),
    .C(_9536_),
    .Y(_9539_)
);

NAND3X1 _19618_ (
    .A(breg_6_bF$buf2),
    .B(areg_30_bF$buf5),
    .C(_9537_),
    .Y(_9540_)
);

NAND2X1 _19619_ (
    .A(breg_6_bF$buf1),
    .B(areg_30_bF$buf4),
    .Y(_9541_)
);

NAND3X1 _19620_ (
    .A(breg_7_bF$buf0),
    .B(areg_29_bF$buf0),
    .C(_9541_),
    .Y(_9542_)
);

NAND3X1 _19621_ (
    .A(_9533_),
    .B(_9540_),
    .C(_9542_),
    .Y(_9544_)
);

NAND3X1 _19622_ (
    .A(_9531_),
    .B(_9544_),
    .C(_9539_),
    .Y(_9545_)
);

AOI21X1 _19623_ (
    .A(_9540_),
    .B(_9542_),
    .C(_9533_),
    .Y(_9546_)
);

AOI21X1 _19624_ (
    .A(_9538_),
    .B(_9536_),
    .C(_9534_),
    .Y(_9547_)
);

OAI21X1 _19625_ (
    .A(_9547_),
    .B(_9546_),
    .C(_9530_),
    .Y(_9548_)
);

AOI21X1 _19626_ (
    .A(_9545_),
    .B(_9548_),
    .C(_9529_),
    .Y(_9549_)
);

OAI21X1 _19627_ (
    .A(_9167_),
    .B(_9149_),
    .C(_9151_),
    .Y(_9550_)
);

NAND3X1 _19628_ (
    .A(_9530_),
    .B(_9544_),
    .C(_9539_),
    .Y(_9551_)
);

OAI21X1 _19629_ (
    .A(_9547_),
    .B(_9546_),
    .C(_9531_),
    .Y(_9552_)
);

AOI21X1 _19630_ (
    .A(_9551_),
    .B(_9552_),
    .C(_9550_),
    .Y(_9553_)
);

NOR3X1 _19631_ (
    .A(_9549_),
    .B(_9173_),
    .C(_9553_),
    .Y(_9555_)
);

INVX1 _19632_ (
    .A(_9173_),
    .Y(_9556_)
);

NAND3X1 _19633_ (
    .A(_9550_),
    .B(_9551_),
    .C(_9552_),
    .Y(_9557_)
);

NOR3X1 _19634_ (
    .A(_9546_),
    .B(_9531_),
    .C(_9547_),
    .Y(_9558_)
);

AOI21X1 _19635_ (
    .A(_9544_),
    .B(_9539_),
    .C(_9530_),
    .Y(_9559_)
);

OAI21X1 _19636_ (
    .A(_9558_),
    .B(_9559_),
    .C(_9529_),
    .Y(_9560_)
);

AOI21X1 _19637_ (
    .A(_9557_),
    .B(_9560_),
    .C(_9556_),
    .Y(_9561_)
);

OAI21X1 _19638_ (
    .A(_9555_),
    .B(_9561_),
    .C(_9183_),
    .Y(_9562_)
);

NOR3X1 _19639_ (
    .A(_9166_),
    .B(_9175_),
    .C(_9172_),
    .Y(_9563_)
);

NAND3X1 _19640_ (
    .A(_9556_),
    .B(_9557_),
    .C(_9560_),
    .Y(_9564_)
);

OAI21X1 _19641_ (
    .A(_9549_),
    .B(_9553_),
    .C(_9173_),
    .Y(_9566_)
);

NAND3X1 _19642_ (
    .A(_9564_),
    .B(_9566_),
    .C(_9563_),
    .Y(_9567_)
);

NAND2X1 _19643_ (
    .A(_9567_),
    .B(_9562_),
    .Y(_9568_)
);

NOR2X1 _19644_ (
    .A(_9528_),
    .B(_9568_),
    .Y(_9569_)
);

AND2X2 _19645_ (
    .A(_9568_),
    .B(_9528_),
    .Y(_9570_)
);

OAI21X1 _19646_ (
    .A(_9570_),
    .B(_9569_),
    .C(_9482_),
    .Y(_9571_)
);

AOI21X1 _19647_ (
    .A(_9195_),
    .B(_9191_),
    .C(_9200_),
    .Y(_9572_)
);

OR2X2 _19648_ (
    .A(_9568_),
    .B(_9528_),
    .Y(_9573_)
);

NAND2X1 _19649_ (
    .A(_9528_),
    .B(_9568_),
    .Y(_9574_)
);

NAND3X1 _19650_ (
    .A(_9574_),
    .B(_9573_),
    .C(_9572_),
    .Y(_9575_)
);

AOI21X1 _19651_ (
    .A(_9571_),
    .B(_9575_),
    .C(_9481_),
    .Y(_9577_)
);

OAI21X1 _19652_ (
    .A(_9479_),
    .B(_9478_),
    .C(_9391_),
    .Y(_9578_)
);

NAND3X1 _19653_ (
    .A(_9474_),
    .B(_9470_),
    .C(_9476_),
    .Y(_9579_)
);

NAND2X1 _19654_ (
    .A(_9579_),
    .B(_9578_),
    .Y(_9580_)
);

NAND3X1 _19655_ (
    .A(_9574_),
    .B(_9573_),
    .C(_9482_),
    .Y(_9581_)
);

OAI21X1 _19656_ (
    .A(_9570_),
    .B(_9569_),
    .C(_9572_),
    .Y(_9582_)
);

AOI21X1 _19657_ (
    .A(_9582_),
    .B(_9581_),
    .C(_9580_),
    .Y(_9583_)
);

OAI21X1 _19658_ (
    .A(_9577_),
    .B(_9583_),
    .C(_9390_),
    .Y(_9584_)
);

NOR3X1 _19659_ (
    .A(_9188_),
    .B(_9196_),
    .C(_9198_),
    .Y(_9585_)
);

AOI21X1 _19660_ (
    .A(_9210_),
    .B(_9208_),
    .C(_9585_),
    .Y(_9586_)
);

NAND3X1 _19661_ (
    .A(_9581_),
    .B(_9582_),
    .C(_9580_),
    .Y(_9588_)
);

NAND3X1 _19662_ (
    .A(_9571_),
    .B(_9575_),
    .C(_9481_),
    .Y(_9589_)
);

NAND3X1 _19663_ (
    .A(_9588_),
    .B(_9589_),
    .C(_9586_),
    .Y(_9590_)
);

AOI21X1 _19664_ (
    .A(_9590_),
    .B(_9584_),
    .C(_9387_),
    .Y(_9591_)
);

NAND3X1 _19665_ (
    .A(_9383_),
    .B(_9376_),
    .C(_9381_),
    .Y(_9592_)
);

NAND3X1 _19666_ (
    .A(_9277_),
    .B(_9384_),
    .C(_9385_),
    .Y(_9593_)
);

NAND2X1 _19667_ (
    .A(_9593_),
    .B(_9592_),
    .Y(_9594_)
);

NAND3X1 _19668_ (
    .A(_9588_),
    .B(_9589_),
    .C(_9390_),
    .Y(_9595_)
);

OAI21X1 _19669_ (
    .A(_9577_),
    .B(_9583_),
    .C(_9586_),
    .Y(_9596_)
);

AOI21X1 _19670_ (
    .A(_9595_),
    .B(_9596_),
    .C(_9594_),
    .Y(_9597_)
);

OAI21X1 _19671_ (
    .A(_9591_),
    .B(_9597_),
    .C(_9276_),
    .Y(_9599_)
);

NOR3X1 _19672_ (
    .A(_9205_),
    .B(_9211_),
    .C(_9215_),
    .Y(_9600_)
);

AOI21X1 _19673_ (
    .A(_9224_),
    .B(_9222_),
    .C(_9600_),
    .Y(_9601_)
);

NAND3X1 _19674_ (
    .A(_9595_),
    .B(_9596_),
    .C(_9594_),
    .Y(_9602_)
);

NAND3X1 _19675_ (
    .A(_9590_),
    .B(_9584_),
    .C(_9387_),
    .Y(_9603_)
);

NAND3X1 _19676_ (
    .A(_9602_),
    .B(_9603_),
    .C(_9601_),
    .Y(_9604_)
);

AOI21X1 _19677_ (
    .A(_9604_),
    .B(_9599_),
    .C(_9274_),
    .Y(_9605_)
);

NAND3X1 _19678_ (
    .A(_9276_),
    .B(_9602_),
    .C(_9603_),
    .Y(_9606_)
);

OAI21X1 _19679_ (
    .A(_9591_),
    .B(_9597_),
    .C(_9601_),
    .Y(_9607_)
);

AOI21X1 _19680_ (
    .A(_9606_),
    .B(_9607_),
    .C(_9273_),
    .Y(_9608_)
);

OAI21X1 _19681_ (
    .A(_9605_),
    .B(_9608_),
    .C(_9272_),
    .Y(_9610_)
);

NOR3X1 _19682_ (
    .A(_9219_),
    .B(_9226_),
    .C(_9229_),
    .Y(_9611_)
);

AOI21X1 _19683_ (
    .A(_8887_),
    .B(_9235_),
    .C(_9611_),
    .Y(_9612_)
);

NAND3X1 _19684_ (
    .A(_9273_),
    .B(_9606_),
    .C(_9607_),
    .Y(_9613_)
);

NOR3X1 _19685_ (
    .A(_9591_),
    .B(_9597_),
    .C(_9601_),
    .Y(_9614_)
);

AOI21X1 _19686_ (
    .A(_9602_),
    .B(_9603_),
    .C(_9276_),
    .Y(_9615_)
);

OAI21X1 _19687_ (
    .A(_9614_),
    .B(_9615_),
    .C(_9274_),
    .Y(_9616_)
);

NAND3X1 _19688_ (
    .A(_9612_),
    .B(_9613_),
    .C(_9616_),
    .Y(_9617_)
);

AOI21X1 _19689_ (
    .A(_9610_),
    .B(_9617_),
    .C(_9270_),
    .Y(_9618_)
);

NAND3X1 _19690_ (
    .A(_9272_),
    .B(_9613_),
    .C(_9616_),
    .Y(_9619_)
);

OAI21X1 _19691_ (
    .A(_9605_),
    .B(_9608_),
    .C(_9612_),
    .Y(_9621_)
);

AOI21X1 _19692_ (
    .A(_9621_),
    .B(_9619_),
    .C(_9269_),
    .Y(_9622_)
);

OAI21X1 _19693_ (
    .A(_9618_),
    .B(_9622_),
    .C(_9267_),
    .Y(_9623_)
);

NOR3X1 _19694_ (
    .A(_9233_),
    .B(_9237_),
    .C(_9240_),
    .Y(_9624_)
);

AOI21X1 _19695_ (
    .A(_8882_),
    .B(_9246_),
    .C(_9624_),
    .Y(_9625_)
);

NAND3X1 _19696_ (
    .A(_9269_),
    .B(_9621_),
    .C(_9619_),
    .Y(_9626_)
);

NAND3X1 _19697_ (
    .A(_9270_),
    .B(_9610_),
    .C(_9617_),
    .Y(_9627_)
);

NAND3X1 _19698_ (
    .A(_9626_),
    .B(_9627_),
    .C(_9625_),
    .Y(_9628_)
);

NAND2X1 _19699_ (
    .A(_9628_),
    .B(_9623_),
    .Y(_9629_)
);

INVX2 _19700_ (
    .A(_9629_),
    .Y(_9630_)
);

XNOR2X1 _19701_ (
    .A(_9265_),
    .B(_9630_),
    .Y(_0_[36])
);

INVX1 _19702_ (
    .A(_9265_),
    .Y(_9632_)
);

NAND3X1 _19703_ (
    .A(_9267_),
    .B(_9626_),
    .C(_9627_),
    .Y(_9633_)
);

OAI21X1 _19704_ (
    .A(_9632_),
    .B(_9630_),
    .C(_9633_),
    .Y(_9634_)
);

AOI21X1 _19705_ (
    .A(_9613_),
    .B(_9616_),
    .C(_9272_),
    .Y(_9635_)
);

OAI21X1 _19706_ (
    .A(_9635_),
    .B(_9270_),
    .C(_9619_),
    .Y(_9636_)
);

OAI21X1 _19707_ (
    .A(_9307_),
    .B(_9280_),
    .C(_9315_),
    .Y(_9637_)
);

INVX2 _19708_ (
    .A(_9637_),
    .Y(_9638_)
);

OAI21X1 _19709_ (
    .A(_9615_),
    .B(_9274_),
    .C(_9606_),
    .Y(_9639_)
);

NAND2X1 _19710_ (
    .A(_9376_),
    .B(_9382_),
    .Y(_9640_)
);

INVX2 _19711_ (
    .A(_9640_),
    .Y(_9642_)
);

AOI21X1 _19712_ (
    .A(_9588_),
    .B(_9589_),
    .C(_9390_),
    .Y(_9643_)
);

OAI21X1 _19713_ (
    .A(_9387_),
    .B(_9643_),
    .C(_9595_),
    .Y(_9644_)
);

NAND2X1 _19714_ (
    .A(_9360_),
    .B(_9370_),
    .Y(_9645_)
);

NOR2X1 _19715_ (
    .A(_3646__bF$buf0),
    .B(_7225__bF$buf3),
    .Y(_9646_)
);

INVX1 _19716_ (
    .A(_9646_),
    .Y(_9647_)
);

OAI21X1 _19717_ (
    .A(_9297_),
    .B(_9283_),
    .C(_9305_),
    .Y(_9648_)
);

NOR2X1 _19718_ (
    .A(_4434__bF$buf2),
    .B(_6815__bF$buf2),
    .Y(_9649_)
);

INVX2 _19719_ (
    .A(_9649_),
    .Y(_9650_)
);

OAI21X1 _19720_ (
    .A(_9295_),
    .B(_9285_),
    .C(_9289_),
    .Y(_9651_)
);

NAND2X1 _19721_ (
    .A(areg_8_bF$buf0),
    .B(breg_29_bF$buf1),
    .Y(_9653_)
);

INVX2 _19722_ (
    .A(_9653_),
    .Y(_9654_)
);

AND2X2 _19723_ (
    .A(areg_9_bF$buf0),
    .B(breg_28_bF$buf4),
    .Y(_9655_)
);

AND2X2 _19724_ (
    .A(areg_10_bF$buf0),
    .B(breg_27_bF$buf4),
    .Y(_9656_)
);

NAND2X1 _19725_ (
    .A(_9655_),
    .B(_9656_),
    .Y(_9657_)
);

OAI22X1 _19726_ (
    .A(_6582__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_7711__bF$buf3),
    .D(_5668__bF$buf3),
    .Y(_9658_)
);

NAND3X1 _19727_ (
    .A(_9654_),
    .B(_9658_),
    .C(_9657_),
    .Y(_9659_)
);

NAND2X1 _19728_ (
    .A(areg_10_bF$buf4),
    .B(breg_28_bF$buf3),
    .Y(_9660_)
);

NOR2X1 _19729_ (
    .A(_9293_),
    .B(_9660_),
    .Y(_9661_)
);

NOR2X1 _19730_ (
    .A(_9655_),
    .B(_9656_),
    .Y(_9662_)
);

OAI21X1 _19731_ (
    .A(_9662_),
    .B(_9661_),
    .C(_9653_),
    .Y(_9664_)
);

AOI21X1 _19732_ (
    .A(_9659_),
    .B(_9664_),
    .C(_9651_),
    .Y(_9665_)
);

AOI21X1 _19733_ (
    .A(_9286_),
    .B(_9291_),
    .C(_9294_),
    .Y(_9666_)
);

OAI21X1 _19734_ (
    .A(_6582__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_9656_),
    .Y(_9667_)
);

OAI21X1 _19735_ (
    .A(_7711__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_9655_),
    .Y(_9668_)
);

AOI21X1 _19736_ (
    .A(_9667_),
    .B(_9668_),
    .C(_9653_),
    .Y(_9669_)
);

AOI21X1 _19737_ (
    .A(_9658_),
    .B(_9657_),
    .C(_9654_),
    .Y(_9670_)
);

NOR3X1 _19738_ (
    .A(_9670_),
    .B(_9666_),
    .C(_9669_),
    .Y(_9671_)
);

OAI21X1 _19739_ (
    .A(_9671_),
    .B(_9665_),
    .C(_9650_),
    .Y(_9672_)
);

OAI21X1 _19740_ (
    .A(_9669_),
    .B(_9670_),
    .C(_9666_),
    .Y(_9673_)
);

NAND3X1 _19741_ (
    .A(_9659_),
    .B(_9651_),
    .C(_9664_),
    .Y(_9675_)
);

NAND3X1 _19742_ (
    .A(_9649_),
    .B(_9673_),
    .C(_9675_),
    .Y(_9676_)
);

AOI21X1 _19743_ (
    .A(_9676_),
    .B(_9672_),
    .C(_9648_),
    .Y(_9677_)
);

AOI21X1 _19744_ (
    .A(_9282_),
    .B(_9304_),
    .C(_9302_),
    .Y(_9678_)
);

AOI21X1 _19745_ (
    .A(_9673_),
    .B(_9675_),
    .C(_9649_),
    .Y(_9679_)
);

NOR3X1 _19746_ (
    .A(_9665_),
    .B(_9650_),
    .C(_9671_),
    .Y(_9680_)
);

NOR3X1 _19747_ (
    .A(_9678_),
    .B(_9679_),
    .C(_9680_),
    .Y(_9681_)
);

OAI21X1 _19748_ (
    .A(_9681_),
    .B(_9677_),
    .C(_9647_),
    .Y(_9682_)
);

OAI21X1 _19749_ (
    .A(_9680_),
    .B(_9679_),
    .C(_9678_),
    .Y(_9683_)
);

NAND3X1 _19750_ (
    .A(_9648_),
    .B(_9676_),
    .C(_9672_),
    .Y(_9684_)
);

NAND3X1 _19751_ (
    .A(_9646_),
    .B(_9684_),
    .C(_9683_),
    .Y(_9686_)
);

AND2X2 _19752_ (
    .A(_9682_),
    .B(_9686_),
    .Y(_9687_)
);

OAI21X1 _19753_ (
    .A(_9355_),
    .B(_9358_),
    .C(_9349_),
    .Y(_9688_)
);

NAND2X1 _19754_ (
    .A(_9336_),
    .B(_9342_),
    .Y(_9689_)
);

OAI21X1 _19755_ (
    .A(_9327_),
    .B(_9322_),
    .C(_9330_),
    .Y(_9690_)
);

NAND2X1 _19756_ (
    .A(areg_11_bF$buf0),
    .B(breg_26_bF$buf3),
    .Y(_9691_)
);

NAND2X1 _19757_ (
    .A(areg_12_bF$buf1),
    .B(breg_25_bF$buf0),
    .Y(_9692_)
);

NAND2X1 _19758_ (
    .A(areg_13_bF$buf4),
    .B(breg_24_bF$buf1),
    .Y(_9693_)
);

NOR2X1 _19759_ (
    .A(_9692_),
    .B(_9693_),
    .Y(_9694_)
);

AND2X2 _19760_ (
    .A(_9692_),
    .B(_9693_),
    .Y(_9695_)
);

OAI21X1 _19761_ (
    .A(_9695_),
    .B(_9694_),
    .C(_9691_),
    .Y(_9697_)
);

INVX1 _19762_ (
    .A(_9691_),
    .Y(_9698_)
);

OR2X2 _19763_ (
    .A(_9692_),
    .B(_9693_),
    .Y(_9699_)
);

OAI21X1 _19764_ (
    .A(_549__bF$buf0),
    .B(_5315__bF$buf1),
    .C(_9692_),
    .Y(_9700_)
);

NAND3X1 _19765_ (
    .A(_9698_),
    .B(_9700_),
    .C(_9699_),
    .Y(_9701_)
);

NAND2X1 _19766_ (
    .A(areg_15_bF$buf1),
    .B(breg_22_bF$buf4),
    .Y(_9702_)
);

OAI22X1 _19767_ (
    .A(_9009_),
    .B(_9702_),
    .C(_9393_),
    .D(_9396_),
    .Y(_9703_)
);

NAND3X1 _19768_ (
    .A(_9697_),
    .B(_9701_),
    .C(_9703_),
    .Y(_9704_)
);

AOI21X1 _19769_ (
    .A(_9700_),
    .B(_9699_),
    .C(_9698_),
    .Y(_9705_)
);

NOR3X1 _19770_ (
    .A(_9691_),
    .B(_9694_),
    .C(_9695_),
    .Y(_9706_)
);

OAI21X1 _19771_ (
    .A(_2465__bF$buf0),
    .B(_3781__bF$buf2),
    .C(_9333_),
    .Y(_9708_)
);

AOI21X1 _19772_ (
    .A(_9392_),
    .B(_9708_),
    .C(_9395_),
    .Y(_9709_)
);

OAI21X1 _19773_ (
    .A(_9706_),
    .B(_9705_),
    .C(_9709_),
    .Y(_9710_)
);

NAND3X1 _19774_ (
    .A(_9690_),
    .B(_9710_),
    .C(_9704_),
    .Y(_9711_)
);

INVX1 _19775_ (
    .A(_9690_),
    .Y(_9712_)
);

NAND3X1 _19776_ (
    .A(_9709_),
    .B(_9697_),
    .C(_9701_),
    .Y(_9713_)
);

OAI21X1 _19777_ (
    .A(_9706_),
    .B(_9705_),
    .C(_9703_),
    .Y(_9714_)
);

NAND3X1 _19778_ (
    .A(_9712_),
    .B(_9713_),
    .C(_9714_),
    .Y(_9715_)
);

OAI21X1 _19779_ (
    .A(_9419_),
    .B(_9421_),
    .C(_9413_),
    .Y(_9716_)
);

NAND3X1 _19780_ (
    .A(_9711_),
    .B(_9715_),
    .C(_9716_),
    .Y(_9717_)
);

AOI21X1 _19781_ (
    .A(_9713_),
    .B(_9714_),
    .C(_9712_),
    .Y(_9719_)
);

AOI21X1 _19782_ (
    .A(_9710_),
    .B(_9704_),
    .C(_9690_),
    .Y(_9720_)
);

AOI21X1 _19783_ (
    .A(_9417_),
    .B(_9398_),
    .C(_9420_),
    .Y(_9721_)
);

OAI21X1 _19784_ (
    .A(_9720_),
    .B(_9719_),
    .C(_9721_),
    .Y(_9722_)
);

NAND3X1 _19785_ (
    .A(_9689_),
    .B(_9722_),
    .C(_9717_),
    .Y(_9723_)
);

AND2X2 _19786_ (
    .A(_9342_),
    .B(_9336_),
    .Y(_9724_)
);

NOR3X1 _19787_ (
    .A(_9720_),
    .B(_9719_),
    .C(_9721_),
    .Y(_9725_)
);

AOI21X1 _19788_ (
    .A(_9711_),
    .B(_9715_),
    .C(_9716_),
    .Y(_9726_)
);

OAI21X1 _19789_ (
    .A(_9725_),
    .B(_9726_),
    .C(_9724_),
    .Y(_9727_)
);

NAND3X1 _19790_ (
    .A(_9688_),
    .B(_9723_),
    .C(_9727_),
    .Y(_9728_)
);

AOI21X1 _19791_ (
    .A(_9320_),
    .B(_9353_),
    .C(_9357_),
    .Y(_9730_)
);

NAND3X1 _19792_ (
    .A(_9711_),
    .B(_9715_),
    .C(_9721_),
    .Y(_9731_)
);

OAI21X1 _19793_ (
    .A(_9720_),
    .B(_9719_),
    .C(_9716_),
    .Y(_9732_)
);

AOI21X1 _19794_ (
    .A(_9732_),
    .B(_9731_),
    .C(_9724_),
    .Y(_9733_)
);

AOI21X1 _19795_ (
    .A(_9722_),
    .B(_9717_),
    .C(_9689_),
    .Y(_9734_)
);

OAI21X1 _19796_ (
    .A(_9733_),
    .B(_9734_),
    .C(_9730_),
    .Y(_9735_)
);

NAND3X1 _19797_ (
    .A(_9735_),
    .B(_9728_),
    .C(_9687_),
    .Y(_9736_)
);

NAND2X1 _19798_ (
    .A(_9686_),
    .B(_9682_),
    .Y(_9737_)
);

OAI21X1 _19799_ (
    .A(_9733_),
    .B(_9734_),
    .C(_9688_),
    .Y(_9738_)
);

NAND3X1 _19800_ (
    .A(_9730_),
    .B(_9723_),
    .C(_9727_),
    .Y(_9739_)
);

NAND3X1 _19801_ (
    .A(_9737_),
    .B(_9738_),
    .C(_9739_),
    .Y(_9741_)
);

OAI21X1 _19802_ (
    .A(_9476_),
    .B(_9478_),
    .C(_9474_),
    .Y(_9742_)
);

NAND3X1 _19803_ (
    .A(_9742_),
    .B(_9741_),
    .C(_9736_),
    .Y(_9743_)
);

AOI21X1 _19804_ (
    .A(_9738_),
    .B(_9739_),
    .C(_9737_),
    .Y(_9744_)
);

AOI21X1 _19805_ (
    .A(_9735_),
    .B(_9728_),
    .C(_9687_),
    .Y(_9745_)
);

AOI21X1 _19806_ (
    .A(_9391_),
    .B(_9470_),
    .C(_9479_),
    .Y(_9746_)
);

OAI21X1 _19807_ (
    .A(_9745_),
    .B(_9744_),
    .C(_9746_),
    .Y(_9747_)
);

NAND3X1 _19808_ (
    .A(_9645_),
    .B(_9743_),
    .C(_9747_),
    .Y(_9748_)
);

AND2X2 _19809_ (
    .A(_9370_),
    .B(_9360_),
    .Y(_9749_)
);

NAND3X1 _19810_ (
    .A(_9741_),
    .B(_9746_),
    .C(_9736_),
    .Y(_9750_)
);

OAI21X1 _19811_ (
    .A(_9745_),
    .B(_9744_),
    .C(_9742_),
    .Y(_9752_)
);

NAND3X1 _19812_ (
    .A(_9750_),
    .B(_9752_),
    .C(_9749_),
    .Y(_9753_)
);

NAND2X1 _19813_ (
    .A(_9748_),
    .B(_9753_),
    .Y(_9754_)
);

AOI21X1 _19814_ (
    .A(_9574_),
    .B(_9573_),
    .C(_9482_),
    .Y(_9755_)
);

OAI21X1 _19815_ (
    .A(_9481_),
    .B(_9755_),
    .C(_9581_),
    .Y(_9756_)
);

NAND2X1 _19816_ (
    .A(_9465_),
    .B(_9471_),
    .Y(_9757_)
);

NAND2X1 _19817_ (
    .A(areg_14_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_9758_)
);

NAND2X1 _19818_ (
    .A(areg_16_bF$buf4),
    .B(breg_21_bF$buf4),
    .Y(_9759_)
);

NOR2X1 _19819_ (
    .A(_9702_),
    .B(_9759_),
    .Y(_9760_)
);

AND2X2 _19820_ (
    .A(_9702_),
    .B(_9759_),
    .Y(_9761_)
);

NOR2X1 _19821_ (
    .A(_9760_),
    .B(_9761_),
    .Y(_9763_)
);

XNOR2X1 _19822_ (
    .A(_9763_),
    .B(_9758_),
    .Y(_9764_)
);

OAI21X1 _19823_ (
    .A(_9410_),
    .B(_9401_),
    .C(_9405_),
    .Y(_9765_)
);

NAND2X1 _19824_ (
    .A(areg_17_bF$buf4),
    .B(breg_20_bF$buf0),
    .Y(_9766_)
);

INVX2 _19825_ (
    .A(_9766_),
    .Y(_9767_)
);

AND2X2 _19826_ (
    .A(areg_18_bF$buf4),
    .B(breg_19_bF$buf4),
    .Y(_9768_)
);

AND2X2 _19827_ (
    .A(breg_18_bF$buf4),
    .B(areg_19_bF$buf1),
    .Y(_9769_)
);

NAND2X1 _19828_ (
    .A(_9768_),
    .B(_9769_),
    .Y(_9770_)
);

OAI21X1 _19829_ (
    .A(_3529__bF$buf4),
    .B(_3402__bF$buf1),
    .C(_9408_),
    .Y(_9771_)
);

NAND3X1 _19830_ (
    .A(_9767_),
    .B(_9771_),
    .C(_9770_),
    .Y(_9772_)
);

NAND2X1 _19831_ (
    .A(breg_18_bF$buf3),
    .B(areg_19_bF$buf0),
    .Y(_9774_)
);

NOR2X1 _19832_ (
    .A(_9408_),
    .B(_9774_),
    .Y(_9775_)
);

NOR2X1 _19833_ (
    .A(_9768_),
    .B(_9769_),
    .Y(_9776_)
);

OAI21X1 _19834_ (
    .A(_9776_),
    .B(_9775_),
    .C(_9766_),
    .Y(_9777_)
);

NAND3X1 _19835_ (
    .A(_9772_),
    .B(_9765_),
    .C(_9777_),
    .Y(_9778_)
);

AOI21X1 _19836_ (
    .A(_9402_),
    .B(_9406_),
    .C(_9409_),
    .Y(_9779_)
);

NOR3X1 _19837_ (
    .A(_9766_),
    .B(_9775_),
    .C(_9776_),
    .Y(_9780_)
);

AOI21X1 _19838_ (
    .A(_9771_),
    .B(_9770_),
    .C(_9767_),
    .Y(_9781_)
);

OAI21X1 _19839_ (
    .A(_9780_),
    .B(_9781_),
    .C(_9779_),
    .Y(_9782_)
);

NAND3X1 _19840_ (
    .A(_9778_),
    .B(_9782_),
    .C(_9764_),
    .Y(_9783_)
);

INVX2 _19841_ (
    .A(_9758_),
    .Y(_9785_)
);

XNOR2X1 _19842_ (
    .A(_9763_),
    .B(_9785_),
    .Y(_9786_)
);

NOR3X1 _19843_ (
    .A(_9779_),
    .B(_9781_),
    .C(_9780_),
    .Y(_9787_)
);

AOI21X1 _19844_ (
    .A(_9772_),
    .B(_9777_),
    .C(_9765_),
    .Y(_9788_)
);

OAI21X1 _19845_ (
    .A(_9787_),
    .B(_9788_),
    .C(_9786_),
    .Y(_9789_)
);

NAND2X1 _19846_ (
    .A(_9783_),
    .B(_9789_),
    .Y(_9790_)
);

OAI21X1 _19847_ (
    .A(_9460_),
    .B(_9427_),
    .C(_9452_),
    .Y(_9791_)
);

AND2X2 _19848_ (
    .A(breg_16_bF$buf4),
    .B(areg_21_bF$buf0),
    .Y(_9792_)
);

AOI21X1 _19849_ (
    .A(_9045_),
    .B(_9792_),
    .C(_9443_),
    .Y(_9793_)
);

NAND2X1 _19850_ (
    .A(breg_17_bF$buf3),
    .B(areg_20_bF$buf2),
    .Y(_9794_)
);

INVX1 _19851_ (
    .A(_9794_),
    .Y(_9796_)
);

AND2X2 _19852_ (
    .A(breg_15_bF$buf5),
    .B(areg_22_bF$buf0),
    .Y(_9797_)
);

NAND2X1 _19853_ (
    .A(_9792_),
    .B(_9797_),
    .Y(_9798_)
);

OAI22X1 _19854_ (
    .A(_2362__bF$buf0),
    .B(_4551__bF$buf0),
    .C(_2560__bF$buf3),
    .D(_3961__bF$buf1),
    .Y(_9799_)
);

NAND3X1 _19855_ (
    .A(_9796_),
    .B(_9799_),
    .C(_9798_),
    .Y(_9800_)
);

OAI21X1 _19856_ (
    .A(_2560__bF$buf2),
    .B(_3961__bF$buf0),
    .C(_9797_),
    .Y(_9801_)
);

OAI21X1 _19857_ (
    .A(_2362__bF$buf5),
    .B(_4551__bF$buf4),
    .C(_9792_),
    .Y(_9802_)
);

NAND3X1 _19858_ (
    .A(_9794_),
    .B(_9801_),
    .C(_9802_),
    .Y(_9803_)
);

NOR2X1 _19859_ (
    .A(_9446_),
    .B(_9485_),
    .Y(_9804_)
);

OAI21X1 _19860_ (
    .A(_2586__bF$buf4),
    .B(_5921__bF$buf0),
    .C(_9446_),
    .Y(_9805_)
);

AOI21X1 _19861_ (
    .A(_9511_),
    .B(_9805_),
    .C(_9804_),
    .Y(_9807_)
);

NAND3X1 _19862_ (
    .A(_9807_),
    .B(_9800_),
    .C(_9803_),
    .Y(_9808_)
);

AOI21X1 _19863_ (
    .A(_9801_),
    .B(_9802_),
    .C(_9794_),
    .Y(_9809_)
);

AOI21X1 _19864_ (
    .A(_9799_),
    .B(_9798_),
    .C(_9796_),
    .Y(_9810_)
);

NAND2X1 _19865_ (
    .A(breg_13_bF$buf0),
    .B(areg_24_bF$buf1),
    .Y(_9811_)
);

AND2X2 _19866_ (
    .A(_9446_),
    .B(_9485_),
    .Y(_9812_)
);

OAI22X1 _19867_ (
    .A(_9100_),
    .B(_9811_),
    .C(_9812_),
    .D(_9484_),
    .Y(_9813_)
);

OAI21X1 _19868_ (
    .A(_9809_),
    .B(_9810_),
    .C(_9813_),
    .Y(_9814_)
);

AOI21X1 _19869_ (
    .A(_9808_),
    .B(_9814_),
    .C(_9793_),
    .Y(_9815_)
);

INVX1 _19870_ (
    .A(_9430_),
    .Y(_9816_)
);

OAI21X1 _19871_ (
    .A(_9432_),
    .B(_9816_),
    .C(_9435_),
    .Y(_9818_)
);

NAND3X1 _19872_ (
    .A(_9800_),
    .B(_9803_),
    .C(_9813_),
    .Y(_9819_)
);

OAI21X1 _19873_ (
    .A(_9809_),
    .B(_9810_),
    .C(_9807_),
    .Y(_9820_)
);

AOI21X1 _19874_ (
    .A(_9819_),
    .B(_9820_),
    .C(_9818_),
    .Y(_9821_)
);

OAI21X1 _19875_ (
    .A(_9815_),
    .B(_9821_),
    .C(_9791_),
    .Y(_9822_)
);

AOI21X1 _19876_ (
    .A(_9451_),
    .B(_9453_),
    .C(_9459_),
    .Y(_9823_)
);

NAND3X1 _19877_ (
    .A(_9818_),
    .B(_9819_),
    .C(_9820_),
    .Y(_9824_)
);

NOR3X1 _19878_ (
    .A(_9810_),
    .B(_9807_),
    .C(_9809_),
    .Y(_9825_)
);

AOI21X1 _19879_ (
    .A(_9800_),
    .B(_9803_),
    .C(_9813_),
    .Y(_9826_)
);

OAI21X1 _19880_ (
    .A(_9825_),
    .B(_9826_),
    .C(_9793_),
    .Y(_9827_)
);

NAND3X1 _19881_ (
    .A(_9823_),
    .B(_9824_),
    .C(_9827_),
    .Y(_9829_)
);

AOI21X1 _19882_ (
    .A(_9822_),
    .B(_9829_),
    .C(_9790_),
    .Y(_9830_)
);

OAI21X1 _19883_ (
    .A(_9780_),
    .B(_9781_),
    .C(_9765_),
    .Y(_9831_)
);

NAND3X1 _19884_ (
    .A(_9779_),
    .B(_9772_),
    .C(_9777_),
    .Y(_9832_)
);

AOI21X1 _19885_ (
    .A(_9831_),
    .B(_9832_),
    .C(_9786_),
    .Y(_9833_)
);

AOI21X1 _19886_ (
    .A(_9782_),
    .B(_9778_),
    .C(_9764_),
    .Y(_9834_)
);

NOR2X1 _19887_ (
    .A(_9833_),
    .B(_9834_),
    .Y(_9835_)
);

NAND3X1 _19888_ (
    .A(_9791_),
    .B(_9824_),
    .C(_9827_),
    .Y(_9836_)
);

OAI21X1 _19889_ (
    .A(_9815_),
    .B(_9821_),
    .C(_9823_),
    .Y(_9837_)
);

AOI21X1 _19890_ (
    .A(_9837_),
    .B(_9836_),
    .C(_9835_),
    .Y(_9838_)
);

NOR3X1 _19891_ (
    .A(_9519_),
    .B(_9520_),
    .C(_9518_),
    .Y(_9840_)
);

AOI21X1 _19892_ (
    .A(_9483_),
    .B(_9522_),
    .C(_9840_),
    .Y(_9841_)
);

OAI21X1 _19893_ (
    .A(_9838_),
    .B(_9830_),
    .C(_9841_),
    .Y(_9842_)
);

NAND3X1 _19894_ (
    .A(_9837_),
    .B(_9836_),
    .C(_9835_),
    .Y(_9843_)
);

NAND3X1 _19895_ (
    .A(_9822_),
    .B(_9790_),
    .C(_9829_),
    .Y(_9844_)
);

AOI21X1 _19896_ (
    .A(_9509_),
    .B(_9515_),
    .C(_9516_),
    .Y(_9845_)
);

OAI21X1 _19897_ (
    .A(_9524_),
    .B(_9845_),
    .C(_9517_),
    .Y(_9846_)
);

NAND3X1 _19898_ (
    .A(_9844_),
    .B(_9843_),
    .C(_9846_),
    .Y(_9847_)
);

NAND3X1 _19899_ (
    .A(_9757_),
    .B(_9847_),
    .C(_9842_),
    .Y(_9848_)
);

AND2X2 _19900_ (
    .A(_9471_),
    .B(_9465_),
    .Y(_9849_)
);

AOI21X1 _19901_ (
    .A(_9844_),
    .B(_9843_),
    .C(_9846_),
    .Y(_9851_)
);

NOR3X1 _19902_ (
    .A(_9830_),
    .B(_9838_),
    .C(_9841_),
    .Y(_9852_)
);

OAI21X1 _19903_ (
    .A(_9852_),
    .B(_9851_),
    .C(_9849_),
    .Y(_9853_)
);

NAND2X1 _19904_ (
    .A(_9848_),
    .B(_9853_),
    .Y(_9854_)
);

OAI21X1 _19905_ (
    .A(_9568_),
    .B(_9528_),
    .C(_9567_),
    .Y(_9855_)
);

AND2X2 _19906_ (
    .A(_9509_),
    .B(_9502_),
    .Y(_9856_)
);

NAND2X1 _19907_ (
    .A(breg_14_bF$buf2),
    .B(areg_23_bF$buf2),
    .Y(_9857_)
);

NAND2X1 _19908_ (
    .A(breg_12_bF$buf3),
    .B(areg_25_bF$buf3),
    .Y(_9858_)
);

XOR2X1 _19909_ (
    .A(_9811_),
    .B(_9858_),
    .Y(_9859_)
);

XNOR2X1 _19910_ (
    .A(_9859_),
    .B(_9857_),
    .Y(_9860_)
);

OAI21X1 _19911_ (
    .A(_9500_),
    .B(_9490_),
    .C(_9494_),
    .Y(_9862_)
);

NAND2X1 _19912_ (
    .A(breg_11_bF$buf0),
    .B(areg_26_bF$buf3),
    .Y(_9863_)
);

INVX2 _19913_ (
    .A(_9863_),
    .Y(_9864_)
);

AND2X2 _19914_ (
    .A(breg_10_bF$buf4),
    .B(areg_27_bF$buf1),
    .Y(_9865_)
);

AND2X2 _19915_ (
    .A(breg_9_bF$buf1),
    .B(areg_28_bF$buf2),
    .Y(_9866_)
);

NAND2X1 _19916_ (
    .A(_9865_),
    .B(_9866_),
    .Y(_9867_)
);

NAND2X1 _19917_ (
    .A(breg_10_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_9868_)
);

OAI21X1 _19918_ (
    .A(_6044__bF$buf3),
    .B(_7520__bF$buf2),
    .C(_9868_),
    .Y(_9869_)
);

NAND3X1 _19919_ (
    .A(_9864_),
    .B(_9869_),
    .C(_9867_),
    .Y(_9870_)
);

NAND2X1 _19920_ (
    .A(breg_9_bF$buf0),
    .B(areg_28_bF$buf1),
    .Y(_9871_)
);

NOR2X1 _19921_ (
    .A(_9868_),
    .B(_9871_),
    .Y(_9873_)
);

NOR2X1 _19922_ (
    .A(_9865_),
    .B(_9866_),
    .Y(_9874_)
);

OAI21X1 _19923_ (
    .A(_9874_),
    .B(_9873_),
    .C(_9863_),
    .Y(_9875_)
);

NAND3X1 _19924_ (
    .A(_9870_),
    .B(_9862_),
    .C(_9875_),
    .Y(_9876_)
);

AOI21X1 _19925_ (
    .A(_9491_),
    .B(_9495_),
    .C(_9498_),
    .Y(_9877_)
);

OAI21X1 _19926_ (
    .A(_7217__bF$buf2),
    .B(_7100__bF$buf0),
    .C(_9866_),
    .Y(_9878_)
);

OAI21X1 _19927_ (
    .A(_6044__bF$buf2),
    .B(_7520__bF$buf1),
    .C(_9865_),
    .Y(_9879_)
);

AOI21X1 _19928_ (
    .A(_9878_),
    .B(_9879_),
    .C(_9863_),
    .Y(_9880_)
);

AOI21X1 _19929_ (
    .A(_9869_),
    .B(_9867_),
    .C(_9864_),
    .Y(_9881_)
);

OAI21X1 _19930_ (
    .A(_9880_),
    .B(_9881_),
    .C(_9877_),
    .Y(_9882_)
);

NAND3X1 _19931_ (
    .A(_9876_),
    .B(_9882_),
    .C(_9860_),
    .Y(_9884_)
);

INVX2 _19932_ (
    .A(_9857_),
    .Y(_9885_)
);

XNOR2X1 _19933_ (
    .A(_9859_),
    .B(_9885_),
    .Y(_9886_)
);

OAI21X1 _19934_ (
    .A(_9880_),
    .B(_9881_),
    .C(_9862_),
    .Y(_9887_)
);

NAND3X1 _19935_ (
    .A(_9877_),
    .B(_9870_),
    .C(_9875_),
    .Y(_9888_)
);

NAND3X1 _19936_ (
    .A(_9887_),
    .B(_9888_),
    .C(_9886_),
    .Y(_9889_)
);

OAI21X1 _19937_ (
    .A(_9559_),
    .B(_9529_),
    .C(_9551_),
    .Y(_9890_)
);

NAND3X1 _19938_ (
    .A(_9890_),
    .B(_9884_),
    .C(_9889_),
    .Y(_9891_)
);

AOI21X1 _19939_ (
    .A(_9887_),
    .B(_9888_),
    .C(_9886_),
    .Y(_9892_)
);

AOI21X1 _19940_ (
    .A(_9876_),
    .B(_9882_),
    .C(_9860_),
    .Y(_9893_)
);

AOI21X1 _19941_ (
    .A(_9550_),
    .B(_9552_),
    .C(_9558_),
    .Y(_9894_)
);

OAI21X1 _19942_ (
    .A(_9892_),
    .B(_9893_),
    .C(_9894_),
    .Y(_9895_)
);

NAND3X1 _19943_ (
    .A(_9891_),
    .B(_9856_),
    .C(_9895_),
    .Y(_9896_)
);

NAND2X1 _19944_ (
    .A(_9502_),
    .B(_9509_),
    .Y(_9897_)
);

NAND3X1 _19945_ (
    .A(_9894_),
    .B(_9884_),
    .C(_9889_),
    .Y(_9898_)
);

OAI21X1 _19946_ (
    .A(_9892_),
    .B(_9893_),
    .C(_9890_),
    .Y(_9899_)
);

NAND3X1 _19947_ (
    .A(_9897_),
    .B(_9898_),
    .C(_9899_),
    .Y(_9900_)
);

NAND2X1 _19948_ (
    .A(breg_7_bF$buf5),
    .B(areg_30_bF$buf3),
    .Y(_9901_)
);

OAI21X1 _19949_ (
    .A(_9149_),
    .B(_9901_),
    .C(_9539_),
    .Y(_9902_)
);

NOR2X1 _19950_ (
    .A(_5420__bF$buf3),
    .B(_9153_),
    .Y(_9903_)
);

NAND2X1 _19951_ (
    .A(breg_6_bF$buf0),
    .B(areg_31_bF$buf4),
    .Y(_9905_)
);

NOR2X1 _19952_ (
    .A(_9905_),
    .B(_9535_),
    .Y(_9906_)
);

AOI21X1 _19953_ (
    .A(breg_6_bF$buf5),
    .B(areg_31_bF$buf3),
    .C(_9901_),
    .Y(_9907_)
);

OAI21X1 _19954_ (
    .A(_9906_),
    .B(_9907_),
    .C(_9903_),
    .Y(_9908_)
);

XNOR2X1 _19955_ (
    .A(_9901_),
    .B(_9905_),
    .Y(_9909_)
);

OAI21X1 _19956_ (
    .A(_5420__bF$buf2),
    .B(_9153_),
    .C(_9909_),
    .Y(_9910_)
);

NAND2X1 _19957_ (
    .A(_9908_),
    .B(_9910_),
    .Y(_9911_)
);

XNOR2X1 _19958_ (
    .A(_9911_),
    .B(_9902_),
    .Y(_9912_)
);

NAND2X1 _19959_ (
    .A(_9912_),
    .B(_9564_),
    .Y(_9913_)
);

XOR2X1 _19960_ (
    .A(_9911_),
    .B(_9902_),
    .Y(_9914_)
);

NAND2X1 _19961_ (
    .A(_9914_),
    .B(_9555_),
    .Y(_9916_)
);

AOI22X1 _19962_ (
    .A(_9913_),
    .B(_9916_),
    .C(_9896_),
    .D(_9900_),
    .Y(_9917_)
);

NAND3X1 _19963_ (
    .A(_9897_),
    .B(_9891_),
    .C(_9895_),
    .Y(_9918_)
);

NAND3X1 _19964_ (
    .A(_9898_),
    .B(_9856_),
    .C(_9899_),
    .Y(_9919_)
);

NAND2X1 _19965_ (
    .A(_9912_),
    .B(_9555_),
    .Y(_9920_)
);

NAND2X1 _19966_ (
    .A(_9914_),
    .B(_9564_),
    .Y(_9921_)
);

AOI22X1 _19967_ (
    .A(_9920_),
    .B(_9921_),
    .C(_9919_),
    .D(_9918_),
    .Y(_9922_)
);

OAI21X1 _19968_ (
    .A(_9917_),
    .B(_9922_),
    .C(_9855_),
    .Y(_9923_)
);

AND2X2 _19969_ (
    .A(_9527_),
    .B(_9523_),
    .Y(_9924_)
);

INVX1 _19970_ (
    .A(_9567_),
    .Y(_9925_)
);

AOI21X1 _19971_ (
    .A(_9562_),
    .B(_9924_),
    .C(_9925_),
    .Y(_9927_)
);

NOR2X1 _19972_ (
    .A(_9922_),
    .B(_9917_),
    .Y(_9928_)
);

NAND2X1 _19973_ (
    .A(_9928_),
    .B(_9927_),
    .Y(_9929_)
);

AOI21X1 _19974_ (
    .A(_9923_),
    .B(_9929_),
    .C(_9854_),
    .Y(_9930_)
);

OAI21X1 _19975_ (
    .A(_9852_),
    .B(_9851_),
    .C(_9757_),
    .Y(_9931_)
);

NAND3X1 _19976_ (
    .A(_9842_),
    .B(_9847_),
    .C(_9849_),
    .Y(_9932_)
);

NAND2X1 _19977_ (
    .A(_9932_),
    .B(_9931_),
    .Y(_9933_)
);

OAI21X1 _19978_ (
    .A(_9569_),
    .B(_9925_),
    .C(_9928_),
    .Y(_9934_)
);

OAI21X1 _19979_ (
    .A(_9917_),
    .B(_9922_),
    .C(_9927_),
    .Y(_9935_)
);

AOI21X1 _19980_ (
    .A(_9934_),
    .B(_9935_),
    .C(_9933_),
    .Y(_9936_)
);

OAI21X1 _19981_ (
    .A(_9930_),
    .B(_9936_),
    .C(_9756_),
    .Y(_9938_)
);

NOR3X1 _19982_ (
    .A(_9570_),
    .B(_9569_),
    .C(_9572_),
    .Y(_9939_)
);

AOI21X1 _19983_ (
    .A(_9582_),
    .B(_9580_),
    .C(_9939_),
    .Y(_9940_)
);

NAND3X1 _19984_ (
    .A(_9934_),
    .B(_9935_),
    .C(_9933_),
    .Y(_9941_)
);

AND2X2 _19985_ (
    .A(_9928_),
    .B(_9855_),
    .Y(_9942_)
);

NOR2X1 _19986_ (
    .A(_9855_),
    .B(_9928_),
    .Y(_9943_)
);

OAI21X1 _19987_ (
    .A(_9942_),
    .B(_9943_),
    .C(_9854_),
    .Y(_9944_)
);

NAND3X1 _19988_ (
    .A(_9941_),
    .B(_9944_),
    .C(_9940_),
    .Y(_9945_)
);

AOI21X1 _19989_ (
    .A(_9938_),
    .B(_9945_),
    .C(_9754_),
    .Y(_9946_)
);

NAND3X1 _19990_ (
    .A(_9743_),
    .B(_9747_),
    .C(_9749_),
    .Y(_9947_)
);

NAND3X1 _19991_ (
    .A(_9645_),
    .B(_9750_),
    .C(_9752_),
    .Y(_9949_)
);

NAND2X1 _19992_ (
    .A(_9949_),
    .B(_9947_),
    .Y(_9950_)
);

NAND3X1 _19993_ (
    .A(_9941_),
    .B(_9944_),
    .C(_9756_),
    .Y(_9951_)
);

OAI21X1 _19994_ (
    .A(_9930_),
    .B(_9936_),
    .C(_9940_),
    .Y(_9952_)
);

AOI21X1 _19995_ (
    .A(_9952_),
    .B(_9951_),
    .C(_9950_),
    .Y(_9953_)
);

OAI21X1 _19996_ (
    .A(_9946_),
    .B(_9953_),
    .C(_9644_),
    .Y(_9954_)
);

NOR3X1 _19997_ (
    .A(_9577_),
    .B(_9583_),
    .C(_9586_),
    .Y(_9955_)
);

AOI21X1 _19998_ (
    .A(_9594_),
    .B(_9596_),
    .C(_9955_),
    .Y(_9956_)
);

NAND3X1 _19999_ (
    .A(_9952_),
    .B(_9951_),
    .C(_9950_),
    .Y(_9957_)
);

NAND3X1 _20000_ (
    .A(_9938_),
    .B(_9945_),
    .C(_9754_),
    .Y(_9958_)
);

NAND3X1 _20001_ (
    .A(_9957_),
    .B(_9958_),
    .C(_9956_),
    .Y(_9960_)
);

AOI21X1 _20002_ (
    .A(_9954_),
    .B(_9960_),
    .C(_9642_),
    .Y(_9961_)
);

NAND3X1 _20003_ (
    .A(_9957_),
    .B(_9958_),
    .C(_9644_),
    .Y(_9962_)
);

OAI21X1 _20004_ (
    .A(_9946_),
    .B(_9953_),
    .C(_9956_),
    .Y(_9963_)
);

AOI21X1 _20005_ (
    .A(_9962_),
    .B(_9963_),
    .C(_9640_),
    .Y(_9964_)
);

OAI21X1 _20006_ (
    .A(_9961_),
    .B(_9964_),
    .C(_9639_),
    .Y(_9965_)
);

AOI21X1 _20007_ (
    .A(_9273_),
    .B(_9607_),
    .C(_9614_),
    .Y(_9966_)
);

NAND3X1 _20008_ (
    .A(_9640_),
    .B(_9962_),
    .C(_9963_),
    .Y(_9967_)
);

NAND3X1 _20009_ (
    .A(_9642_),
    .B(_9954_),
    .C(_9960_),
    .Y(_9968_)
);

NAND3X1 _20010_ (
    .A(_9967_),
    .B(_9968_),
    .C(_9966_),
    .Y(_9969_)
);

AOI21X1 _20011_ (
    .A(_9965_),
    .B(_9969_),
    .C(_9638_),
    .Y(_9971_)
);

NAND3X1 _20012_ (
    .A(_9967_),
    .B(_9968_),
    .C(_9639_),
    .Y(_9972_)
);

OAI21X1 _20013_ (
    .A(_9961_),
    .B(_9964_),
    .C(_9966_),
    .Y(_9973_)
);

AOI21X1 _20014_ (
    .A(_9972_),
    .B(_9973_),
    .C(_9637_),
    .Y(_9974_)
);

OAI21X1 _20015_ (
    .A(_9971_),
    .B(_9974_),
    .C(_9636_),
    .Y(_9975_)
);

NOR3X1 _20016_ (
    .A(_9605_),
    .B(_9608_),
    .C(_9612_),
    .Y(_9976_)
);

AOI21X1 _20017_ (
    .A(_9269_),
    .B(_9621_),
    .C(_9976_),
    .Y(_9977_)
);

NAND3X1 _20018_ (
    .A(_9637_),
    .B(_9972_),
    .C(_9973_),
    .Y(_9978_)
);

NAND3X1 _20019_ (
    .A(_9638_),
    .B(_9965_),
    .C(_9969_),
    .Y(_9979_)
);

NAND3X1 _20020_ (
    .A(_9978_),
    .B(_9979_),
    .C(_9977_),
    .Y(_9980_)
);

NAND2X1 _20021_ (
    .A(_9975_),
    .B(_9980_),
    .Y(_9982_)
);

XOR2X1 _20022_ (
    .A(_9634_),
    .B(_9982_),
    .Y(_0_[37])
);

NOR3X1 _20023_ (
    .A(_9618_),
    .B(_9622_),
    .C(_9625_),
    .Y(_9983_)
);

NOR3X1 _20024_ (
    .A(_9971_),
    .B(_9974_),
    .C(_9977_),
    .Y(_9984_)
);

OAI21X1 _20025_ (
    .A(_9971_),
    .B(_9974_),
    .C(_9977_),
    .Y(_9985_)
);

OAI21X1 _20026_ (
    .A(_9983_),
    .B(_9984_),
    .C(_9985_),
    .Y(_9986_)
);

AOI22X1 _20027_ (
    .A(_9975_),
    .B(_9980_),
    .C(_9623_),
    .D(_9628_),
    .Y(_9987_)
);

INVX1 _20028_ (
    .A(_9987_),
    .Y(_9988_)
);

OAI21X1 _20029_ (
    .A(_9632_),
    .B(_9988_),
    .C(_9986_),
    .Y(_9989_)
);

NOR3X1 _20030_ (
    .A(_9961_),
    .B(_9964_),
    .C(_9966_),
    .Y(_9990_)
);

AOI21X1 _20031_ (
    .A(_9637_),
    .B(_9973_),
    .C(_9990_),
    .Y(_9992_)
);

OAI21X1 _20032_ (
    .A(_9677_),
    .B(_9647_),
    .C(_9684_),
    .Y(_9993_)
);

AOI21X1 _20033_ (
    .A(_9957_),
    .B(_9958_),
    .C(_9644_),
    .Y(_9994_)
);

OAI21X1 _20034_ (
    .A(_9994_),
    .B(_9642_),
    .C(_9962_),
    .Y(_9995_)
);

NAND2X1 _20035_ (
    .A(_9743_),
    .B(_9748_),
    .Y(_9996_)
);

AOI21X1 _20036_ (
    .A(_9941_),
    .B(_9944_),
    .C(_9756_),
    .Y(_9997_)
);

OAI21X1 _20037_ (
    .A(_9754_),
    .B(_9997_),
    .C(_9951_),
    .Y(_9998_)
);

AND2X2 _20038_ (
    .A(_9736_),
    .B(_9728_),
    .Y(_9999_)
);

NOR2X1 _20039_ (
    .A(_4434__bF$buf1),
    .B(_7225__bF$buf2),
    .Y(_10000_)
);

INVX1 _20040_ (
    .A(_10000_),
    .Y(_10001_)
);

OAI21X1 _20041_ (
    .A(_9665_),
    .B(_9650_),
    .C(_9675_),
    .Y(_10003_)
);

NOR2X1 _20042_ (
    .A(_5190__bF$buf1),
    .B(_6815__bF$buf1),
    .Y(_10004_)
);

INVX2 _20043_ (
    .A(_10004_),
    .Y(_10005_)
);

OAI21X1 _20044_ (
    .A(_9662_),
    .B(_9653_),
    .C(_9657_),
    .Y(_10006_)
);

NAND2X1 _20045_ (
    .A(areg_9_bF$buf4),
    .B(breg_29_bF$buf0),
    .Y(_10007_)
);

INVX2 _20046_ (
    .A(_10007_),
    .Y(_10008_)
);

AND2X2 _20047_ (
    .A(areg_10_bF$buf3),
    .B(breg_28_bF$buf2),
    .Y(_10009_)
);

AND2X2 _20048_ (
    .A(areg_11_bF$buf4),
    .B(breg_27_bF$buf3),
    .Y(_10010_)
);

NAND2X1 _20049_ (
    .A(_10009_),
    .B(_10010_),
    .Y(_10011_)
);

OAI21X1 _20050_ (
    .A(_9104__bF$buf1),
    .B(_5668__bF$buf1),
    .C(_9660_),
    .Y(_10012_)
);

NAND3X1 _20051_ (
    .A(_10008_),
    .B(_10012_),
    .C(_10011_),
    .Y(_10014_)
);

NAND2X1 _20052_ (
    .A(areg_11_bF$buf3),
    .B(breg_27_bF$buf2),
    .Y(_10015_)
);

NOR2X1 _20053_ (
    .A(_9660_),
    .B(_10015_),
    .Y(_10016_)
);

NOR2X1 _20054_ (
    .A(_10009_),
    .B(_10010_),
    .Y(_10017_)
);

OAI21X1 _20055_ (
    .A(_10017_),
    .B(_10016_),
    .C(_10007_),
    .Y(_10018_)
);

AOI21X1 _20056_ (
    .A(_10014_),
    .B(_10018_),
    .C(_10006_),
    .Y(_10019_)
);

AOI21X1 _20057_ (
    .A(_9654_),
    .B(_9658_),
    .C(_9661_),
    .Y(_10020_)
);

OAI21X1 _20058_ (
    .A(_7711__bF$buf1),
    .B(_6050__bF$buf0),
    .C(_10010_),
    .Y(_10021_)
);

OAI21X1 _20059_ (
    .A(_9104__bF$buf0),
    .B(_5668__bF$buf0),
    .C(_10009_),
    .Y(_10022_)
);

AOI21X1 _20060_ (
    .A(_10021_),
    .B(_10022_),
    .C(_10007_),
    .Y(_10023_)
);

AOI21X1 _20061_ (
    .A(_10012_),
    .B(_10011_),
    .C(_10008_),
    .Y(_10025_)
);

NOR3X1 _20062_ (
    .A(_10025_),
    .B(_10020_),
    .C(_10023_),
    .Y(_10026_)
);

OAI21X1 _20063_ (
    .A(_10026_),
    .B(_10019_),
    .C(_10005_),
    .Y(_10027_)
);

OAI21X1 _20064_ (
    .A(_10023_),
    .B(_10025_),
    .C(_10020_),
    .Y(_10028_)
);

NAND3X1 _20065_ (
    .A(_10014_),
    .B(_10006_),
    .C(_10018_),
    .Y(_10029_)
);

NAND3X1 _20066_ (
    .A(_10004_),
    .B(_10028_),
    .C(_10029_),
    .Y(_10030_)
);

AOI21X1 _20067_ (
    .A(_10030_),
    .B(_10027_),
    .C(_10003_),
    .Y(_10031_)
);

AOI21X1 _20068_ (
    .A(_9649_),
    .B(_9673_),
    .C(_9671_),
    .Y(_10032_)
);

AOI21X1 _20069_ (
    .A(_10028_),
    .B(_10029_),
    .C(_10004_),
    .Y(_10033_)
);

NOR3X1 _20070_ (
    .A(_10019_),
    .B(_10005_),
    .C(_10026_),
    .Y(_10034_)
);

NOR3X1 _20071_ (
    .A(_10032_),
    .B(_10033_),
    .C(_10034_),
    .Y(_10036_)
);

OAI21X1 _20072_ (
    .A(_10036_),
    .B(_10031_),
    .C(_10001_),
    .Y(_10037_)
);

OAI21X1 _20073_ (
    .A(_10034_),
    .B(_10033_),
    .C(_10032_),
    .Y(_10038_)
);

NAND3X1 _20074_ (
    .A(_10003_),
    .B(_10030_),
    .C(_10027_),
    .Y(_10039_)
);

NAND3X1 _20075_ (
    .A(_10000_),
    .B(_10039_),
    .C(_10038_),
    .Y(_10040_)
);

AND2X2 _20076_ (
    .A(_10037_),
    .B(_10040_),
    .Y(_10041_)
);

OAI21X1 _20077_ (
    .A(_9726_),
    .B(_9724_),
    .C(_9717_),
    .Y(_10042_)
);

NAND2X1 _20078_ (
    .A(_9704_),
    .B(_9711_),
    .Y(_10043_)
);

OAI21X1 _20079_ (
    .A(_9695_),
    .B(_9691_),
    .C(_9699_),
    .Y(_10044_)
);

NAND2X1 _20080_ (
    .A(areg_12_bF$buf0),
    .B(breg_26_bF$buf2),
    .Y(_10045_)
);

NAND2X1 _20081_ (
    .A(areg_13_bF$buf3),
    .B(breg_25_bF$buf5),
    .Y(_10047_)
);

NAND2X1 _20082_ (
    .A(areg_14_bF$buf2),
    .B(breg_24_bF$buf0),
    .Y(_10048_)
);

NOR2X1 _20083_ (
    .A(_10047_),
    .B(_10048_),
    .Y(_10049_)
);

AND2X2 _20084_ (
    .A(_10047_),
    .B(_10048_),
    .Y(_10050_)
);

OAI21X1 _20085_ (
    .A(_10050_),
    .B(_10049_),
    .C(_10045_),
    .Y(_10051_)
);

INVX1 _20086_ (
    .A(_10045_),
    .Y(_10052_)
);

OR2X2 _20087_ (
    .A(_10047_),
    .B(_10048_),
    .Y(_10053_)
);

OAI21X1 _20088_ (
    .A(_2287__bF$buf3),
    .B(_5315__bF$buf0),
    .C(_10047_),
    .Y(_10054_)
);

NAND3X1 _20089_ (
    .A(_10052_),
    .B(_10054_),
    .C(_10053_),
    .Y(_10055_)
);

NAND2X1 _20090_ (
    .A(areg_16_bF$buf3),
    .B(breg_22_bF$buf3),
    .Y(_10056_)
);

OAI22X1 _20091_ (
    .A(_9394_),
    .B(_10056_),
    .C(_9761_),
    .D(_9758_),
    .Y(_10058_)
);

NAND3X1 _20092_ (
    .A(_10051_),
    .B(_10055_),
    .C(_10058_),
    .Y(_10059_)
);

AOI21X1 _20093_ (
    .A(_10054_),
    .B(_10053_),
    .C(_10052_),
    .Y(_10060_)
);

NOR3X1 _20094_ (
    .A(_10045_),
    .B(_10049_),
    .C(_10050_),
    .Y(_10061_)
);

OAI21X1 _20095_ (
    .A(_2669__bF$buf1),
    .B(_3781__bF$buf1),
    .C(_9702_),
    .Y(_10062_)
);

AOI21X1 _20096_ (
    .A(_9785_),
    .B(_10062_),
    .C(_9760_),
    .Y(_10063_)
);

OAI21X1 _20097_ (
    .A(_10061_),
    .B(_10060_),
    .C(_10063_),
    .Y(_10064_)
);

NAND3X1 _20098_ (
    .A(_10044_),
    .B(_10059_),
    .C(_10064_),
    .Y(_10065_)
);

INVX1 _20099_ (
    .A(_10044_),
    .Y(_10066_)
);

NAND3X1 _20100_ (
    .A(_10063_),
    .B(_10051_),
    .C(_10055_),
    .Y(_10067_)
);

OAI21X1 _20101_ (
    .A(_10061_),
    .B(_10060_),
    .C(_10058_),
    .Y(_10069_)
);

NAND3X1 _20102_ (
    .A(_10066_),
    .B(_10067_),
    .C(_10069_),
    .Y(_10070_)
);

OAI21X1 _20103_ (
    .A(_9786_),
    .B(_9788_),
    .C(_9778_),
    .Y(_10071_)
);

NAND3X1 _20104_ (
    .A(_10065_),
    .B(_10070_),
    .C(_10071_),
    .Y(_10072_)
);

AOI21X1 _20105_ (
    .A(_10067_),
    .B(_10069_),
    .C(_10066_),
    .Y(_10073_)
);

AOI21X1 _20106_ (
    .A(_10059_),
    .B(_10064_),
    .C(_10044_),
    .Y(_10074_)
);

AOI21X1 _20107_ (
    .A(_9782_),
    .B(_9764_),
    .C(_9787_),
    .Y(_10075_)
);

OAI21X1 _20108_ (
    .A(_10073_),
    .B(_10074_),
    .C(_10075_),
    .Y(_10076_)
);

NAND3X1 _20109_ (
    .A(_10043_),
    .B(_10076_),
    .C(_10072_),
    .Y(_10077_)
);

AND2X2 _20110_ (
    .A(_9711_),
    .B(_9704_),
    .Y(_10078_)
);

NOR3X1 _20111_ (
    .A(_10073_),
    .B(_10074_),
    .C(_10075_),
    .Y(_10080_)
);

AOI21X1 _20112_ (
    .A(_10065_),
    .B(_10070_),
    .C(_10071_),
    .Y(_10081_)
);

OAI21X1 _20113_ (
    .A(_10080_),
    .B(_10081_),
    .C(_10078_),
    .Y(_10082_)
);

NAND3X1 _20114_ (
    .A(_10077_),
    .B(_10042_),
    .C(_10082_),
    .Y(_10083_)
);

AOI21X1 _20115_ (
    .A(_9689_),
    .B(_9722_),
    .C(_9725_),
    .Y(_10084_)
);

NAND3X1 _20116_ (
    .A(_10065_),
    .B(_10070_),
    .C(_10075_),
    .Y(_10085_)
);

OAI21X1 _20117_ (
    .A(_10073_),
    .B(_10074_),
    .C(_10071_),
    .Y(_10086_)
);

AOI21X1 _20118_ (
    .A(_10086_),
    .B(_10085_),
    .C(_10078_),
    .Y(_10087_)
);

AOI21X1 _20119_ (
    .A(_10076_),
    .B(_10072_),
    .C(_10043_),
    .Y(_10088_)
);

OAI21X1 _20120_ (
    .A(_10087_),
    .B(_10088_),
    .C(_10084_),
    .Y(_10089_)
);

NAND3X1 _20121_ (
    .A(_10089_),
    .B(_10083_),
    .C(_10041_),
    .Y(_10091_)
);

NAND2X1 _20122_ (
    .A(_10040_),
    .B(_10037_),
    .Y(_10092_)
);

OAI21X1 _20123_ (
    .A(_10087_),
    .B(_10088_),
    .C(_10042_),
    .Y(_10093_)
);

NAND3X1 _20124_ (
    .A(_10084_),
    .B(_10077_),
    .C(_10082_),
    .Y(_10094_)
);

NAND3X1 _20125_ (
    .A(_10092_),
    .B(_10093_),
    .C(_10094_),
    .Y(_10095_)
);

OAI21X1 _20126_ (
    .A(_9849_),
    .B(_9851_),
    .C(_9847_),
    .Y(_10096_)
);

NAND3X1 _20127_ (
    .A(_10096_),
    .B(_10095_),
    .C(_10091_),
    .Y(_10097_)
);

AOI21X1 _20128_ (
    .A(_10093_),
    .B(_10094_),
    .C(_10092_),
    .Y(_10098_)
);

AOI21X1 _20129_ (
    .A(_10089_),
    .B(_10083_),
    .C(_10041_),
    .Y(_10099_)
);

AOI21X1 _20130_ (
    .A(_9757_),
    .B(_9842_),
    .C(_9852_),
    .Y(_10100_)
);

OAI21X1 _20131_ (
    .A(_10099_),
    .B(_10098_),
    .C(_10100_),
    .Y(_10102_)
);

NAND3X1 _20132_ (
    .A(_10097_),
    .B(_9999_),
    .C(_10102_),
    .Y(_10103_)
);

NAND2X1 _20133_ (
    .A(_9728_),
    .B(_9736_),
    .Y(_10104_)
);

NAND3X1 _20134_ (
    .A(_10100_),
    .B(_10095_),
    .C(_10091_),
    .Y(_10105_)
);

OAI21X1 _20135_ (
    .A(_10099_),
    .B(_10098_),
    .C(_10096_),
    .Y(_10106_)
);

NAND3X1 _20136_ (
    .A(_10104_),
    .B(_10105_),
    .C(_10106_),
    .Y(_10107_)
);

NAND2X1 _20137_ (
    .A(_10107_),
    .B(_10103_),
    .Y(_10108_)
);

OAI21X1 _20138_ (
    .A(_9854_),
    .B(_9943_),
    .C(_9934_),
    .Y(_10109_)
);

NAND2X1 _20139_ (
    .A(_9836_),
    .B(_9843_),
    .Y(_10110_)
);

NAND2X1 _20140_ (
    .A(areg_15_bF$buf0),
    .B(breg_23_bF$buf0),
    .Y(_10111_)
);

INVX2 _20141_ (
    .A(_10111_),
    .Y(_10113_)
);

NAND2X1 _20142_ (
    .A(areg_17_bF$buf3),
    .B(breg_21_bF$buf3),
    .Y(_10114_)
);

XOR2X1 _20143_ (
    .A(_10056_),
    .B(_10114_),
    .Y(_10115_)
);

XNOR2X1 _20144_ (
    .A(_10115_),
    .B(_10113_),
    .Y(_10116_)
);

OAI21X1 _20145_ (
    .A(_9776_),
    .B(_9766_),
    .C(_9770_),
    .Y(_10117_)
);

NAND2X1 _20146_ (
    .A(areg_18_bF$buf3),
    .B(breg_20_bF$buf4),
    .Y(_10118_)
);

NAND2X1 _20147_ (
    .A(breg_19_bF$buf3),
    .B(areg_20_bF$buf1),
    .Y(_10119_)
);

NOR2X1 _20148_ (
    .A(_9774_),
    .B(_10119_),
    .Y(_10120_)
);

AND2X2 _20149_ (
    .A(areg_19_bF$buf5),
    .B(breg_19_bF$buf2),
    .Y(_10121_)
);

AND2X2 _20150_ (
    .A(breg_18_bF$buf2),
    .B(areg_20_bF$buf0),
    .Y(_10122_)
);

NOR2X1 _20151_ (
    .A(_10121_),
    .B(_10122_),
    .Y(_10124_)
);

NOR3X1 _20152_ (
    .A(_10118_),
    .B(_10120_),
    .C(_10124_),
    .Y(_10125_)
);

INVX2 _20153_ (
    .A(_10118_),
    .Y(_10126_)
);

NAND2X1 _20154_ (
    .A(_10121_),
    .B(_10122_),
    .Y(_10127_)
);

OAI22X1 _20155_ (
    .A(_3529__bF$buf3),
    .B(_3958__bF$buf3),
    .C(_3402__bF$buf0),
    .D(_3253__bF$buf0),
    .Y(_10128_)
);

AOI21X1 _20156_ (
    .A(_10128_),
    .B(_10127_),
    .C(_10126_),
    .Y(_10129_)
);

OAI21X1 _20157_ (
    .A(_10125_),
    .B(_10129_),
    .C(_10117_),
    .Y(_10130_)
);

AOI21X1 _20158_ (
    .A(_9767_),
    .B(_9771_),
    .C(_9775_),
    .Y(_10131_)
);

NAND3X1 _20159_ (
    .A(_10126_),
    .B(_10128_),
    .C(_10127_),
    .Y(_10132_)
);

OAI21X1 _20160_ (
    .A(_10124_),
    .B(_10120_),
    .C(_10118_),
    .Y(_10133_)
);

NAND3X1 _20161_ (
    .A(_10131_),
    .B(_10132_),
    .C(_10133_),
    .Y(_10135_)
);

AOI21X1 _20162_ (
    .A(_10135_),
    .B(_10130_),
    .C(_10116_),
    .Y(_10136_)
);

XNOR2X1 _20163_ (
    .A(_10115_),
    .B(_10111_),
    .Y(_10137_)
);

NAND3X1 _20164_ (
    .A(_10132_),
    .B(_10117_),
    .C(_10133_),
    .Y(_10138_)
);

OAI21X1 _20165_ (
    .A(_10125_),
    .B(_10129_),
    .C(_10131_),
    .Y(_10139_)
);

AOI21X1 _20166_ (
    .A(_10138_),
    .B(_10139_),
    .C(_10137_),
    .Y(_10140_)
);

NOR2X1 _20167_ (
    .A(_10136_),
    .B(_10140_),
    .Y(_10141_)
);

OAI21X1 _20168_ (
    .A(_9826_),
    .B(_9793_),
    .C(_9819_),
    .Y(_10142_)
);

NAND2X1 _20169_ (
    .A(breg_16_bF$buf3),
    .B(areg_22_bF$buf4),
    .Y(_10143_)
);

OAI21X1 _20170_ (
    .A(_9816_),
    .B(_10143_),
    .C(_9800_),
    .Y(_10144_)
);

NAND2X1 _20171_ (
    .A(breg_17_bF$buf2),
    .B(areg_21_bF$buf4),
    .Y(_10146_)
);

INVX1 _20172_ (
    .A(_10146_),
    .Y(_10147_)
);

AND2X2 _20173_ (
    .A(breg_16_bF$buf2),
    .B(areg_22_bF$buf3),
    .Y(_10148_)
);

AND2X2 _20174_ (
    .A(breg_15_bF$buf4),
    .B(areg_23_bF$buf1),
    .Y(_10149_)
);

NAND2X1 _20175_ (
    .A(_10148_),
    .B(_10149_),
    .Y(_10150_)
);

OAI21X1 _20176_ (
    .A(_2362__bF$buf4),
    .B(_4541__bF$buf2),
    .C(_10143_),
    .Y(_10151_)
);

NAND3X1 _20177_ (
    .A(_10147_),
    .B(_10151_),
    .C(_10150_),
    .Y(_10152_)
);

OAI21X1 _20178_ (
    .A(_2560__bF$buf1),
    .B(_4551__bF$buf3),
    .C(_10149_),
    .Y(_10153_)
);

OAI21X1 _20179_ (
    .A(_2362__bF$buf3),
    .B(_4541__bF$buf1),
    .C(_10148_),
    .Y(_10154_)
);

NAND3X1 _20180_ (
    .A(_10146_),
    .B(_10153_),
    .C(_10154_),
    .Y(_10155_)
);

NAND2X1 _20181_ (
    .A(breg_13_bF$buf4),
    .B(areg_25_bF$buf2),
    .Y(_10157_)
);

AND2X2 _20182_ (
    .A(_9811_),
    .B(_9858_),
    .Y(_10158_)
);

OAI22X1 _20183_ (
    .A(_9485_),
    .B(_10157_),
    .C(_10158_),
    .D(_9857_),
    .Y(_10159_)
);

NAND3X1 _20184_ (
    .A(_10152_),
    .B(_10155_),
    .C(_10159_),
    .Y(_10160_)
);

AOI21X1 _20185_ (
    .A(_10153_),
    .B(_10154_),
    .C(_10146_),
    .Y(_10161_)
);

AOI21X1 _20186_ (
    .A(_10151_),
    .B(_10150_),
    .C(_10147_),
    .Y(_10162_)
);

NOR2X1 _20187_ (
    .A(_9811_),
    .B(_9858_),
    .Y(_10163_)
);

OAI21X1 _20188_ (
    .A(_2586__bF$buf3),
    .B(_6300__bF$buf3),
    .C(_9811_),
    .Y(_10164_)
);

AOI21X1 _20189_ (
    .A(_9885_),
    .B(_10164_),
    .C(_10163_),
    .Y(_10165_)
);

OAI21X1 _20190_ (
    .A(_10161_),
    .B(_10162_),
    .C(_10165_),
    .Y(_10166_)
);

NAND3X1 _20191_ (
    .A(_10144_),
    .B(_10160_),
    .C(_10166_),
    .Y(_10168_)
);

AOI21X1 _20192_ (
    .A(_9430_),
    .B(_10148_),
    .C(_9809_),
    .Y(_10169_)
);

NOR3X1 _20193_ (
    .A(_10162_),
    .B(_10165_),
    .C(_10161_),
    .Y(_10170_)
);

AOI21X1 _20194_ (
    .A(_10152_),
    .B(_10155_),
    .C(_10159_),
    .Y(_10171_)
);

OAI21X1 _20195_ (
    .A(_10170_),
    .B(_10171_),
    .C(_10169_),
    .Y(_10172_)
);

NAND3X1 _20196_ (
    .A(_10142_),
    .B(_10168_),
    .C(_10172_),
    .Y(_10173_)
);

AOI21X1 _20197_ (
    .A(_9818_),
    .B(_9820_),
    .C(_9825_),
    .Y(_10174_)
);

NAND3X1 _20198_ (
    .A(_10165_),
    .B(_10152_),
    .C(_10155_),
    .Y(_10175_)
);

OAI21X1 _20199_ (
    .A(_10161_),
    .B(_10162_),
    .C(_10159_),
    .Y(_10176_)
);

AOI21X1 _20200_ (
    .A(_10175_),
    .B(_10176_),
    .C(_10169_),
    .Y(_10177_)
);

AOI21X1 _20201_ (
    .A(_10160_),
    .B(_10166_),
    .C(_10144_),
    .Y(_10179_)
);

OAI21X1 _20202_ (
    .A(_10177_),
    .B(_10179_),
    .C(_10174_),
    .Y(_10180_)
);

NAND3X1 _20203_ (
    .A(_10180_),
    .B(_10141_),
    .C(_10173_),
    .Y(_10181_)
);

NAND3X1 _20204_ (
    .A(_10138_),
    .B(_10139_),
    .C(_10137_),
    .Y(_10182_)
);

NOR3X1 _20205_ (
    .A(_10131_),
    .B(_10129_),
    .C(_10125_),
    .Y(_10183_)
);

AOI21X1 _20206_ (
    .A(_10132_),
    .B(_10133_),
    .C(_10117_),
    .Y(_10184_)
);

OAI21X1 _20207_ (
    .A(_10183_),
    .B(_10184_),
    .C(_10116_),
    .Y(_10185_)
);

NAND2X1 _20208_ (
    .A(_10182_),
    .B(_10185_),
    .Y(_10186_)
);

OAI21X1 _20209_ (
    .A(_10177_),
    .B(_10179_),
    .C(_10142_),
    .Y(_10187_)
);

NAND3X1 _20210_ (
    .A(_10174_),
    .B(_10168_),
    .C(_10172_),
    .Y(_10188_)
);

NAND3X1 _20211_ (
    .A(_10187_),
    .B(_10186_),
    .C(_10188_),
    .Y(_10190_)
);

AOI21X1 _20212_ (
    .A(_9884_),
    .B(_9889_),
    .C(_9890_),
    .Y(_10191_)
);

OAI21X1 _20213_ (
    .A(_10191_),
    .B(_9856_),
    .C(_9891_),
    .Y(_10192_)
);

AOI21X1 _20214_ (
    .A(_10190_),
    .B(_10181_),
    .C(_10192_),
    .Y(_10193_)
);

AOI21X1 _20215_ (
    .A(_10187_),
    .B(_10188_),
    .C(_10186_),
    .Y(_10194_)
);

AOI21X1 _20216_ (
    .A(_10180_),
    .B(_10173_),
    .C(_10141_),
    .Y(_10195_)
);

NOR3X1 _20217_ (
    .A(_9893_),
    .B(_9894_),
    .C(_9892_),
    .Y(_10196_)
);

AOI21X1 _20218_ (
    .A(_9897_),
    .B(_9895_),
    .C(_10196_),
    .Y(_10197_)
);

NOR3X1 _20219_ (
    .A(_10194_),
    .B(_10195_),
    .C(_10197_),
    .Y(_10198_)
);

OAI21X1 _20220_ (
    .A(_10198_),
    .B(_10193_),
    .C(_10110_),
    .Y(_10199_)
);

AND2X2 _20221_ (
    .A(_9843_),
    .B(_9836_),
    .Y(_10201_)
);

OAI21X1 _20222_ (
    .A(_10195_),
    .B(_10194_),
    .C(_10197_),
    .Y(_10202_)
);

NAND3X1 _20223_ (
    .A(_10190_),
    .B(_10181_),
    .C(_10192_),
    .Y(_10203_)
);

NAND3X1 _20224_ (
    .A(_10201_),
    .B(_10203_),
    .C(_10202_),
    .Y(_10204_)
);

NAND2X1 _20225_ (
    .A(_10204_),
    .B(_10199_),
    .Y(_10205_)
);

NAND2X1 _20226_ (
    .A(_9918_),
    .B(_9919_),
    .Y(_10206_)
);

NAND2X1 _20227_ (
    .A(_9921_),
    .B(_9920_),
    .Y(_10207_)
);

OAI21X1 _20228_ (
    .A(_10206_),
    .B(_10207_),
    .C(_9920_),
    .Y(_10208_)
);

AND2X2 _20229_ (
    .A(_9884_),
    .B(_9876_),
    .Y(_10209_)
);

NAND3X1 _20230_ (
    .A(_9908_),
    .B(_9910_),
    .C(_9902_),
    .Y(_10210_)
);

NAND2X1 _20231_ (
    .A(breg_14_bF$buf1),
    .B(areg_24_bF$buf0),
    .Y(_10211_)
);

NAND2X1 _20232_ (
    .A(breg_12_bF$buf2),
    .B(areg_26_bF$buf2),
    .Y(_10212_)
);

XOR2X1 _20233_ (
    .A(_10157_),
    .B(_10212_),
    .Y(_10213_)
);

XNOR2X1 _20234_ (
    .A(_10213_),
    .B(_10211_),
    .Y(_10214_)
);

OAI21X1 _20235_ (
    .A(_9874_),
    .B(_9863_),
    .C(_9867_),
    .Y(_10215_)
);

NAND2X1 _20236_ (
    .A(breg_11_bF$buf4),
    .B(areg_27_bF$buf5),
    .Y(_10216_)
);

INVX2 _20237_ (
    .A(_10216_),
    .Y(_10217_)
);

AND2X2 _20238_ (
    .A(breg_10_bF$buf2),
    .B(areg_28_bF$buf0),
    .Y(_10218_)
);

AND2X2 _20239_ (
    .A(breg_9_bF$buf5),
    .B(areg_29_bF$buf5),
    .Y(_10219_)
);

NAND2X1 _20240_ (
    .A(_10218_),
    .B(_10219_),
    .Y(_10220_)
);

NAND2X1 _20241_ (
    .A(breg_9_bF$buf4),
    .B(areg_29_bF$buf4),
    .Y(_10222_)
);

OAI21X1 _20242_ (
    .A(_7217__bF$buf1),
    .B(_7520__bF$buf0),
    .C(_10222_),
    .Y(_10223_)
);

NAND3X1 _20243_ (
    .A(_10217_),
    .B(_10223_),
    .C(_10220_),
    .Y(_10224_)
);

NAND2X1 _20244_ (
    .A(breg_10_bF$buf1),
    .B(areg_29_bF$buf3),
    .Y(_10225_)
);

NOR2X1 _20245_ (
    .A(_9871_),
    .B(_10225_),
    .Y(_10226_)
);

NOR2X1 _20246_ (
    .A(_10218_),
    .B(_10219_),
    .Y(_10227_)
);

OAI21X1 _20247_ (
    .A(_10227_),
    .B(_10226_),
    .C(_10216_),
    .Y(_10228_)
);

NAND3X1 _20248_ (
    .A(_10224_),
    .B(_10215_),
    .C(_10228_),
    .Y(_10229_)
);

AOI21X1 _20249_ (
    .A(_9864_),
    .B(_9869_),
    .C(_9873_),
    .Y(_10230_)
);

OAI21X1 _20250_ (
    .A(_7217__bF$buf0),
    .B(_7520__bF$buf3),
    .C(_10219_),
    .Y(_10231_)
);

OAI21X1 _20251_ (
    .A(_6044__bF$buf1),
    .B(_9153_),
    .C(_10218_),
    .Y(_10234_)
);

AOI21X1 _20252_ (
    .A(_10231_),
    .B(_10234_),
    .C(_10216_),
    .Y(_10235_)
);

AOI21X1 _20253_ (
    .A(_10223_),
    .B(_10220_),
    .C(_10217_),
    .Y(_10236_)
);

OAI21X1 _20254_ (
    .A(_10235_),
    .B(_10236_),
    .C(_10230_),
    .Y(_10237_)
);

NAND3X1 _20255_ (
    .A(_10229_),
    .B(_10237_),
    .C(_10214_),
    .Y(_10238_)
);

INVX2 _20256_ (
    .A(_10211_),
    .Y(_10239_)
);

XNOR2X1 _20257_ (
    .A(_10213_),
    .B(_10239_),
    .Y(_10240_)
);

OAI21X1 _20258_ (
    .A(_10235_),
    .B(_10236_),
    .C(_10215_),
    .Y(_10241_)
);

NAND3X1 _20259_ (
    .A(_10230_),
    .B(_10224_),
    .C(_10228_),
    .Y(_10242_)
);

NAND3X1 _20260_ (
    .A(_10241_),
    .B(_10242_),
    .C(_10240_),
    .Y(_10243_)
);

NAND3X1 _20261_ (
    .A(_10210_),
    .B(_10238_),
    .C(_10243_),
    .Y(_10245_)
);

AOI21X1 _20262_ (
    .A(_9536_),
    .B(_9539_),
    .C(_9911_),
    .Y(_10246_)
);

AOI21X1 _20263_ (
    .A(_10241_),
    .B(_10242_),
    .C(_10240_),
    .Y(_10247_)
);

AOI21X1 _20264_ (
    .A(_10229_),
    .B(_10237_),
    .C(_10214_),
    .Y(_10248_)
);

OAI21X1 _20265_ (
    .A(_10247_),
    .B(_10248_),
    .C(_10246_),
    .Y(_10249_)
);

AOI21X1 _20266_ (
    .A(_10245_),
    .B(_10249_),
    .C(_10209_),
    .Y(_10250_)
);

NAND2X1 _20267_ (
    .A(_9876_),
    .B(_9884_),
    .Y(_10251_)
);

NAND3X1 _20268_ (
    .A(_10246_),
    .B(_10238_),
    .C(_10243_),
    .Y(_10252_)
);

OAI21X1 _20269_ (
    .A(_10247_),
    .B(_10248_),
    .C(_10210_),
    .Y(_10253_)
);

AOI21X1 _20270_ (
    .A(_10252_),
    .B(_10253_),
    .C(_10251_),
    .Y(_10254_)
);

OAI21X1 _20271_ (
    .A(_9901_),
    .B(_9905_),
    .C(_9908_),
    .Y(_10256_)
);

NAND2X1 _20272_ (
    .A(breg[8]),
    .B(areg_31_bF$buf2),
    .Y(_10257_)
);

NOR2X1 _20273_ (
    .A(_9901_),
    .B(_10257_),
    .Y(_10258_)
);

AOI22X1 _20274_ (
    .A(breg_7_bF$buf4),
    .B(areg_31_bF$buf1),
    .C(breg[8]),
    .D(areg_30_bF$buf2),
    .Y(_10259_)
);

NOR2X1 _20275_ (
    .A(_10259_),
    .B(_10258_),
    .Y(_10260_)
);

NOR2X1 _20276_ (
    .A(_10260_),
    .B(_10256_),
    .Y(_10261_)
);

NAND2X1 _20277_ (
    .A(_10260_),
    .B(_10256_),
    .Y(_10262_)
);

INVX2 _20278_ (
    .A(_10262_),
    .Y(_10263_)
);

NOR2X1 _20279_ (
    .A(_10261_),
    .B(_10263_),
    .Y(_10264_)
);

INVX1 _20280_ (
    .A(_10264_),
    .Y(_10265_)
);

OAI21X1 _20281_ (
    .A(_10250_),
    .B(_10254_),
    .C(_10265_),
    .Y(_10267_)
);

NAND3X1 _20282_ (
    .A(_10251_),
    .B(_10252_),
    .C(_10253_),
    .Y(_10268_)
);

NAND3X1 _20283_ (
    .A(_10245_),
    .B(_10209_),
    .C(_10249_),
    .Y(_10269_)
);

NAND3X1 _20284_ (
    .A(_10264_),
    .B(_10268_),
    .C(_10269_),
    .Y(_10270_)
);

NAND3X1 _20285_ (
    .A(_10267_),
    .B(_10270_),
    .C(_10208_),
    .Y(_10271_)
);

AOI21X1 _20286_ (
    .A(_9555_),
    .B(_9912_),
    .C(_9917_),
    .Y(_10272_)
);

NAND2X1 _20287_ (
    .A(_10270_),
    .B(_10267_),
    .Y(_10273_)
);

NAND2X1 _20288_ (
    .A(_10273_),
    .B(_10272_),
    .Y(_10274_)
);

NAND3X1 _20289_ (
    .A(_10271_),
    .B(_10274_),
    .C(_10205_),
    .Y(_10275_)
);

NAND3X1 _20290_ (
    .A(_10110_),
    .B(_10203_),
    .C(_10202_),
    .Y(_10276_)
);

OAI21X1 _20291_ (
    .A(_10198_),
    .B(_10193_),
    .C(_10201_),
    .Y(_10278_)
);

NAND2X1 _20292_ (
    .A(_10276_),
    .B(_10278_),
    .Y(_10279_)
);

NOR2X1 _20293_ (
    .A(_10273_),
    .B(_10272_),
    .Y(_10280_)
);

AOI21X1 _20294_ (
    .A(_10267_),
    .B(_10270_),
    .C(_10208_),
    .Y(_10281_)
);

OAI21X1 _20295_ (
    .A(_10280_),
    .B(_10281_),
    .C(_10279_),
    .Y(_10282_)
);

NAND3X1 _20296_ (
    .A(_10282_),
    .B(_10275_),
    .C(_10109_),
    .Y(_10283_)
);

AOI21X1 _20297_ (
    .A(_9935_),
    .B(_9933_),
    .C(_9942_),
    .Y(_10284_)
);

NAND2X1 _20298_ (
    .A(_10208_),
    .B(_10273_),
    .Y(_10285_)
);

OR2X2 _20299_ (
    .A(_10273_),
    .B(_10208_),
    .Y(_10286_)
);

AOI21X1 _20300_ (
    .A(_10285_),
    .B(_10286_),
    .C(_10279_),
    .Y(_10287_)
);

AOI21X1 _20301_ (
    .A(_10271_),
    .B(_10274_),
    .C(_10205_),
    .Y(_10289_)
);

OAI21X1 _20302_ (
    .A(_10287_),
    .B(_10289_),
    .C(_10284_),
    .Y(_10290_)
);

NAND3X1 _20303_ (
    .A(_10283_),
    .B(_10290_),
    .C(_10108_),
    .Y(_10291_)
);

NAND3X1 _20304_ (
    .A(_10104_),
    .B(_10097_),
    .C(_10102_),
    .Y(_10292_)
);

NAND3X1 _20305_ (
    .A(_10105_),
    .B(_9999_),
    .C(_10106_),
    .Y(_10293_)
);

NAND2X1 _20306_ (
    .A(_10292_),
    .B(_10293_),
    .Y(_10294_)
);

OAI21X1 _20307_ (
    .A(_10287_),
    .B(_10289_),
    .C(_10109_),
    .Y(_10295_)
);

NAND3X1 _20308_ (
    .A(_10282_),
    .B(_10275_),
    .C(_10284_),
    .Y(_10296_)
);

NAND3X1 _20309_ (
    .A(_10296_),
    .B(_10295_),
    .C(_10294_),
    .Y(_10297_)
);

NAND3X1 _20310_ (
    .A(_10291_),
    .B(_10297_),
    .C(_9998_),
    .Y(_10298_)
);

NOR3X1 _20311_ (
    .A(_9930_),
    .B(_9936_),
    .C(_9940_),
    .Y(_10300_)
);

AOI21X1 _20312_ (
    .A(_9950_),
    .B(_9952_),
    .C(_10300_),
    .Y(_10301_)
);

AOI21X1 _20313_ (
    .A(_10296_),
    .B(_10295_),
    .C(_10294_),
    .Y(_10302_)
);

AOI21X1 _20314_ (
    .A(_10283_),
    .B(_10290_),
    .C(_10108_),
    .Y(_10303_)
);

OAI21X1 _20315_ (
    .A(_10302_),
    .B(_10303_),
    .C(_10301_),
    .Y(_10304_)
);

NAND3X1 _20316_ (
    .A(_9996_),
    .B(_10304_),
    .C(_10298_),
    .Y(_10305_)
);

INVX2 _20317_ (
    .A(_9996_),
    .Y(_10306_)
);

OAI21X1 _20318_ (
    .A(_10302_),
    .B(_10303_),
    .C(_9998_),
    .Y(_10307_)
);

NAND3X1 _20319_ (
    .A(_10291_),
    .B(_10297_),
    .C(_10301_),
    .Y(_10308_)
);

NAND3X1 _20320_ (
    .A(_10306_),
    .B(_10307_),
    .C(_10308_),
    .Y(_10309_)
);

NAND3X1 _20321_ (
    .A(_10305_),
    .B(_10309_),
    .C(_9995_),
    .Y(_10311_)
);

NOR3X1 _20322_ (
    .A(_9946_),
    .B(_9953_),
    .C(_9956_),
    .Y(_10312_)
);

AOI21X1 _20323_ (
    .A(_9640_),
    .B(_9963_),
    .C(_10312_),
    .Y(_10313_)
);

AOI21X1 _20324_ (
    .A(_10307_),
    .B(_10308_),
    .C(_10306_),
    .Y(_10314_)
);

AOI21X1 _20325_ (
    .A(_10304_),
    .B(_10298_),
    .C(_9996_),
    .Y(_10315_)
);

OAI21X1 _20326_ (
    .A(_10314_),
    .B(_10315_),
    .C(_10313_),
    .Y(_10316_)
);

NAND3X1 _20327_ (
    .A(_9993_),
    .B(_10311_),
    .C(_10316_),
    .Y(_10317_)
);

INVX2 _20328_ (
    .A(_9993_),
    .Y(_10318_)
);

OAI21X1 _20329_ (
    .A(_10314_),
    .B(_10315_),
    .C(_9995_),
    .Y(_10319_)
);

NAND3X1 _20330_ (
    .A(_10305_),
    .B(_10309_),
    .C(_10313_),
    .Y(_10320_)
);

NAND3X1 _20331_ (
    .A(_10318_),
    .B(_10319_),
    .C(_10320_),
    .Y(_10322_)
);

AOI21X1 _20332_ (
    .A(_10317_),
    .B(_10322_),
    .C(_9992_),
    .Y(_10323_)
);

AOI21X1 _20333_ (
    .A(_9967_),
    .B(_9968_),
    .C(_9639_),
    .Y(_10324_)
);

OAI21X1 _20334_ (
    .A(_10324_),
    .B(_9638_),
    .C(_9972_),
    .Y(_10325_)
);

AOI21X1 _20335_ (
    .A(_10319_),
    .B(_10320_),
    .C(_10318_),
    .Y(_10326_)
);

AOI21X1 _20336_ (
    .A(_10311_),
    .B(_10316_),
    .C(_9993_),
    .Y(_10327_)
);

NOR3X1 _20337_ (
    .A(_10327_),
    .B(_10325_),
    .C(_10326_),
    .Y(_10328_)
);

OAI21X1 _20338_ (
    .A(_10323_),
    .B(_10328_),
    .C(_9989_),
    .Y(_10329_)
);

INVX1 _20339_ (
    .A(_10329_),
    .Y(_10330_)
);

OAI21X1 _20340_ (
    .A(_10326_),
    .B(_10327_),
    .C(_10325_),
    .Y(_10331_)
);

NAND3X1 _20341_ (
    .A(_10317_),
    .B(_10322_),
    .C(_9992_),
    .Y(_10333_)
);

NAND2X1 _20342_ (
    .A(_10331_),
    .B(_10333_),
    .Y(_10334_)
);

NOR2X1 _20343_ (
    .A(_10334_),
    .B(_9989_),
    .Y(_10335_)
);

NOR2X1 _20344_ (
    .A(_10335_),
    .B(_10330_),
    .Y(_0_[38])
);

NAND2X1 _20345_ (
    .A(_10317_),
    .B(_10322_),
    .Y(_10336_)
);

OAI21X1 _20346_ (
    .A(_9992_),
    .B(_10336_),
    .C(_10329_),
    .Y(_10337_)
);

AOI21X1 _20347_ (
    .A(_10305_),
    .B(_10309_),
    .C(_9995_),
    .Y(_10338_)
);

OAI21X1 _20348_ (
    .A(_10338_),
    .B(_10318_),
    .C(_10311_),
    .Y(_10339_)
);

OAI21X1 _20349_ (
    .A(_10031_),
    .B(_10001_),
    .C(_10039_),
    .Y(_10340_)
);

INVX1 _20350_ (
    .A(_10340_),
    .Y(_10341_)
);

AOI21X1 _20351_ (
    .A(_10291_),
    .B(_10297_),
    .C(_9998_),
    .Y(_10343_)
);

OAI21X1 _20352_ (
    .A(_10343_),
    .B(_10306_),
    .C(_10298_),
    .Y(_10344_)
);

NAND2X1 _20353_ (
    .A(_10097_),
    .B(_10292_),
    .Y(_10345_)
);

INVX2 _20354_ (
    .A(_10345_),
    .Y(_10346_)
);

AOI21X1 _20355_ (
    .A(_10282_),
    .B(_10275_),
    .C(_10109_),
    .Y(_10347_)
);

OAI21X1 _20356_ (
    .A(_10294_),
    .B(_10347_),
    .C(_10283_),
    .Y(_10348_)
);

NAND2X1 _20357_ (
    .A(_10083_),
    .B(_10091_),
    .Y(_10349_)
);

NOR2X1 _20358_ (
    .A(_5190__bF$buf0),
    .B(_7225__bF$buf1),
    .Y(_10350_)
);

INVX1 _20359_ (
    .A(_10350_),
    .Y(_10351_)
);

OAI21X1 _20360_ (
    .A(_10019_),
    .B(_10005_),
    .C(_10029_),
    .Y(_10352_)
);

NOR2X1 _20361_ (
    .A(_6582__bF$buf0),
    .B(_6815__bF$buf0),
    .Y(_10354_)
);

INVX2 _20362_ (
    .A(_10354_),
    .Y(_10355_)
);

OAI21X1 _20363_ (
    .A(_10017_),
    .B(_10007_),
    .C(_10011_),
    .Y(_10356_)
);

NAND2X1 _20364_ (
    .A(areg_10_bF$buf2),
    .B(breg_29_bF$buf4),
    .Y(_10357_)
);

INVX2 _20365_ (
    .A(_10357_),
    .Y(_10358_)
);

AND2X2 _20366_ (
    .A(areg_11_bF$buf2),
    .B(breg_28_bF$buf1),
    .Y(_10359_)
);

AND2X2 _20367_ (
    .A(areg_12_bF$buf4),
    .B(breg_27_bF$buf1),
    .Y(_10360_)
);

NAND2X1 _20368_ (
    .A(_10359_),
    .B(_10360_),
    .Y(_10361_)
);

OAI22X1 _20369_ (
    .A(_9104__bF$buf3),
    .B(_6050__bF$buf3),
    .C(_10869__bF$buf1),
    .D(_5668__bF$buf5),
    .Y(_10362_)
);

NAND3X1 _20370_ (
    .A(_10358_),
    .B(_10362_),
    .C(_10361_),
    .Y(_10363_)
);

NAND2X1 _20371_ (
    .A(areg_12_bF$buf3),
    .B(breg_28_bF$buf0),
    .Y(_10365_)
);

NOR2X1 _20372_ (
    .A(_10015_),
    .B(_10365_),
    .Y(_10366_)
);

NOR2X1 _20373_ (
    .A(_10359_),
    .B(_10360_),
    .Y(_10367_)
);

OAI21X1 _20374_ (
    .A(_10367_),
    .B(_10366_),
    .C(_10357_),
    .Y(_10368_)
);

AOI21X1 _20375_ (
    .A(_10363_),
    .B(_10368_),
    .C(_10356_),
    .Y(_10369_)
);

AOI21X1 _20376_ (
    .A(_10008_),
    .B(_10012_),
    .C(_10016_),
    .Y(_10370_)
);

OAI21X1 _20377_ (
    .A(_9104__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_10360_),
    .Y(_10371_)
);

OAI21X1 _20378_ (
    .A(_10869__bF$buf0),
    .B(_5668__bF$buf4),
    .C(_10359_),
    .Y(_10372_)
);

AOI21X1 _20379_ (
    .A(_10371_),
    .B(_10372_),
    .C(_10357_),
    .Y(_10373_)
);

AOI21X1 _20380_ (
    .A(_10362_),
    .B(_10361_),
    .C(_10358_),
    .Y(_10374_)
);

NOR3X1 _20381_ (
    .A(_10374_),
    .B(_10370_),
    .C(_10373_),
    .Y(_10376_)
);

OAI21X1 _20382_ (
    .A(_10376_),
    .B(_10369_),
    .C(_10355_),
    .Y(_10377_)
);

OAI21X1 _20383_ (
    .A(_10373_),
    .B(_10374_),
    .C(_10370_),
    .Y(_10378_)
);

NAND3X1 _20384_ (
    .A(_10363_),
    .B(_10356_),
    .C(_10368_),
    .Y(_10379_)
);

NAND3X1 _20385_ (
    .A(_10354_),
    .B(_10378_),
    .C(_10379_),
    .Y(_10380_)
);

AOI21X1 _20386_ (
    .A(_10380_),
    .B(_10377_),
    .C(_10352_),
    .Y(_10381_)
);

AOI21X1 _20387_ (
    .A(_10004_),
    .B(_10028_),
    .C(_10026_),
    .Y(_10382_)
);

AOI21X1 _20388_ (
    .A(_10378_),
    .B(_10379_),
    .C(_10354_),
    .Y(_10383_)
);

NOR3X1 _20389_ (
    .A(_10369_),
    .B(_10355_),
    .C(_10376_),
    .Y(_10384_)
);

NOR3X1 _20390_ (
    .A(_10382_),
    .B(_10383_),
    .C(_10384_),
    .Y(_10385_)
);

OAI21X1 _20391_ (
    .A(_10385_),
    .B(_10381_),
    .C(_10351_),
    .Y(_10387_)
);

OAI21X1 _20392_ (
    .A(_10384_),
    .B(_10383_),
    .C(_10382_),
    .Y(_10388_)
);

NAND3X1 _20393_ (
    .A(_10352_),
    .B(_10380_),
    .C(_10377_),
    .Y(_10389_)
);

NAND3X1 _20394_ (
    .A(_10350_),
    .B(_10389_),
    .C(_10388_),
    .Y(_10390_)
);

AND2X2 _20395_ (
    .A(_10387_),
    .B(_10390_),
    .Y(_10391_)
);

OAI21X1 _20396_ (
    .A(_10081_),
    .B(_10078_),
    .C(_10072_),
    .Y(_10392_)
);

NAND2X1 _20397_ (
    .A(_10059_),
    .B(_10065_),
    .Y(_10393_)
);

OAI21X1 _20398_ (
    .A(_10050_),
    .B(_10045_),
    .C(_10053_),
    .Y(_10394_)
);

NAND2X1 _20399_ (
    .A(areg_13_bF$buf2),
    .B(breg_26_bF$buf1),
    .Y(_10395_)
);

NAND2X1 _20400_ (
    .A(areg_14_bF$buf1),
    .B(breg_25_bF$buf4),
    .Y(_10396_)
);

NAND2X1 _20401_ (
    .A(areg_15_bF$buf4),
    .B(breg_24_bF$buf5),
    .Y(_10398_)
);

NOR2X1 _20402_ (
    .A(_10396_),
    .B(_10398_),
    .Y(_10399_)
);

AND2X2 _20403_ (
    .A(_10396_),
    .B(_10398_),
    .Y(_10400_)
);

OAI21X1 _20404_ (
    .A(_10400_),
    .B(_10399_),
    .C(_10395_),
    .Y(_10401_)
);

INVX1 _20405_ (
    .A(_10395_),
    .Y(_10402_)
);

OR2X2 _20406_ (
    .A(_10396_),
    .B(_10398_),
    .Y(_10403_)
);

OAI21X1 _20407_ (
    .A(_2465__bF$buf4),
    .B(_5315__bF$buf4),
    .C(_10396_),
    .Y(_10404_)
);

NAND3X1 _20408_ (
    .A(_10402_),
    .B(_10404_),
    .C(_10403_),
    .Y(_10405_)
);

NAND2X1 _20409_ (
    .A(areg_17_bF$buf2),
    .B(breg_22_bF$buf2),
    .Y(_10406_)
);

AND2X2 _20410_ (
    .A(_10056_),
    .B(_10114_),
    .Y(_10407_)
);

OAI22X1 _20411_ (
    .A(_9759_),
    .B(_10406_),
    .C(_10407_),
    .D(_10111_),
    .Y(_10409_)
);

NAND3X1 _20412_ (
    .A(_10401_),
    .B(_10405_),
    .C(_10409_),
    .Y(_10410_)
);

AOI21X1 _20413_ (
    .A(_10404_),
    .B(_10403_),
    .C(_10402_),
    .Y(_10411_)
);

NOR3X1 _20414_ (
    .A(_10395_),
    .B(_10399_),
    .C(_10400_),
    .Y(_10412_)
);

NOR2X1 _20415_ (
    .A(_10056_),
    .B(_10114_),
    .Y(_10413_)
);

OAI21X1 _20416_ (
    .A(_2884__bF$buf3),
    .B(_3781__bF$buf0),
    .C(_10056_),
    .Y(_10414_)
);

AOI21X1 _20417_ (
    .A(_10113_),
    .B(_10414_),
    .C(_10413_),
    .Y(_10415_)
);

OAI21X1 _20418_ (
    .A(_10412_),
    .B(_10411_),
    .C(_10415_),
    .Y(_10416_)
);

NAND3X1 _20419_ (
    .A(_10394_),
    .B(_10410_),
    .C(_10416_),
    .Y(_10417_)
);

INVX1 _20420_ (
    .A(_10394_),
    .Y(_10418_)
);

NAND3X1 _20421_ (
    .A(_10415_),
    .B(_10401_),
    .C(_10405_),
    .Y(_10420_)
);

OAI21X1 _20422_ (
    .A(_10412_),
    .B(_10411_),
    .C(_10409_),
    .Y(_10421_)
);

NAND3X1 _20423_ (
    .A(_10418_),
    .B(_10420_),
    .C(_10421_),
    .Y(_10422_)
);

OAI21X1 _20424_ (
    .A(_10116_),
    .B(_10184_),
    .C(_10138_),
    .Y(_10423_)
);

NAND3X1 _20425_ (
    .A(_10417_),
    .B(_10422_),
    .C(_10423_),
    .Y(_10424_)
);

AOI21X1 _20426_ (
    .A(_10420_),
    .B(_10421_),
    .C(_10418_),
    .Y(_10425_)
);

AOI21X1 _20427_ (
    .A(_10410_),
    .B(_10416_),
    .C(_10394_),
    .Y(_10426_)
);

AOI21X1 _20428_ (
    .A(_10139_),
    .B(_10137_),
    .C(_10183_),
    .Y(_10427_)
);

OAI21X1 _20429_ (
    .A(_10425_),
    .B(_10426_),
    .C(_10427_),
    .Y(_10428_)
);

NAND3X1 _20430_ (
    .A(_10393_),
    .B(_10428_),
    .C(_10424_),
    .Y(_10429_)
);

INVX2 _20431_ (
    .A(_10393_),
    .Y(_10431_)
);

NOR3X1 _20432_ (
    .A(_10425_),
    .B(_10426_),
    .C(_10427_),
    .Y(_10432_)
);

AOI21X1 _20433_ (
    .A(_10417_),
    .B(_10422_),
    .C(_10423_),
    .Y(_10433_)
);

OAI21X1 _20434_ (
    .A(_10432_),
    .B(_10433_),
    .C(_10431_),
    .Y(_10434_)
);

NAND3X1 _20435_ (
    .A(_10429_),
    .B(_10392_),
    .C(_10434_),
    .Y(_10435_)
);

AOI21X1 _20436_ (
    .A(_10043_),
    .B(_10076_),
    .C(_10080_),
    .Y(_10436_)
);

NAND3X1 _20437_ (
    .A(_10417_),
    .B(_10422_),
    .C(_10427_),
    .Y(_10437_)
);

OAI21X1 _20438_ (
    .A(_10425_),
    .B(_10426_),
    .C(_10423_),
    .Y(_10438_)
);

AOI21X1 _20439_ (
    .A(_10438_),
    .B(_10437_),
    .C(_10431_),
    .Y(_10439_)
);

AOI21X1 _20440_ (
    .A(_10428_),
    .B(_10424_),
    .C(_10393_),
    .Y(_10440_)
);

OAI21X1 _20441_ (
    .A(_10439_),
    .B(_10440_),
    .C(_10436_),
    .Y(_10442_)
);

NAND3X1 _20442_ (
    .A(_10435_),
    .B(_10442_),
    .C(_10391_),
    .Y(_10443_)
);

NAND2X1 _20443_ (
    .A(_10390_),
    .B(_10387_),
    .Y(_10444_)
);

OAI21X1 _20444_ (
    .A(_10439_),
    .B(_10440_),
    .C(_10392_),
    .Y(_10445_)
);

NAND3X1 _20445_ (
    .A(_10429_),
    .B(_10434_),
    .C(_10436_),
    .Y(_10446_)
);

NAND3X1 _20446_ (
    .A(_10444_),
    .B(_10445_),
    .C(_10446_),
    .Y(_10447_)
);

OAI21X1 _20447_ (
    .A(_10201_),
    .B(_10193_),
    .C(_10203_),
    .Y(_10448_)
);

NAND3X1 _20448_ (
    .A(_10447_),
    .B(_10448_),
    .C(_10443_),
    .Y(_10449_)
);

AOI21X1 _20449_ (
    .A(_10445_),
    .B(_10446_),
    .C(_10444_),
    .Y(_10450_)
);

AOI21X1 _20450_ (
    .A(_10435_),
    .B(_10442_),
    .C(_10391_),
    .Y(_10451_)
);

AOI21X1 _20451_ (
    .A(_10110_),
    .B(_10202_),
    .C(_10198_),
    .Y(_10453_)
);

OAI21X1 _20452_ (
    .A(_10451_),
    .B(_10450_),
    .C(_10453_),
    .Y(_10454_)
);

NAND3X1 _20453_ (
    .A(_10349_),
    .B(_10449_),
    .C(_10454_),
    .Y(_10455_)
);

AND2X2 _20454_ (
    .A(_10091_),
    .B(_10083_),
    .Y(_10456_)
);

NAND3X1 _20455_ (
    .A(_10447_),
    .B(_10453_),
    .C(_10443_),
    .Y(_10457_)
);

OAI21X1 _20456_ (
    .A(_10451_),
    .B(_10450_),
    .C(_10448_),
    .Y(_10458_)
);

NAND3X1 _20457_ (
    .A(_10457_),
    .B(_10458_),
    .C(_10456_),
    .Y(_10459_)
);

NAND2X1 _20458_ (
    .A(_10455_),
    .B(_10459_),
    .Y(_10460_)
);

OAI21X1 _20459_ (
    .A(_10279_),
    .B(_10281_),
    .C(_10271_),
    .Y(_10461_)
);

NAND2X1 _20460_ (
    .A(_10173_),
    .B(_10181_),
    .Y(_10462_)
);

NAND2X1 _20461_ (
    .A(areg_16_bF$buf2),
    .B(breg_23_bF$buf3),
    .Y(_10464_)
);

INVX2 _20462_ (
    .A(_10464_),
    .Y(_10465_)
);

NAND2X1 _20463_ (
    .A(areg_18_bF$buf2),
    .B(breg_21_bF$buf2),
    .Y(_10466_)
);

XOR2X1 _20464_ (
    .A(_10406_),
    .B(_10466_),
    .Y(_10467_)
);

XNOR2X1 _20465_ (
    .A(_10467_),
    .B(_10465_),
    .Y(_10468_)
);

OAI21X1 _20466_ (
    .A(_10124_),
    .B(_10118_),
    .C(_10127_),
    .Y(_10469_)
);

NAND2X1 _20467_ (
    .A(areg_19_bF$buf4),
    .B(breg_20_bF$buf3),
    .Y(_10470_)
);

AND2X2 _20468_ (
    .A(breg_18_bF$buf1),
    .B(areg_21_bF$buf3),
    .Y(_10471_)
);

OAI21X1 _20469_ (
    .A(_3253__bF$buf3),
    .B(_3958__bF$buf2),
    .C(_10471_),
    .Y(_10472_)
);

AND2X2 _20470_ (
    .A(breg_19_bF$buf1),
    .B(areg_20_bF$buf4),
    .Y(_10473_)
);

OAI21X1 _20471_ (
    .A(_3529__bF$buf2),
    .B(_3961__bF$buf4),
    .C(_10473_),
    .Y(_10475_)
);

AOI21X1 _20472_ (
    .A(_10472_),
    .B(_10475_),
    .C(_10470_),
    .Y(_10476_)
);

INVX2 _20473_ (
    .A(_10470_),
    .Y(_10477_)
);

NAND2X1 _20474_ (
    .A(_10473_),
    .B(_10471_),
    .Y(_10478_)
);

OAI21X1 _20475_ (
    .A(_3529__bF$buf1),
    .B(_3961__bF$buf3),
    .C(_10119_),
    .Y(_10479_)
);

AOI21X1 _20476_ (
    .A(_10479_),
    .B(_10478_),
    .C(_10477_),
    .Y(_10480_)
);

OAI21X1 _20477_ (
    .A(_10476_),
    .B(_10480_),
    .C(_10469_),
    .Y(_10481_)
);

AOI21X1 _20478_ (
    .A(_10126_),
    .B(_10128_),
    .C(_10120_),
    .Y(_10482_)
);

NAND3X1 _20479_ (
    .A(_10477_),
    .B(_10479_),
    .C(_10478_),
    .Y(_10483_)
);

NAND2X1 _20480_ (
    .A(breg_18_bF$buf0),
    .B(areg_21_bF$buf2),
    .Y(_10484_)
);

NOR2X1 _20481_ (
    .A(_10119_),
    .B(_10484_),
    .Y(_10486_)
);

NOR2X1 _20482_ (
    .A(_10473_),
    .B(_10471_),
    .Y(_10487_)
);

OAI21X1 _20483_ (
    .A(_10487_),
    .B(_10486_),
    .C(_10470_),
    .Y(_10488_)
);

NAND3X1 _20484_ (
    .A(_10482_),
    .B(_10483_),
    .C(_10488_),
    .Y(_10489_)
);

AOI21X1 _20485_ (
    .A(_10481_),
    .B(_10489_),
    .C(_10468_),
    .Y(_10490_)
);

XNOR2X1 _20486_ (
    .A(_10467_),
    .B(_10464_),
    .Y(_10491_)
);

NAND3X1 _20487_ (
    .A(_10483_),
    .B(_10469_),
    .C(_10488_),
    .Y(_10492_)
);

OAI21X1 _20488_ (
    .A(_10476_),
    .B(_10480_),
    .C(_10482_),
    .Y(_10493_)
);

AOI21X1 _20489_ (
    .A(_10493_),
    .B(_10492_),
    .C(_10491_),
    .Y(_10494_)
);

NOR2X1 _20490_ (
    .A(_10490_),
    .B(_10494_),
    .Y(_10495_)
);

OAI21X1 _20491_ (
    .A(_10171_),
    .B(_10169_),
    .C(_10160_),
    .Y(_10497_)
);

INVX1 _20492_ (
    .A(_10149_),
    .Y(_10498_)
);

OAI21X1 _20493_ (
    .A(_10143_),
    .B(_10498_),
    .C(_10152_),
    .Y(_10499_)
);

NAND2X1 _20494_ (
    .A(breg_17_bF$buf1),
    .B(areg_22_bF$buf2),
    .Y(_10500_)
);

INVX1 _20495_ (
    .A(_10500_),
    .Y(_10501_)
);

AND2X2 _20496_ (
    .A(breg_16_bF$buf1),
    .B(areg_23_bF$buf0),
    .Y(_10502_)
);

AND2X2 _20497_ (
    .A(breg_15_bF$buf3),
    .B(areg_24_bF$buf4),
    .Y(_10503_)
);

NAND2X1 _20498_ (
    .A(_10502_),
    .B(_10503_),
    .Y(_10504_)
);

OAI22X1 _20499_ (
    .A(_2362__bF$buf2),
    .B(_5921__bF$buf3),
    .C(_2560__bF$buf0),
    .D(_4541__bF$buf0),
    .Y(_10505_)
);

NAND3X1 _20500_ (
    .A(_10501_),
    .B(_10505_),
    .C(_10504_),
    .Y(_10506_)
);

OAI21X1 _20501_ (
    .A(_2560__bF$buf4),
    .B(_4541__bF$buf4),
    .C(_10503_),
    .Y(_10508_)
);

OAI21X1 _20502_ (
    .A(_2362__bF$buf1),
    .B(_5921__bF$buf2),
    .C(_10502_),
    .Y(_10509_)
);

NAND3X1 _20503_ (
    .A(_10500_),
    .B(_10508_),
    .C(_10509_),
    .Y(_10510_)
);

NAND2X1 _20504_ (
    .A(breg_13_bF$buf3),
    .B(areg_26_bF$buf1),
    .Y(_10511_)
);

AND2X2 _20505_ (
    .A(_10157_),
    .B(_10212_),
    .Y(_10512_)
);

OAI22X1 _20506_ (
    .A(_9858_),
    .B(_10511_),
    .C(_10512_),
    .D(_10211_),
    .Y(_10513_)
);

NAND3X1 _20507_ (
    .A(_10506_),
    .B(_10510_),
    .C(_10513_),
    .Y(_10514_)
);

AOI21X1 _20508_ (
    .A(_10508_),
    .B(_10509_),
    .C(_10500_),
    .Y(_10515_)
);

AOI21X1 _20509_ (
    .A(_10505_),
    .B(_10504_),
    .C(_10501_),
    .Y(_10516_)
);

NOR2X1 _20510_ (
    .A(_10157_),
    .B(_10212_),
    .Y(_10517_)
);

OAI21X1 _20511_ (
    .A(_2586__bF$buf2),
    .B(_6686__bF$buf1),
    .C(_10157_),
    .Y(_10519_)
);

AOI21X1 _20512_ (
    .A(_10239_),
    .B(_10519_),
    .C(_10517_),
    .Y(_10520_)
);

OAI21X1 _20513_ (
    .A(_10515_),
    .B(_10516_),
    .C(_10520_),
    .Y(_10521_)
);

NAND3X1 _20514_ (
    .A(_10499_),
    .B(_10514_),
    .C(_10521_),
    .Y(_10522_)
);

AOI21X1 _20515_ (
    .A(_9797_),
    .B(_10502_),
    .C(_10161_),
    .Y(_10523_)
);

NOR3X1 _20516_ (
    .A(_10516_),
    .B(_10520_),
    .C(_10515_),
    .Y(_10524_)
);

AOI21X1 _20517_ (
    .A(_10506_),
    .B(_10510_),
    .C(_10513_),
    .Y(_10525_)
);

OAI21X1 _20518_ (
    .A(_10524_),
    .B(_10525_),
    .C(_10523_),
    .Y(_10526_)
);

NAND3X1 _20519_ (
    .A(_10497_),
    .B(_10522_),
    .C(_10526_),
    .Y(_10527_)
);

AOI21X1 _20520_ (
    .A(_10144_),
    .B(_10166_),
    .C(_10170_),
    .Y(_10528_)
);

NAND3X1 _20521_ (
    .A(_10520_),
    .B(_10506_),
    .C(_10510_),
    .Y(_10530_)
);

OAI21X1 _20522_ (
    .A(_10515_),
    .B(_10516_),
    .C(_10513_),
    .Y(_10531_)
);

AOI21X1 _20523_ (
    .A(_10530_),
    .B(_10531_),
    .C(_10523_),
    .Y(_10532_)
);

AOI21X1 _20524_ (
    .A(_10514_),
    .B(_10521_),
    .C(_10499_),
    .Y(_10533_)
);

OAI21X1 _20525_ (
    .A(_10532_),
    .B(_10533_),
    .C(_10528_),
    .Y(_10534_)
);

NAND3X1 _20526_ (
    .A(_10495_),
    .B(_10534_),
    .C(_10527_),
    .Y(_10535_)
);

OR2X2 _20527_ (
    .A(_10490_),
    .B(_10494_),
    .Y(_10536_)
);

OAI21X1 _20528_ (
    .A(_10532_),
    .B(_10533_),
    .C(_10497_),
    .Y(_10537_)
);

NAND3X1 _20529_ (
    .A(_10528_),
    .B(_10522_),
    .C(_10526_),
    .Y(_10538_)
);

NAND3X1 _20530_ (
    .A(_10537_),
    .B(_10538_),
    .C(_10536_),
    .Y(_10539_)
);

AOI21X1 _20531_ (
    .A(_10238_),
    .B(_10243_),
    .C(_10246_),
    .Y(_10541_)
);

OAI21X1 _20532_ (
    .A(_10541_),
    .B(_10209_),
    .C(_10252_),
    .Y(_10542_)
);

NAND3X1 _20533_ (
    .A(_10535_),
    .B(_10539_),
    .C(_10542_),
    .Y(_10543_)
);

AOI21X1 _20534_ (
    .A(_10538_),
    .B(_10537_),
    .C(_10536_),
    .Y(_10544_)
);

AOI21X1 _20535_ (
    .A(_10534_),
    .B(_10527_),
    .C(_10495_),
    .Y(_10545_)
);

NOR3X1 _20536_ (
    .A(_10248_),
    .B(_10210_),
    .C(_10247_),
    .Y(_10546_)
);

AOI21X1 _20537_ (
    .A(_10251_),
    .B(_10253_),
    .C(_10546_),
    .Y(_10547_)
);

OAI21X1 _20538_ (
    .A(_10544_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10548_)
);

NAND3X1 _20539_ (
    .A(_10462_),
    .B(_10543_),
    .C(_10548_),
    .Y(_10549_)
);

AND2X2 _20540_ (
    .A(_10181_),
    .B(_10173_),
    .Y(_10550_)
);

NOR3X1 _20541_ (
    .A(_10544_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10552_)
);

AOI21X1 _20542_ (
    .A(_10535_),
    .B(_10539_),
    .C(_10542_),
    .Y(_10553_)
);

OAI21X1 _20543_ (
    .A(_10552_),
    .B(_10553_),
    .C(_10550_),
    .Y(_10554_)
);

NAND2X1 _20544_ (
    .A(_10549_),
    .B(_10554_),
    .Y(_10555_)
);

NAND2X1 _20545_ (
    .A(_10229_),
    .B(_10238_),
    .Y(_10556_)
);

NAND2X1 _20546_ (
    .A(breg_14_bF$buf0),
    .B(areg_25_bF$buf1),
    .Y(_10557_)
);

NAND2X1 _20547_ (
    .A(breg_12_bF$buf1),
    .B(areg_27_bF$buf4),
    .Y(_10558_)
);

XOR2X1 _20548_ (
    .A(_10511_),
    .B(_10558_),
    .Y(_10559_)
);

XNOR2X1 _20549_ (
    .A(_10559_),
    .B(_10557_),
    .Y(_10560_)
);

OAI21X1 _20550_ (
    .A(_10227_),
    .B(_10216_),
    .C(_10220_),
    .Y(_10561_)
);

NAND2X1 _20551_ (
    .A(breg_11_bF$buf3),
    .B(areg_28_bF$buf5),
    .Y(_10563_)
);

INVX2 _20552_ (
    .A(_10563_),
    .Y(_10564_)
);

AND2X2 _20553_ (
    .A(breg_10_bF$buf0),
    .B(areg_30_bF$buf1),
    .Y(_10565_)
);

NAND2X1 _20554_ (
    .A(_10219_),
    .B(_10565_),
    .Y(_10566_)
);

AOI22X1 _20555_ (
    .A(breg_9_bF$buf3),
    .B(areg_30_bF$buf0),
    .C(breg_10_bF$buf5),
    .D(areg_29_bF$buf2),
    .Y(_10567_)
);

INVX2 _20556_ (
    .A(_10567_),
    .Y(_10568_)
);

NAND3X1 _20557_ (
    .A(_10564_),
    .B(_10568_),
    .C(_10566_),
    .Y(_10569_)
);

NAND2X1 _20558_ (
    .A(breg_10_bF$buf4),
    .B(areg_30_bF$buf5),
    .Y(_10570_)
);

NOR2X1 _20559_ (
    .A(_10222_),
    .B(_10570_),
    .Y(_10571_)
);

OAI21X1 _20560_ (
    .A(_10571_),
    .B(_10567_),
    .C(_10563_),
    .Y(_10572_)
);

NAND3X1 _20561_ (
    .A(_10569_),
    .B(_10572_),
    .C(_10561_),
    .Y(_10574_)
);

AOI21X1 _20562_ (
    .A(_10217_),
    .B(_10223_),
    .C(_10226_),
    .Y(_10575_)
);

NOR3X1 _20563_ (
    .A(_10563_),
    .B(_10567_),
    .C(_10571_),
    .Y(_10576_)
);

AOI21X1 _20564_ (
    .A(_10568_),
    .B(_10566_),
    .C(_10564_),
    .Y(_10577_)
);

OAI21X1 _20565_ (
    .A(_10577_),
    .B(_10576_),
    .C(_10575_),
    .Y(_10578_)
);

NAND3X1 _20566_ (
    .A(_10574_),
    .B(_10578_),
    .C(_10560_),
    .Y(_10579_)
);

INVX2 _20567_ (
    .A(_10557_),
    .Y(_10580_)
);

XNOR2X1 _20568_ (
    .A(_10559_),
    .B(_10580_),
    .Y(_10581_)
);

OAI21X1 _20569_ (
    .A(_10577_),
    .B(_10576_),
    .C(_10561_),
    .Y(_10582_)
);

NAND3X1 _20570_ (
    .A(_10575_),
    .B(_10572_),
    .C(_10569_),
    .Y(_10583_)
);

NAND3X1 _20571_ (
    .A(_10582_),
    .B(_10583_),
    .C(_10581_),
    .Y(_10585_)
);

NAND3X1 _20572_ (
    .A(_10579_),
    .B(_10585_),
    .C(_10263_),
    .Y(_10586_)
);

AOI21X1 _20573_ (
    .A(_10582_),
    .B(_10583_),
    .C(_10581_),
    .Y(_10587_)
);

AOI21X1 _20574_ (
    .A(_10574_),
    .B(_10578_),
    .C(_10560_),
    .Y(_10588_)
);

OAI21X1 _20575_ (
    .A(_10587_),
    .B(_10588_),
    .C(_10262_),
    .Y(_10589_)
);

NAND3X1 _20576_ (
    .A(_10556_),
    .B(_10586_),
    .C(_10589_),
    .Y(_10590_)
);

AND2X2 _20577_ (
    .A(_10238_),
    .B(_10229_),
    .Y(_10591_)
);

NAND3X1 _20578_ (
    .A(_10262_),
    .B(_10579_),
    .C(_10585_),
    .Y(_10592_)
);

OAI21X1 _20579_ (
    .A(_10587_),
    .B(_10588_),
    .C(_10263_),
    .Y(_10593_)
);

NAND3X1 _20580_ (
    .A(_10592_),
    .B(_10591_),
    .C(_10593_),
    .Y(_10594_)
);

NOR2X1 _20581_ (
    .A(_10257_),
    .B(_9535_),
    .Y(_10596_)
);

AOI21X1 _20582_ (
    .A(_10594_),
    .B(_10590_),
    .C(_10596_),
    .Y(_10597_)
);

AOI21X1 _20583_ (
    .A(_10592_),
    .B(_10593_),
    .C(_10591_),
    .Y(_10598_)
);

AOI21X1 _20584_ (
    .A(_10586_),
    .B(_10589_),
    .C(_10556_),
    .Y(_10599_)
);

INVX1 _20585_ (
    .A(_10596_),
    .Y(_10600_)
);

NOR3X1 _20586_ (
    .A(_10598_),
    .B(_10600_),
    .C(_10599_),
    .Y(_10601_)
);

OAI21X1 _20587_ (
    .A(_10601_),
    .B(_10597_),
    .C(_10270_),
    .Y(_10602_)
);

NOR3X1 _20588_ (
    .A(_10250_),
    .B(_10265_),
    .C(_10254_),
    .Y(_10603_)
);

OAI21X1 _20589_ (
    .A(_10599_),
    .B(_10598_),
    .C(_10600_),
    .Y(_10604_)
);

NAND3X1 _20590_ (
    .A(_10596_),
    .B(_10594_),
    .C(_10590_),
    .Y(_10605_)
);

NAND3X1 _20591_ (
    .A(_10604_),
    .B(_10605_),
    .C(_10603_),
    .Y(_10607_)
);

NAND2X1 _20592_ (
    .A(_10607_),
    .B(_10602_),
    .Y(_10608_)
);

NOR2X1 _20593_ (
    .A(_10555_),
    .B(_10608_),
    .Y(_10609_)
);

NAND3X1 _20594_ (
    .A(_10535_),
    .B(_10539_),
    .C(_10547_),
    .Y(_10610_)
);

OAI21X1 _20595_ (
    .A(_10544_),
    .B(_10545_),
    .C(_10542_),
    .Y(_10611_)
);

AOI21X1 _20596_ (
    .A(_10611_),
    .B(_10610_),
    .C(_10550_),
    .Y(_10612_)
);

AOI21X1 _20597_ (
    .A(_10543_),
    .B(_10548_),
    .C(_10462_),
    .Y(_10613_)
);

NOR2X1 _20598_ (
    .A(_10613_),
    .B(_10612_),
    .Y(_10614_)
);

AOI21X1 _20599_ (
    .A(_10602_),
    .B(_10607_),
    .C(_10614_),
    .Y(_10615_)
);

OAI21X1 _20600_ (
    .A(_10609_),
    .B(_10615_),
    .C(_10461_),
    .Y(_10616_)
);

AOI21X1 _20601_ (
    .A(_10274_),
    .B(_10205_),
    .C(_10280_),
    .Y(_10618_)
);

NAND3X1 _20602_ (
    .A(_10602_),
    .B(_10607_),
    .C(_10614_),
    .Y(_10619_)
);

OAI21X1 _20603_ (
    .A(_10612_),
    .B(_10613_),
    .C(_10608_),
    .Y(_10620_)
);

NAND3X1 _20604_ (
    .A(_10619_),
    .B(_10620_),
    .C(_10618_),
    .Y(_10621_)
);

AOI21X1 _20605_ (
    .A(_10616_),
    .B(_10621_),
    .C(_10460_),
    .Y(_10622_)
);

NAND3X1 _20606_ (
    .A(_10449_),
    .B(_10454_),
    .C(_10456_),
    .Y(_10623_)
);

NAND3X1 _20607_ (
    .A(_10349_),
    .B(_10457_),
    .C(_10458_),
    .Y(_10624_)
);

NAND2X1 _20608_ (
    .A(_10624_),
    .B(_10623_),
    .Y(_10625_)
);

NAND3X1 _20609_ (
    .A(_10619_),
    .B(_10620_),
    .C(_10461_),
    .Y(_10626_)
);

OAI21X1 _20610_ (
    .A(_10609_),
    .B(_10615_),
    .C(_10618_),
    .Y(_10627_)
);

AOI21X1 _20611_ (
    .A(_10627_),
    .B(_10626_),
    .C(_10625_),
    .Y(_10629_)
);

OAI21X1 _20612_ (
    .A(_10622_),
    .B(_10629_),
    .C(_10348_),
    .Y(_10630_)
);

NOR3X1 _20613_ (
    .A(_10287_),
    .B(_10289_),
    .C(_10284_),
    .Y(_10631_)
);

AOI21X1 _20614_ (
    .A(_10108_),
    .B(_10290_),
    .C(_10631_),
    .Y(_10632_)
);

NAND3X1 _20615_ (
    .A(_10627_),
    .B(_10626_),
    .C(_10625_),
    .Y(_10633_)
);

NAND3X1 _20616_ (
    .A(_10616_),
    .B(_10621_),
    .C(_10460_),
    .Y(_10634_)
);

NAND3X1 _20617_ (
    .A(_10633_),
    .B(_10634_),
    .C(_10632_),
    .Y(_10635_)
);

AOI21X1 _20618_ (
    .A(_10630_),
    .B(_10635_),
    .C(_10346_),
    .Y(_10636_)
);

NAND3X1 _20619_ (
    .A(_10633_),
    .B(_10634_),
    .C(_10348_),
    .Y(_10637_)
);

OAI21X1 _20620_ (
    .A(_10622_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10638_)
);

AOI21X1 _20621_ (
    .A(_10637_),
    .B(_10638_),
    .C(_10345_),
    .Y(_10640_)
);

OAI21X1 _20622_ (
    .A(_10636_),
    .B(_10640_),
    .C(_10344_),
    .Y(_10641_)
);

NOR3X1 _20623_ (
    .A(_10302_),
    .B(_10303_),
    .C(_10301_),
    .Y(_10642_)
);

AOI21X1 _20624_ (
    .A(_10304_),
    .B(_9996_),
    .C(_10642_),
    .Y(_10643_)
);

NAND3X1 _20625_ (
    .A(_10345_),
    .B(_10637_),
    .C(_10638_),
    .Y(_10644_)
);

NOR3X1 _20626_ (
    .A(_10622_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10645_)
);

AOI21X1 _20627_ (
    .A(_10633_),
    .B(_10634_),
    .C(_10348_),
    .Y(_10646_)
);

OAI21X1 _20628_ (
    .A(_10645_),
    .B(_10646_),
    .C(_10346_),
    .Y(_10647_)
);

NAND3X1 _20629_ (
    .A(_10644_),
    .B(_10643_),
    .C(_10647_),
    .Y(_10648_)
);

AOI21X1 _20630_ (
    .A(_10641_),
    .B(_10648_),
    .C(_10341_),
    .Y(_10649_)
);

NAND3X1 _20631_ (
    .A(_10344_),
    .B(_10644_),
    .C(_10647_),
    .Y(_10651_)
);

OAI21X1 _20632_ (
    .A(_10636_),
    .B(_10640_),
    .C(_10643_),
    .Y(_10652_)
);

AOI21X1 _20633_ (
    .A(_10652_),
    .B(_10651_),
    .C(_10340_),
    .Y(_10653_)
);

OAI21X1 _20634_ (
    .A(_10649_),
    .B(_10653_),
    .C(_10339_),
    .Y(_10654_)
);

NOR3X1 _20635_ (
    .A(_10314_),
    .B(_10315_),
    .C(_10313_),
    .Y(_10655_)
);

AOI21X1 _20636_ (
    .A(_9993_),
    .B(_10316_),
    .C(_10655_),
    .Y(_10656_)
);

NAND3X1 _20637_ (
    .A(_10340_),
    .B(_10652_),
    .C(_10651_),
    .Y(_10657_)
);

NAND3X1 _20638_ (
    .A(_10341_),
    .B(_10641_),
    .C(_10648_),
    .Y(_10658_)
);

NAND3X1 _20639_ (
    .A(_10657_),
    .B(_10658_),
    .C(_10656_),
    .Y(_10659_)
);

NAND2X1 _20640_ (
    .A(_10659_),
    .B(_10654_),
    .Y(_10660_)
);

XOR2X1 _20641_ (
    .A(_10337_),
    .B(_10660_),
    .Y(_0_[39])
);

NOR3X1 _20642_ (
    .A(_8453_),
    .B(_8456_),
    .C(_8459_),
    .Y(_10662_)
);

OAI21X1 _20643_ (
    .A(_8068_),
    .B(_10662_),
    .C(_8466_),
    .Y(_10663_)
);

AOI21X1 _20644_ (
    .A(_8872_),
    .B(_8873_),
    .C(_8871_),
    .Y(_10664_)
);

NOR3X1 _20645_ (
    .A(_8868_),
    .B(_8473_),
    .C(_8865_),
    .Y(_10665_)
);

AOI21X1 _20646_ (
    .A(_9252_),
    .B(_9253_),
    .C(_9251_),
    .Y(_10666_)
);

NOR3X1 _20647_ (
    .A(_9244_),
    .B(_8881_),
    .C(_9248_),
    .Y(_10667_)
);

OAI22X1 _20648_ (
    .A(_10665_),
    .B(_10664_),
    .C(_10667_),
    .D(_10666_),
    .Y(_10668_)
);

NOR2X1 _20649_ (
    .A(_9251_),
    .B(_9258_),
    .Y(_10669_)
);

AOI21X1 _20650_ (
    .A(_9260_),
    .B(_8878_),
    .C(_10669_),
    .Y(_10670_)
);

OAI21X1 _20651_ (
    .A(_10668_),
    .B(_10663_),
    .C(_10670_),
    .Y(_10672_)
);

AOI22X1 _20652_ (
    .A(_10333_),
    .B(_10331_),
    .C(_10654_),
    .D(_10659_),
    .Y(_10673_)
);

AND2X2 _20653_ (
    .A(_9987_),
    .B(_10673_),
    .Y(_10674_)
);

AOI21X1 _20654_ (
    .A(_10657_),
    .B(_10658_),
    .C(_10339_),
    .Y(_10675_)
);

AOI21X1 _20655_ (
    .A(_10657_),
    .B(_10658_),
    .C(_10656_),
    .Y(_10676_)
);

NOR3X1 _20656_ (
    .A(_10649_),
    .B(_10339_),
    .C(_10653_),
    .Y(_10677_)
);

OAI22X1 _20657_ (
    .A(_10323_),
    .B(_10328_),
    .C(_10677_),
    .D(_10676_),
    .Y(_10678_)
);

NOR2X1 _20658_ (
    .A(_9992_),
    .B(_10336_),
    .Y(_10679_)
);

NOR3X1 _20659_ (
    .A(_10649_),
    .B(_10653_),
    .C(_10656_),
    .Y(_10680_)
);

NOR2X1 _20660_ (
    .A(_10680_),
    .B(_10679_),
    .Y(_10681_)
);

OAI22X1 _20661_ (
    .A(_9986_),
    .B(_10678_),
    .C(_10681_),
    .D(_10675_),
    .Y(_10683_)
);

AOI21X1 _20662_ (
    .A(_10674_),
    .B(_10672_),
    .C(_10683_),
    .Y(_10684_)
);

NAND2X1 _20663_ (
    .A(_10673_),
    .B(_9987_),
    .Y(_10685_)
);

NOR2X1 _20664_ (
    .A(_9264_),
    .B(_10685_),
    .Y(_10686_)
);

INVX1 _20665_ (
    .A(_10686_),
    .Y(_10687_)
);

OAI21X1 _20666_ (
    .A(_7651_),
    .B(_10687_),
    .C(_10684_),
    .Y(_10688_)
);

NOR3X1 _20667_ (
    .A(_10640_),
    .B(_10636_),
    .C(_10643_),
    .Y(_10689_)
);

OAI21X1 _20668_ (
    .A(_10381_),
    .B(_10351_),
    .C(_10389_),
    .Y(_10690_)
);

INVX2 _20669_ (
    .A(_10690_),
    .Y(_10691_)
);

OAI21X1 _20670_ (
    .A(_10646_),
    .B(_10346_),
    .C(_10637_),
    .Y(_10692_)
);

NAND2X1 _20671_ (
    .A(_10449_),
    .B(_10455_),
    .Y(_10694_)
);

INVX2 _20672_ (
    .A(_10694_),
    .Y(_10695_)
);

AOI21X1 _20673_ (
    .A(_10620_),
    .B(_10619_),
    .C(_10461_),
    .Y(_10696_)
);

OAI21X1 _20674_ (
    .A(_10460_),
    .B(_10696_),
    .C(_10626_),
    .Y(_10697_)
);

NAND2X1 _20675_ (
    .A(_10435_),
    .B(_10443_),
    .Y(_10698_)
);

NOR2X1 _20676_ (
    .A(_6582__bF$buf3),
    .B(_7225__bF$buf0),
    .Y(_10699_)
);

INVX1 _20677_ (
    .A(_10699_),
    .Y(_10700_)
);

OAI21X1 _20678_ (
    .A(_10369_),
    .B(_10355_),
    .C(_10379_),
    .Y(_10701_)
);

NOR2X1 _20679_ (
    .A(_7711__bF$buf0),
    .B(_6815__bF$buf4),
    .Y(_10702_)
);

INVX2 _20680_ (
    .A(_10702_),
    .Y(_10703_)
);

OAI21X1 _20681_ (
    .A(_10367_),
    .B(_10357_),
    .C(_10361_),
    .Y(_10705_)
);

NAND2X1 _20682_ (
    .A(areg_11_bF$buf1),
    .B(breg_29_bF$buf3),
    .Y(_10706_)
);

INVX2 _20683_ (
    .A(_10706_),
    .Y(_10707_)
);

AND2X2 _20684_ (
    .A(areg_12_bF$buf2),
    .B(breg_28_bF$buf5),
    .Y(_10708_)
);

AND2X2 _20685_ (
    .A(areg_13_bF$buf1),
    .B(breg_27_bF$buf0),
    .Y(_10709_)
);

NAND2X1 _20686_ (
    .A(_10708_),
    .B(_10709_),
    .Y(_10710_)
);

OAI21X1 _20687_ (
    .A(_549__bF$buf4),
    .B(_5668__bF$buf3),
    .C(_10365_),
    .Y(_10711_)
);

NAND3X1 _20688_ (
    .A(_10707_),
    .B(_10711_),
    .C(_10710_),
    .Y(_10712_)
);

NAND2X1 _20689_ (
    .A(areg_13_bF$buf0),
    .B(breg_27_bF$buf5),
    .Y(_10713_)
);

NOR2X1 _20690_ (
    .A(_10365_),
    .B(_10713_),
    .Y(_10714_)
);

NOR2X1 _20691_ (
    .A(_10708_),
    .B(_10709_),
    .Y(_10716_)
);

OAI21X1 _20692_ (
    .A(_10716_),
    .B(_10714_),
    .C(_10706_),
    .Y(_10717_)
);

AOI21X1 _20693_ (
    .A(_10712_),
    .B(_10717_),
    .C(_10705_),
    .Y(_10718_)
);

AOI21X1 _20694_ (
    .A(_10358_),
    .B(_10362_),
    .C(_10366_),
    .Y(_10719_)
);

OAI21X1 _20695_ (
    .A(_10869__bF$buf3),
    .B(_6050__bF$buf1),
    .C(_10709_),
    .Y(_10720_)
);

OAI21X1 _20696_ (
    .A(_549__bF$buf3),
    .B(_5668__bF$buf2),
    .C(_10708_),
    .Y(_10721_)
);

AOI21X1 _20697_ (
    .A(_10720_),
    .B(_10721_),
    .C(_10706_),
    .Y(_10722_)
);

AOI21X1 _20698_ (
    .A(_10711_),
    .B(_10710_),
    .C(_10707_),
    .Y(_10723_)
);

NOR3X1 _20699_ (
    .A(_10723_),
    .B(_10719_),
    .C(_10722_),
    .Y(_10724_)
);

OAI21X1 _20700_ (
    .A(_10724_),
    .B(_10718_),
    .C(_10703_),
    .Y(_10725_)
);

OAI21X1 _20701_ (
    .A(_10722_),
    .B(_10723_),
    .C(_10719_),
    .Y(_10727_)
);

NAND3X1 _20702_ (
    .A(_10712_),
    .B(_10705_),
    .C(_10717_),
    .Y(_10728_)
);

NAND3X1 _20703_ (
    .A(_10702_),
    .B(_10727_),
    .C(_10728_),
    .Y(_10729_)
);

AOI21X1 _20704_ (
    .A(_10729_),
    .B(_10725_),
    .C(_10701_),
    .Y(_10730_)
);

AOI21X1 _20705_ (
    .A(_10354_),
    .B(_10378_),
    .C(_10376_),
    .Y(_10731_)
);

AOI21X1 _20706_ (
    .A(_10727_),
    .B(_10728_),
    .C(_10702_),
    .Y(_10732_)
);

NOR3X1 _20707_ (
    .A(_10718_),
    .B(_10703_),
    .C(_10724_),
    .Y(_10733_)
);

NOR3X1 _20708_ (
    .A(_10731_),
    .B(_10732_),
    .C(_10733_),
    .Y(_10734_)
);

OAI21X1 _20709_ (
    .A(_10734_),
    .B(_10730_),
    .C(_10700_),
    .Y(_10735_)
);

OAI21X1 _20710_ (
    .A(_10733_),
    .B(_10732_),
    .C(_10731_),
    .Y(_10736_)
);

NAND3X1 _20711_ (
    .A(_10701_),
    .B(_10729_),
    .C(_10725_),
    .Y(_10738_)
);

NAND3X1 _20712_ (
    .A(_10699_),
    .B(_10738_),
    .C(_10736_),
    .Y(_10739_)
);

AND2X2 _20713_ (
    .A(_10735_),
    .B(_10739_),
    .Y(_10740_)
);

OAI21X1 _20714_ (
    .A(_10431_),
    .B(_10433_),
    .C(_10424_),
    .Y(_10741_)
);

NAND2X1 _20715_ (
    .A(_10410_),
    .B(_10417_),
    .Y(_10742_)
);

OAI21X1 _20716_ (
    .A(_10400_),
    .B(_10395_),
    .C(_10403_),
    .Y(_10743_)
);

NAND2X1 _20717_ (
    .A(areg_14_bF$buf0),
    .B(breg_26_bF$buf0),
    .Y(_10744_)
);

NAND2X1 _20718_ (
    .A(areg_15_bF$buf3),
    .B(breg_25_bF$buf3),
    .Y(_10745_)
);

NAND2X1 _20719_ (
    .A(areg_16_bF$buf1),
    .B(breg_24_bF$buf4),
    .Y(_10746_)
);

NOR2X1 _20720_ (
    .A(_10745_),
    .B(_10746_),
    .Y(_10747_)
);

AND2X2 _20721_ (
    .A(_10745_),
    .B(_10746_),
    .Y(_10749_)
);

OAI21X1 _20722_ (
    .A(_10749_),
    .B(_10747_),
    .C(_10744_),
    .Y(_10750_)
);

INVX1 _20723_ (
    .A(_10744_),
    .Y(_10751_)
);

OR2X2 _20724_ (
    .A(_10745_),
    .B(_10746_),
    .Y(_10752_)
);

OAI21X1 _20725_ (
    .A(_2669__bF$buf0),
    .B(_5315__bF$buf3),
    .C(_10745_),
    .Y(_10753_)
);

NAND3X1 _20726_ (
    .A(_10751_),
    .B(_10753_),
    .C(_10752_),
    .Y(_10754_)
);

NAND2X1 _20727_ (
    .A(areg_18_bF$buf1),
    .B(breg_22_bF$buf1),
    .Y(_10755_)
);

AND2X2 _20728_ (
    .A(_10406_),
    .B(_10466_),
    .Y(_10756_)
);

OAI22X1 _20729_ (
    .A(_10114_),
    .B(_10755_),
    .C(_10756_),
    .D(_10464_),
    .Y(_10757_)
);

NAND3X1 _20730_ (
    .A(_10750_),
    .B(_10754_),
    .C(_10757_),
    .Y(_10758_)
);

AOI21X1 _20731_ (
    .A(_10753_),
    .B(_10752_),
    .C(_10751_),
    .Y(_10760_)
);

NOR3X1 _20732_ (
    .A(_10744_),
    .B(_10747_),
    .C(_10749_),
    .Y(_10761_)
);

NOR2X1 _20733_ (
    .A(_10406_),
    .B(_10466_),
    .Y(_10762_)
);

OAI21X1 _20734_ (
    .A(_3146__bF$buf0),
    .B(_3781__bF$buf3),
    .C(_10406_),
    .Y(_10763_)
);

AOI21X1 _20735_ (
    .A(_10465_),
    .B(_10763_),
    .C(_10762_),
    .Y(_10764_)
);

OAI21X1 _20736_ (
    .A(_10761_),
    .B(_10760_),
    .C(_10764_),
    .Y(_10765_)
);

NAND3X1 _20737_ (
    .A(_10743_),
    .B(_10758_),
    .C(_10765_),
    .Y(_10766_)
);

INVX1 _20738_ (
    .A(_10743_),
    .Y(_10767_)
);

NAND3X1 _20739_ (
    .A(_10764_),
    .B(_10750_),
    .C(_10754_),
    .Y(_10768_)
);

OAI21X1 _20740_ (
    .A(_10761_),
    .B(_10760_),
    .C(_10757_),
    .Y(_10769_)
);

NAND3X1 _20741_ (
    .A(_10767_),
    .B(_10768_),
    .C(_10769_),
    .Y(_10771_)
);

AOI21X1 _20742_ (
    .A(_10483_),
    .B(_10488_),
    .C(_10469_),
    .Y(_10772_)
);

OAI21X1 _20743_ (
    .A(_10468_),
    .B(_10772_),
    .C(_10492_),
    .Y(_10773_)
);

NAND3X1 _20744_ (
    .A(_10766_),
    .B(_10771_),
    .C(_10773_),
    .Y(_10774_)
);

AOI21X1 _20745_ (
    .A(_10768_),
    .B(_10769_),
    .C(_10767_),
    .Y(_10775_)
);

AOI21X1 _20746_ (
    .A(_10758_),
    .B(_10765_),
    .C(_10743_),
    .Y(_10776_)
);

NOR3X1 _20747_ (
    .A(_10480_),
    .B(_10482_),
    .C(_10476_),
    .Y(_10777_)
);

AOI21X1 _20748_ (
    .A(_10493_),
    .B(_10491_),
    .C(_10777_),
    .Y(_10778_)
);

OAI21X1 _20749_ (
    .A(_10775_),
    .B(_10776_),
    .C(_10778_),
    .Y(_10779_)
);

NAND3X1 _20750_ (
    .A(_10742_),
    .B(_10779_),
    .C(_10774_),
    .Y(_10780_)
);

INVX2 _20751_ (
    .A(_10742_),
    .Y(_10782_)
);

NOR3X1 _20752_ (
    .A(_10775_),
    .B(_10776_),
    .C(_10778_),
    .Y(_10783_)
);

AOI21X1 _20753_ (
    .A(_10766_),
    .B(_10771_),
    .C(_10773_),
    .Y(_10784_)
);

OAI21X1 _20754_ (
    .A(_10783_),
    .B(_10784_),
    .C(_10782_),
    .Y(_10785_)
);

NAND3X1 _20755_ (
    .A(_10780_),
    .B(_10785_),
    .C(_10741_),
    .Y(_10786_)
);

AOI21X1 _20756_ (
    .A(_10393_),
    .B(_10428_),
    .C(_10432_),
    .Y(_10787_)
);

NAND3X1 _20757_ (
    .A(_10766_),
    .B(_10771_),
    .C(_10778_),
    .Y(_10788_)
);

OAI21X1 _20758_ (
    .A(_10775_),
    .B(_10776_),
    .C(_10773_),
    .Y(_10789_)
);

AOI21X1 _20759_ (
    .A(_10789_),
    .B(_10788_),
    .C(_10782_),
    .Y(_10790_)
);

AOI21X1 _20760_ (
    .A(_10779_),
    .B(_10774_),
    .C(_10742_),
    .Y(_10791_)
);

OAI21X1 _20761_ (
    .A(_10790_),
    .B(_10791_),
    .C(_10787_),
    .Y(_10793_)
);

NAND3X1 _20762_ (
    .A(_10786_),
    .B(_10793_),
    .C(_10740_),
    .Y(_10794_)
);

NAND2X1 _20763_ (
    .A(_10739_),
    .B(_10735_),
    .Y(_10795_)
);

OAI21X1 _20764_ (
    .A(_10790_),
    .B(_10791_),
    .C(_10741_),
    .Y(_10796_)
);

NAND3X1 _20765_ (
    .A(_10787_),
    .B(_10780_),
    .C(_10785_),
    .Y(_10797_)
);

NAND3X1 _20766_ (
    .A(_10795_),
    .B(_10796_),
    .C(_10797_),
    .Y(_10798_)
);

OAI21X1 _20767_ (
    .A(_10553_),
    .B(_10550_),
    .C(_10543_),
    .Y(_10799_)
);

NAND3X1 _20768_ (
    .A(_10798_),
    .B(_10799_),
    .C(_10794_),
    .Y(_10800_)
);

AOI21X1 _20769_ (
    .A(_10796_),
    .B(_10797_),
    .C(_10795_),
    .Y(_10801_)
);

AOI21X1 _20770_ (
    .A(_10786_),
    .B(_10793_),
    .C(_10740_),
    .Y(_10802_)
);

AOI21X1 _20771_ (
    .A(_10462_),
    .B(_10548_),
    .C(_10552_),
    .Y(_10804_)
);

OAI21X1 _20772_ (
    .A(_10802_),
    .B(_10801_),
    .C(_10804_),
    .Y(_10805_)
);

NAND3X1 _20773_ (
    .A(_10698_),
    .B(_10800_),
    .C(_10805_),
    .Y(_10806_)
);

AND2X2 _20774_ (
    .A(_10443_),
    .B(_10435_),
    .Y(_10807_)
);

NAND3X1 _20775_ (
    .A(_10798_),
    .B(_10804_),
    .C(_10794_),
    .Y(_10808_)
);

OAI21X1 _20776_ (
    .A(_10802_),
    .B(_10801_),
    .C(_10799_),
    .Y(_10809_)
);

NAND3X1 _20777_ (
    .A(_10808_),
    .B(_10809_),
    .C(_10807_),
    .Y(_10810_)
);

NAND2X1 _20778_ (
    .A(_10806_),
    .B(_10810_),
    .Y(_10811_)
);

INVX1 _20779_ (
    .A(_10602_),
    .Y(_10812_)
);

OAI21X1 _20780_ (
    .A(_10555_),
    .B(_10812_),
    .C(_10607_),
    .Y(_10813_)
);

NAND2X1 _20781_ (
    .A(_10527_),
    .B(_10535_),
    .Y(_10815_)
);

NAND2X1 _20782_ (
    .A(areg_17_bF$buf1),
    .B(breg_23_bF$buf2),
    .Y(_10816_)
);

INVX2 _20783_ (
    .A(_10816_),
    .Y(_10817_)
);

NAND2X1 _20784_ (
    .A(areg_19_bF$buf3),
    .B(breg_21_bF$buf1),
    .Y(_10818_)
);

XOR2X1 _20785_ (
    .A(_10755_),
    .B(_10818_),
    .Y(_10819_)
);

XNOR2X1 _20786_ (
    .A(_10819_),
    .B(_10817_),
    .Y(_10820_)
);

OAI21X1 _20787_ (
    .A(_10487_),
    .B(_10470_),
    .C(_10478_),
    .Y(_10821_)
);

NAND2X1 _20788_ (
    .A(areg_20_bF$buf3),
    .B(breg_20_bF$buf2),
    .Y(_10822_)
);

AND2X2 _20789_ (
    .A(breg_18_bF$buf5),
    .B(areg_22_bF$buf1),
    .Y(_10823_)
);

OAI21X1 _20790_ (
    .A(_3253__bF$buf2),
    .B(_3961__bF$buf2),
    .C(_10823_),
    .Y(_10824_)
);

AND2X2 _20791_ (
    .A(breg_19_bF$buf0),
    .B(areg_21_bF$buf1),
    .Y(_10826_)
);

OAI21X1 _20792_ (
    .A(_3529__bF$buf0),
    .B(_4551__bF$buf2),
    .C(_10826_),
    .Y(_10827_)
);

AOI21X1 _20793_ (
    .A(_10824_),
    .B(_10827_),
    .C(_10822_),
    .Y(_10828_)
);

INVX2 _20794_ (
    .A(_10822_),
    .Y(_10829_)
);

NAND2X1 _20795_ (
    .A(_10826_),
    .B(_10823_),
    .Y(_10830_)
);

NAND2X1 _20796_ (
    .A(breg_19_bF$buf5),
    .B(areg_21_bF$buf0),
    .Y(_10831_)
);

OAI21X1 _20797_ (
    .A(_3529__bF$buf4),
    .B(_4551__bF$buf1),
    .C(_10831_),
    .Y(_10832_)
);

AOI21X1 _20798_ (
    .A(_10832_),
    .B(_10830_),
    .C(_10829_),
    .Y(_10833_)
);

OAI21X1 _20799_ (
    .A(_10828_),
    .B(_10833_),
    .C(_10821_),
    .Y(_10834_)
);

AOI21X1 _20800_ (
    .A(_10477_),
    .B(_10479_),
    .C(_10486_),
    .Y(_10835_)
);

NAND3X1 _20801_ (
    .A(_10829_),
    .B(_10832_),
    .C(_10830_),
    .Y(_10837_)
);

NAND2X1 _20802_ (
    .A(breg_18_bF$buf4),
    .B(areg_22_bF$buf0),
    .Y(_10838_)
);

NOR2X1 _20803_ (
    .A(_10831_),
    .B(_10838_),
    .Y(_10839_)
);

NOR2X1 _20804_ (
    .A(_10826_),
    .B(_10823_),
    .Y(_10840_)
);

OAI21X1 _20805_ (
    .A(_10840_),
    .B(_10839_),
    .C(_10822_),
    .Y(_10841_)
);

NAND3X1 _20806_ (
    .A(_10835_),
    .B(_10837_),
    .C(_10841_),
    .Y(_10842_)
);

AOI21X1 _20807_ (
    .A(_10834_),
    .B(_10842_),
    .C(_10820_),
    .Y(_10843_)
);

XNOR2X1 _20808_ (
    .A(_10819_),
    .B(_10816_),
    .Y(_10844_)
);

NAND3X1 _20809_ (
    .A(_10837_),
    .B(_10821_),
    .C(_10841_),
    .Y(_10845_)
);

OAI21X1 _20810_ (
    .A(_10828_),
    .B(_10833_),
    .C(_10835_),
    .Y(_10846_)
);

AOI21X1 _20811_ (
    .A(_10846_),
    .B(_10845_),
    .C(_10844_),
    .Y(_10848_)
);

NOR2X1 _20812_ (
    .A(_10843_),
    .B(_10848_),
    .Y(_10849_)
);

OAI21X1 _20813_ (
    .A(_10525_),
    .B(_10523_),
    .C(_10514_),
    .Y(_10850_)
);

NAND2X1 _20814_ (
    .A(breg_16_bF$buf0),
    .B(areg_24_bF$buf3),
    .Y(_10851_)
);

OAI21X1 _20815_ (
    .A(_10498_),
    .B(_10851_),
    .C(_10506_),
    .Y(_10852_)
);

NAND2X1 _20816_ (
    .A(breg_17_bF$buf0),
    .B(areg_23_bF$buf4),
    .Y(_10853_)
);

INVX1 _20817_ (
    .A(_10853_),
    .Y(_10854_)
);

AND2X2 _20818_ (
    .A(breg_16_bF$buf5),
    .B(areg_24_bF$buf2),
    .Y(_10855_)
);

AND2X2 _20819_ (
    .A(breg_15_bF$buf2),
    .B(areg_25_bF$buf0),
    .Y(_10856_)
);

NAND2X1 _20820_ (
    .A(_10855_),
    .B(_10856_),
    .Y(_10857_)
);

OAI21X1 _20821_ (
    .A(_2362__bF$buf0),
    .B(_6300__bF$buf2),
    .C(_10851_),
    .Y(_10859_)
);

NAND3X1 _20822_ (
    .A(_10854_),
    .B(_10859_),
    .C(_10857_),
    .Y(_10860_)
);

NAND2X1 _20823_ (
    .A(breg_15_bF$buf1),
    .B(areg_25_bF$buf4),
    .Y(_10861_)
);

NOR2X1 _20824_ (
    .A(_10851_),
    .B(_10861_),
    .Y(_10862_)
);

NOR2X1 _20825_ (
    .A(_10855_),
    .B(_10856_),
    .Y(_10863_)
);

OAI21X1 _20826_ (
    .A(_10863_),
    .B(_10862_),
    .C(_10853_),
    .Y(_10864_)
);

NAND2X1 _20827_ (
    .A(breg_13_bF$buf2),
    .B(areg_27_bF$buf3),
    .Y(_10865_)
);

AND2X2 _20828_ (
    .A(_10511_),
    .B(_10558_),
    .Y(_10866_)
);

OAI22X1 _20829_ (
    .A(_10212_),
    .B(_10865_),
    .C(_10866_),
    .D(_10557_),
    .Y(_10867_)
);

NAND3X1 _20830_ (
    .A(_10860_),
    .B(_10867_),
    .C(_10864_),
    .Y(_10868_)
);

NOR3X1 _20831_ (
    .A(_10853_),
    .B(_10862_),
    .C(_10863_),
    .Y(_10870_)
);

AOI21X1 _20832_ (
    .A(_10859_),
    .B(_10857_),
    .C(_10854_),
    .Y(_10871_)
);

NOR2X1 _20833_ (
    .A(_10511_),
    .B(_10558_),
    .Y(_10872_)
);

OAI21X1 _20834_ (
    .A(_2586__bF$buf1),
    .B(_7100__bF$buf3),
    .C(_10511_),
    .Y(_10873_)
);

AOI21X1 _20835_ (
    .A(_10580_),
    .B(_10873_),
    .C(_10872_),
    .Y(_10874_)
);

OAI21X1 _20836_ (
    .A(_10870_),
    .B(_10871_),
    .C(_10874_),
    .Y(_10875_)
);

NAND3X1 _20837_ (
    .A(_10852_),
    .B(_10868_),
    .C(_10875_),
    .Y(_10876_)
);

AOI21X1 _20838_ (
    .A(_10149_),
    .B(_10855_),
    .C(_10515_),
    .Y(_10877_)
);

NOR3X1 _20839_ (
    .A(_10871_),
    .B(_10874_),
    .C(_10870_),
    .Y(_10878_)
);

AOI21X1 _20840_ (
    .A(_10860_),
    .B(_10864_),
    .C(_10867_),
    .Y(_10879_)
);

OAI21X1 _20841_ (
    .A(_10878_),
    .B(_10879_),
    .C(_10877_),
    .Y(_10881_)
);

NAND3X1 _20842_ (
    .A(_10850_),
    .B(_10876_),
    .C(_10881_),
    .Y(_10882_)
);

AOI21X1 _20843_ (
    .A(_10499_),
    .B(_10521_),
    .C(_10524_),
    .Y(_10883_)
);

NAND3X1 _20844_ (
    .A(_10860_),
    .B(_10874_),
    .C(_10864_),
    .Y(_10884_)
);

OAI21X1 _20845_ (
    .A(_10870_),
    .B(_10871_),
    .C(_10867_),
    .Y(_10885_)
);

AOI21X1 _20846_ (
    .A(_10884_),
    .B(_10885_),
    .C(_10877_),
    .Y(_10886_)
);

AOI21X1 _20847_ (
    .A(_10868_),
    .B(_10875_),
    .C(_10852_),
    .Y(_10887_)
);

OAI21X1 _20848_ (
    .A(_10887_),
    .B(_10886_),
    .C(_10883_),
    .Y(_10888_)
);

NAND3X1 _20849_ (
    .A(_10849_),
    .B(_10888_),
    .C(_10882_),
    .Y(_10889_)
);

OR2X2 _20850_ (
    .A(_10843_),
    .B(_10848_),
    .Y(_10890_)
);

OAI21X1 _20851_ (
    .A(_10887_),
    .B(_10886_),
    .C(_10850_),
    .Y(_10892_)
);

NAND3X1 _20852_ (
    .A(_10883_),
    .B(_10876_),
    .C(_10881_),
    .Y(_10893_)
);

NAND3X1 _20853_ (
    .A(_10890_),
    .B(_10892_),
    .C(_10893_),
    .Y(_10894_)
);

AOI21X1 _20854_ (
    .A(_10579_),
    .B(_10585_),
    .C(_10263_),
    .Y(_10895_)
);

OAI21X1 _20855_ (
    .A(_10895_),
    .B(_10591_),
    .C(_10586_),
    .Y(_10896_)
);

NAND3X1 _20856_ (
    .A(_10896_),
    .B(_10889_),
    .C(_10894_),
    .Y(_10897_)
);

AOI21X1 _20857_ (
    .A(_10892_),
    .B(_10893_),
    .C(_10890_),
    .Y(_10898_)
);

AOI21X1 _20858_ (
    .A(_10888_),
    .B(_10882_),
    .C(_10849_),
    .Y(_10899_)
);

NOR3X1 _20859_ (
    .A(_10588_),
    .B(_10262_),
    .C(_10587_),
    .Y(_10900_)
);

AOI21X1 _20860_ (
    .A(_10556_),
    .B(_10589_),
    .C(_10900_),
    .Y(_10901_)
);

OAI21X1 _20861_ (
    .A(_10898_),
    .B(_10899_),
    .C(_10901_),
    .Y(_10903_)
);

NAND3X1 _20862_ (
    .A(_10815_),
    .B(_10897_),
    .C(_10903_),
    .Y(_10904_)
);

AND2X2 _20863_ (
    .A(_10535_),
    .B(_10527_),
    .Y(_10905_)
);

NAND3X1 _20864_ (
    .A(_10889_),
    .B(_10894_),
    .C(_10901_),
    .Y(_10906_)
);

OAI21X1 _20865_ (
    .A(_10898_),
    .B(_10899_),
    .C(_10896_),
    .Y(_10907_)
);

NAND3X1 _20866_ (
    .A(_10905_),
    .B(_10906_),
    .C(_10907_),
    .Y(_10908_)
);

NAND2X1 _20867_ (
    .A(_10904_),
    .B(_10908_),
    .Y(_10909_)
);

NAND2X1 _20868_ (
    .A(_10574_),
    .B(_10579_),
    .Y(_10910_)
);

NAND2X1 _20869_ (
    .A(breg_14_bF$buf3),
    .B(areg_26_bF$buf0),
    .Y(_10911_)
);

NAND2X1 _20870_ (
    .A(breg_12_bF$buf0),
    .B(areg_28_bF$buf4),
    .Y(_10912_)
);

XOR2X1 _20871_ (
    .A(_10865_),
    .B(_10912_),
    .Y(_10914_)
);

XNOR2X1 _20872_ (
    .A(_10914_),
    .B(_10911_),
    .Y(_10915_)
);

OAI21X1 _20873_ (
    .A(_10567_),
    .B(_10563_),
    .C(_10566_),
    .Y(_10916_)
);

NAND2X1 _20874_ (
    .A(breg_11_bF$buf2),
    .B(areg_29_bF$buf1),
    .Y(_10917_)
);

INVX1 _20875_ (
    .A(_10917_),
    .Y(_10918_)
);

AND2X2 _20876_ (
    .A(breg_9_bF$buf2),
    .B(areg_31_bF$buf0),
    .Y(_10919_)
);

NAND2X1 _20877_ (
    .A(_10565_),
    .B(_10919_),
    .Y(_10920_)
);

OAI21X1 _20878_ (
    .A(_6044__bF$buf0),
    .B(_8773_),
    .C(_10570_),
    .Y(_10921_)
);

NAND3X1 _20879_ (
    .A(_10918_),
    .B(_10921_),
    .C(_10920_),
    .Y(_10922_)
);

OAI21X1 _20880_ (
    .A(_7217__bF$buf4),
    .B(_8759_),
    .C(_10919_),
    .Y(_10923_)
);

OAI21X1 _20881_ (
    .A(_6044__bF$buf5),
    .B(_8773_),
    .C(_10565_),
    .Y(_10925_)
);

NAND3X1 _20882_ (
    .A(_10917_),
    .B(_10923_),
    .C(_10925_),
    .Y(_10926_)
);

NAND3X1 _20883_ (
    .A(_10916_),
    .B(_10922_),
    .C(_10926_),
    .Y(_10927_)
);

AOI21X1 _20884_ (
    .A(_10564_),
    .B(_10568_),
    .C(_10571_),
    .Y(_10928_)
);

AOI21X1 _20885_ (
    .A(_10923_),
    .B(_10925_),
    .C(_10917_),
    .Y(_10929_)
);

AOI21X1 _20886_ (
    .A(_10921_),
    .B(_10920_),
    .C(_10918_),
    .Y(_10930_)
);

OAI21X1 _20887_ (
    .A(_10929_),
    .B(_10930_),
    .C(_10928_),
    .Y(_10931_)
);

NAND3X1 _20888_ (
    .A(_10927_),
    .B(_10931_),
    .C(_10915_),
    .Y(_10932_)
);

INVX2 _20889_ (
    .A(_10911_),
    .Y(_10933_)
);

XNOR2X1 _20890_ (
    .A(_10914_),
    .B(_10933_),
    .Y(_10934_)
);

OAI21X1 _20891_ (
    .A(_10929_),
    .B(_10930_),
    .C(_10916_),
    .Y(_10936_)
);

NAND3X1 _20892_ (
    .A(_10928_),
    .B(_10922_),
    .C(_10926_),
    .Y(_10937_)
);

NAND3X1 _20893_ (
    .A(_10936_),
    .B(_10937_),
    .C(_10934_),
    .Y(_10938_)
);

NAND3X1 _20894_ (
    .A(_10258_),
    .B(_10932_),
    .C(_10938_),
    .Y(_10939_)
);

INVX2 _20895_ (
    .A(_10258_),
    .Y(_10940_)
);

AOI21X1 _20896_ (
    .A(_10936_),
    .B(_10937_),
    .C(_10934_),
    .Y(_10941_)
);

AOI21X1 _20897_ (
    .A(_10927_),
    .B(_10931_),
    .C(_10915_),
    .Y(_10942_)
);

OAI21X1 _20898_ (
    .A(_10941_),
    .B(_10942_),
    .C(_10940_),
    .Y(_10943_)
);

NAND3X1 _20899_ (
    .A(_10910_),
    .B(_10939_),
    .C(_10943_),
    .Y(_10944_)
);

AND2X2 _20900_ (
    .A(_10579_),
    .B(_10574_),
    .Y(_10945_)
);

NAND3X1 _20901_ (
    .A(_10940_),
    .B(_10932_),
    .C(_10938_),
    .Y(_10947_)
);

OAI21X1 _20902_ (
    .A(_10941_),
    .B(_10942_),
    .C(_10258_),
    .Y(_10948_)
);

NAND3X1 _20903_ (
    .A(_10947_),
    .B(_10945_),
    .C(_10948_),
    .Y(_10949_)
);

NAND2X1 _20904_ (
    .A(_10944_),
    .B(_10949_),
    .Y(_10950_)
);

XNOR2X1 _20905_ (
    .A(_10605_),
    .B(_10950_),
    .Y(_10951_)
);

NOR2X1 _20906_ (
    .A(_10951_),
    .B(_10909_),
    .Y(_10952_)
);

AOI21X1 _20907_ (
    .A(_10906_),
    .B(_10907_),
    .C(_10905_),
    .Y(_10953_)
);

AOI21X1 _20908_ (
    .A(_10897_),
    .B(_10903_),
    .C(_10815_),
    .Y(_10954_)
);

OAI21X1 _20909_ (
    .A(_10953_),
    .B(_10954_),
    .C(_10951_),
    .Y(_10955_)
);

INVX1 _20910_ (
    .A(_10955_),
    .Y(_10956_)
);

OAI21X1 _20911_ (
    .A(_10956_),
    .B(_10952_),
    .C(_10813_),
    .Y(_10958_)
);

INVX1 _20912_ (
    .A(_10607_),
    .Y(_10959_)
);

AOI21X1 _20913_ (
    .A(_10602_),
    .B(_10614_),
    .C(_10959_),
    .Y(_10960_)
);

XOR2X1 _20914_ (
    .A(_10605_),
    .B(_10950_),
    .Y(_10961_)
);

NAND3X1 _20915_ (
    .A(_10904_),
    .B(_10908_),
    .C(_10961_),
    .Y(_10962_)
);

NAND3X1 _20916_ (
    .A(_10962_),
    .B(_10955_),
    .C(_10960_),
    .Y(_10963_)
);

AOI21X1 _20917_ (
    .A(_10963_),
    .B(_10958_),
    .C(_10811_),
    .Y(_10964_)
);

NAND3X1 _20918_ (
    .A(_10800_),
    .B(_10805_),
    .C(_10807_),
    .Y(_10965_)
);

NAND3X1 _20919_ (
    .A(_10698_),
    .B(_10808_),
    .C(_10809_),
    .Y(_10966_)
);

NAND2X1 _20920_ (
    .A(_10966_),
    .B(_10965_),
    .Y(_10967_)
);

NAND3X1 _20921_ (
    .A(_10962_),
    .B(_10955_),
    .C(_10813_),
    .Y(_10969_)
);

OAI21X1 _20922_ (
    .A(_10956_),
    .B(_10952_),
    .C(_10960_),
    .Y(_10970_)
);

AOI21X1 _20923_ (
    .A(_10969_),
    .B(_10970_),
    .C(_10967_),
    .Y(_10971_)
);

OAI21X1 _20924_ (
    .A(_10964_),
    .B(_10971_),
    .C(_10697_),
    .Y(_10972_)
);

NOR3X1 _20925_ (
    .A(_10609_),
    .B(_10615_),
    .C(_10618_),
    .Y(_10973_)
);

AOI21X1 _20926_ (
    .A(_10625_),
    .B(_10627_),
    .C(_10973_),
    .Y(_10974_)
);

NAND3X1 _20927_ (
    .A(_10969_),
    .B(_10967_),
    .C(_10970_),
    .Y(_10975_)
);

NAND3X1 _20928_ (
    .A(_10963_),
    .B(_10811_),
    .C(_10958_),
    .Y(_10976_)
);

NAND3X1 _20929_ (
    .A(_10975_),
    .B(_10976_),
    .C(_10974_),
    .Y(_10977_)
);

AOI21X1 _20930_ (
    .A(_10977_),
    .B(_10972_),
    .C(_10695_),
    .Y(_10978_)
);

NAND3X1 _20931_ (
    .A(_10976_),
    .B(_10975_),
    .C(_10697_),
    .Y(_10980_)
);

OAI21X1 _20932_ (
    .A(_10964_),
    .B(_10971_),
    .C(_10974_),
    .Y(_10981_)
);

AOI21X1 _20933_ (
    .A(_10980_),
    .B(_10981_),
    .C(_10694_),
    .Y(_10982_)
);

OAI21X1 _20934_ (
    .A(_10982_),
    .B(_10978_),
    .C(_10692_),
    .Y(_10983_)
);

AOI21X1 _20935_ (
    .A(_10638_),
    .B(_10345_),
    .C(_10645_),
    .Y(_10984_)
);

NAND3X1 _20936_ (
    .A(_10694_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10985_)
);

NAND3X1 _20937_ (
    .A(_10695_),
    .B(_10977_),
    .C(_10972_),
    .Y(_10986_)
);

NAND3X1 _20938_ (
    .A(_10986_),
    .B(_10985_),
    .C(_10984_),
    .Y(_10987_)
);

AOI21X1 _20939_ (
    .A(_10987_),
    .B(_10983_),
    .C(_10691_),
    .Y(_10988_)
);

NAND3X1 _20940_ (
    .A(_10985_),
    .B(_10692_),
    .C(_10986_),
    .Y(_10989_)
);

OAI21X1 _20941_ (
    .A(_10982_),
    .B(_10978_),
    .C(_10984_),
    .Y(_10991_)
);

AOI21X1 _20942_ (
    .A(_10989_),
    .B(_10991_),
    .C(_10690_),
    .Y(_10992_)
);

OAI22X1 _20943_ (
    .A(_10988_),
    .B(_10992_),
    .C(_10649_),
    .D(_10689_),
    .Y(_10993_)
);

AOI21X1 _20944_ (
    .A(_10340_),
    .B(_10652_),
    .C(_10689_),
    .Y(_10994_)
);

NAND3X1 _20945_ (
    .A(_10690_),
    .B(_10989_),
    .C(_10991_),
    .Y(_10995_)
);

NAND3X1 _20946_ (
    .A(_10691_),
    .B(_10987_),
    .C(_10983_),
    .Y(_10996_)
);

NAND3X1 _20947_ (
    .A(_10995_),
    .B(_10996_),
    .C(_10994_),
    .Y(_10997_)
);

NAND2X1 _20948_ (
    .A(_10997_),
    .B(_10993_),
    .Y(_10998_)
);

INVX1 _20949_ (
    .A(_10998_),
    .Y(_10999_)
);

XNOR2X1 _20950_ (
    .A(_10688_),
    .B(_10999_),
    .Y(_0_[40])
);

NAND2X1 _20951_ (
    .A(_10995_),
    .B(_10996_),
    .Y(_11001_)
);

NOR2X1 _20952_ (
    .A(_10994_),
    .B(_11001_),
    .Y(_11002_)
);

AOI21X1 _20953_ (
    .A(_10998_),
    .B(_10688_),
    .C(_11002_),
    .Y(_11003_)
);

AOI21X1 _20954_ (
    .A(_10985_),
    .B(_10986_),
    .C(_10692_),
    .Y(_11004_)
);

OAI21X1 _20955_ (
    .A(_11004_),
    .B(_10691_),
    .C(_10989_),
    .Y(_11005_)
);

OAI21X1 _20956_ (
    .A(_10730_),
    .B(_10700_),
    .C(_10738_),
    .Y(_11006_)
);

INVX2 _20957_ (
    .A(_11006_),
    .Y(_11007_)
);

AOI21X1 _20958_ (
    .A(_10976_),
    .B(_10975_),
    .C(_10697_),
    .Y(_11008_)
);

OAI21X1 _20959_ (
    .A(_11008_),
    .B(_10695_),
    .C(_10980_),
    .Y(_11009_)
);

NAND2X1 _20960_ (
    .A(_10800_),
    .B(_10806_),
    .Y(_11010_)
);

INVX2 _20961_ (
    .A(_11010_),
    .Y(_11012_)
);

AOI21X1 _20962_ (
    .A(_10962_),
    .B(_10955_),
    .C(_10813_),
    .Y(_11013_)
);

OAI21X1 _20963_ (
    .A(_10811_),
    .B(_11013_),
    .C(_10969_),
    .Y(_11014_)
);

NAND2X1 _20964_ (
    .A(_10786_),
    .B(_10794_),
    .Y(_11015_)
);

NOR2X1 _20965_ (
    .A(_7711__bF$buf3),
    .B(_7225__bF$buf4),
    .Y(_11016_)
);

INVX1 _20966_ (
    .A(_11016_),
    .Y(_11017_)
);

OAI21X1 _20967_ (
    .A(_10718_),
    .B(_10703_),
    .C(_10728_),
    .Y(_11018_)
);

NOR2X1 _20968_ (
    .A(_9104__bF$buf1),
    .B(_6815__bF$buf3),
    .Y(_11019_)
);

INVX2 _20969_ (
    .A(_11019_),
    .Y(_11020_)
);

OAI21X1 _20970_ (
    .A(_10716_),
    .B(_10706_),
    .C(_10710_),
    .Y(_11021_)
);

NAND2X1 _20971_ (
    .A(areg_12_bF$buf1),
    .B(breg_29_bF$buf2),
    .Y(_11023_)
);

INVX2 _20972_ (
    .A(_11023_),
    .Y(_11024_)
);

AND2X2 _20973_ (
    .A(areg_13_bF$buf4),
    .B(breg_28_bF$buf4),
    .Y(_11025_)
);

AND2X2 _20974_ (
    .A(areg_14_bF$buf4),
    .B(breg_27_bF$buf4),
    .Y(_11026_)
);

NAND2X1 _20975_ (
    .A(_11025_),
    .B(_11026_),
    .Y(_11027_)
);

OAI22X1 _20976_ (
    .A(_549__bF$buf2),
    .B(_6050__bF$buf0),
    .C(_2287__bF$buf2),
    .D(_5668__bF$buf1),
    .Y(_11028_)
);

NAND3X1 _20977_ (
    .A(_11024_),
    .B(_11028_),
    .C(_11027_),
    .Y(_11029_)
);

NAND2X1 _20978_ (
    .A(areg_14_bF$buf3),
    .B(breg_28_bF$buf3),
    .Y(_11030_)
);

NOR2X1 _20979_ (
    .A(_10713_),
    .B(_11030_),
    .Y(_11031_)
);

NOR2X1 _20980_ (
    .A(_11025_),
    .B(_11026_),
    .Y(_11032_)
);

OAI21X1 _20981_ (
    .A(_11032_),
    .B(_11031_),
    .C(_11023_),
    .Y(_11033_)
);

AOI21X1 _20982_ (
    .A(_11029_),
    .B(_11033_),
    .C(_11021_),
    .Y(_11034_)
);

AOI21X1 _20983_ (
    .A(_10707_),
    .B(_10711_),
    .C(_10714_),
    .Y(_11035_)
);

OAI21X1 _20984_ (
    .A(_549__bF$buf1),
    .B(_6050__bF$buf3),
    .C(_11026_),
    .Y(_11036_)
);

OAI21X1 _20985_ (
    .A(_2287__bF$buf1),
    .B(_5668__bF$buf0),
    .C(_11025_),
    .Y(_11037_)
);

AOI21X1 _20986_ (
    .A(_11036_),
    .B(_11037_),
    .C(_11023_),
    .Y(_11038_)
);

AOI21X1 _20987_ (
    .A(_11028_),
    .B(_11027_),
    .C(_11024_),
    .Y(_11039_)
);

NOR3X1 _20988_ (
    .A(_11039_),
    .B(_11035_),
    .C(_11038_),
    .Y(_11040_)
);

OAI21X1 _20989_ (
    .A(_11040_),
    .B(_11034_),
    .C(_11020_),
    .Y(_11041_)
);

OAI21X1 _20990_ (
    .A(_11038_),
    .B(_11039_),
    .C(_11035_),
    .Y(_11042_)
);

NAND3X1 _20991_ (
    .A(_11029_),
    .B(_11021_),
    .C(_11033_),
    .Y(_11045_)
);

NAND3X1 _20992_ (
    .A(_11019_),
    .B(_11042_),
    .C(_11045_),
    .Y(_11046_)
);

AOI21X1 _20993_ (
    .A(_11046_),
    .B(_11041_),
    .C(_11018_),
    .Y(_11047_)
);

AOI21X1 _20994_ (
    .A(_10702_),
    .B(_10727_),
    .C(_10724_),
    .Y(_11048_)
);

AOI21X1 _20995_ (
    .A(_11042_),
    .B(_11045_),
    .C(_11019_),
    .Y(_11049_)
);

NOR3X1 _20996_ (
    .A(_11034_),
    .B(_11020_),
    .C(_11040_),
    .Y(_11050_)
);

NOR3X1 _20997_ (
    .A(_11048_),
    .B(_11049_),
    .C(_11050_),
    .Y(_11051_)
);

OAI21X1 _20998_ (
    .A(_11051_),
    .B(_11047_),
    .C(_11017_),
    .Y(_11052_)
);

OAI21X1 _20999_ (
    .A(_11050_),
    .B(_11049_),
    .C(_11048_),
    .Y(_11053_)
);

NAND3X1 _21000_ (
    .A(_11018_),
    .B(_11046_),
    .C(_11041_),
    .Y(_11054_)
);

NAND3X1 _21001_ (
    .A(_11016_),
    .B(_11054_),
    .C(_11053_),
    .Y(_11056_)
);

AND2X2 _21002_ (
    .A(_11052_),
    .B(_11056_),
    .Y(_11057_)
);

OAI21X1 _21003_ (
    .A(_10782_),
    .B(_10784_),
    .C(_10774_),
    .Y(_11058_)
);

NAND2X1 _21004_ (
    .A(_10758_),
    .B(_10766_),
    .Y(_11059_)
);

OAI21X1 _21005_ (
    .A(_10749_),
    .B(_10744_),
    .C(_10752_),
    .Y(_11060_)
);

NAND2X1 _21006_ (
    .A(areg_15_bF$buf2),
    .B(breg_26_bF$buf4),
    .Y(_11061_)
);

NAND2X1 _21007_ (
    .A(areg_16_bF$buf0),
    .B(breg_25_bF$buf2),
    .Y(_11062_)
);

NAND2X1 _21008_ (
    .A(areg_17_bF$buf0),
    .B(breg_24_bF$buf3),
    .Y(_11063_)
);

NOR2X1 _21009_ (
    .A(_11062_),
    .B(_11063_),
    .Y(_11064_)
);

AND2X2 _21010_ (
    .A(_11062_),
    .B(_11063_),
    .Y(_11065_)
);

OAI21X1 _21011_ (
    .A(_11065_),
    .B(_11064_),
    .C(_11061_),
    .Y(_11067_)
);

INVX1 _21012_ (
    .A(_11061_),
    .Y(_11068_)
);

OR2X2 _21013_ (
    .A(_11062_),
    .B(_11063_),
    .Y(_11069_)
);

OAI21X1 _21014_ (
    .A(_2884__bF$buf2),
    .B(_5315__bF$buf2),
    .C(_11062_),
    .Y(_11070_)
);

NAND3X1 _21015_ (
    .A(_11068_),
    .B(_11070_),
    .C(_11069_),
    .Y(_11071_)
);

NAND2X1 _21016_ (
    .A(areg_19_bF$buf2),
    .B(breg_22_bF$buf0),
    .Y(_11072_)
);

AND2X2 _21017_ (
    .A(_10755_),
    .B(_10818_),
    .Y(_11073_)
);

OAI22X1 _21018_ (
    .A(_10466_),
    .B(_11072_),
    .C(_11073_),
    .D(_10816_),
    .Y(_11074_)
);

NAND3X1 _21019_ (
    .A(_11067_),
    .B(_11071_),
    .C(_11074_),
    .Y(_11075_)
);

AOI21X1 _21020_ (
    .A(_11070_),
    .B(_11069_),
    .C(_11068_),
    .Y(_11076_)
);

NOR3X1 _21021_ (
    .A(_11061_),
    .B(_11064_),
    .C(_11065_),
    .Y(_11078_)
);

NOR2X1 _21022_ (
    .A(_10755_),
    .B(_10818_),
    .Y(_11079_)
);

OAI21X1 _21023_ (
    .A(_3402__bF$buf3),
    .B(_3781__bF$buf2),
    .C(_10755_),
    .Y(_11080_)
);

AOI21X1 _21024_ (
    .A(_10817_),
    .B(_11080_),
    .C(_11079_),
    .Y(_11081_)
);

OAI21X1 _21025_ (
    .A(_11078_),
    .B(_11076_),
    .C(_11081_),
    .Y(_11082_)
);

NAND3X1 _21026_ (
    .A(_11060_),
    .B(_11075_),
    .C(_11082_),
    .Y(_11083_)
);

INVX1 _21027_ (
    .A(_11060_),
    .Y(_11084_)
);

NAND3X1 _21028_ (
    .A(_11081_),
    .B(_11067_),
    .C(_11071_),
    .Y(_11085_)
);

OAI21X1 _21029_ (
    .A(_11078_),
    .B(_11076_),
    .C(_11074_),
    .Y(_11086_)
);

NAND3X1 _21030_ (
    .A(_11084_),
    .B(_11085_),
    .C(_11086_),
    .Y(_11087_)
);

AOI21X1 _21031_ (
    .A(_10837_),
    .B(_10841_),
    .C(_10821_),
    .Y(_11089_)
);

OAI21X1 _21032_ (
    .A(_10820_),
    .B(_11089_),
    .C(_10845_),
    .Y(_11090_)
);

NAND3X1 _21033_ (
    .A(_11083_),
    .B(_11087_),
    .C(_11090_),
    .Y(_11091_)
);

AOI21X1 _21034_ (
    .A(_11085_),
    .B(_11086_),
    .C(_11084_),
    .Y(_11092_)
);

AOI21X1 _21035_ (
    .A(_11075_),
    .B(_11082_),
    .C(_11060_),
    .Y(_11093_)
);

NOR3X1 _21036_ (
    .A(_10833_),
    .B(_10835_),
    .C(_10828_),
    .Y(_11094_)
);

AOI21X1 _21037_ (
    .A(_10846_),
    .B(_10844_),
    .C(_11094_),
    .Y(_11095_)
);

OAI21X1 _21038_ (
    .A(_11092_),
    .B(_11093_),
    .C(_11095_),
    .Y(_11096_)
);

NAND3X1 _21039_ (
    .A(_11059_),
    .B(_11096_),
    .C(_11091_),
    .Y(_11097_)
);

AND2X2 _21040_ (
    .A(_10766_),
    .B(_10758_),
    .Y(_11098_)
);

NOR3X1 _21041_ (
    .A(_11092_),
    .B(_11093_),
    .C(_11095_),
    .Y(_11100_)
);

AOI21X1 _21042_ (
    .A(_11083_),
    .B(_11087_),
    .C(_11090_),
    .Y(_11101_)
);

OAI21X1 _21043_ (
    .A(_11100_),
    .B(_11101_),
    .C(_11098_),
    .Y(_11102_)
);

NAND3X1 _21044_ (
    .A(_11097_),
    .B(_11102_),
    .C(_11058_),
    .Y(_11103_)
);

AOI21X1 _21045_ (
    .A(_10742_),
    .B(_10779_),
    .C(_10783_),
    .Y(_11104_)
);

NAND3X1 _21046_ (
    .A(_11083_),
    .B(_11087_),
    .C(_11095_),
    .Y(_11105_)
);

OAI21X1 _21047_ (
    .A(_11092_),
    .B(_11093_),
    .C(_11090_),
    .Y(_11106_)
);

AOI21X1 _21048_ (
    .A(_11106_),
    .B(_11105_),
    .C(_11098_),
    .Y(_11107_)
);

AOI21X1 _21049_ (
    .A(_11096_),
    .B(_11091_),
    .C(_11059_),
    .Y(_11108_)
);

OAI21X1 _21050_ (
    .A(_11107_),
    .B(_11108_),
    .C(_11104_),
    .Y(_11109_)
);

NAND3X1 _21051_ (
    .A(_11103_),
    .B(_11109_),
    .C(_11057_),
    .Y(_11111_)
);

NAND2X1 _21052_ (
    .A(_11056_),
    .B(_11052_),
    .Y(_11112_)
);

OAI21X1 _21053_ (
    .A(_11107_),
    .B(_11108_),
    .C(_11058_),
    .Y(_11113_)
);

NAND3X1 _21054_ (
    .A(_11104_),
    .B(_11097_),
    .C(_11102_),
    .Y(_11114_)
);

NAND3X1 _21055_ (
    .A(_11113_),
    .B(_11112_),
    .C(_11114_),
    .Y(_11115_)
);

AOI21X1 _21056_ (
    .A(_10889_),
    .B(_10894_),
    .C(_10896_),
    .Y(_11116_)
);

OAI21X1 _21057_ (
    .A(_11116_),
    .B(_10905_),
    .C(_10897_),
    .Y(_11117_)
);

NAND3X1 _21058_ (
    .A(_11115_),
    .B(_11117_),
    .C(_11111_),
    .Y(_11118_)
);

AOI21X1 _21059_ (
    .A(_11113_),
    .B(_11114_),
    .C(_11112_),
    .Y(_11119_)
);

AOI21X1 _21060_ (
    .A(_11103_),
    .B(_11109_),
    .C(_11057_),
    .Y(_11120_)
);

NOR3X1 _21061_ (
    .A(_10898_),
    .B(_10901_),
    .C(_10899_),
    .Y(_11122_)
);

AOI21X1 _21062_ (
    .A(_10815_),
    .B(_10903_),
    .C(_11122_),
    .Y(_11123_)
);

OAI21X1 _21063_ (
    .A(_11120_),
    .B(_11119_),
    .C(_11123_),
    .Y(_11124_)
);

NAND3X1 _21064_ (
    .A(_11015_),
    .B(_11118_),
    .C(_11124_),
    .Y(_11125_)
);

AND2X2 _21065_ (
    .A(_10794_),
    .B(_10786_),
    .Y(_11126_)
);

NAND3X1 _21066_ (
    .A(_11115_),
    .B(_11111_),
    .C(_11123_),
    .Y(_11127_)
);

OAI21X1 _21067_ (
    .A(_11120_),
    .B(_11119_),
    .C(_11117_),
    .Y(_11128_)
);

NAND3X1 _21068_ (
    .A(_11128_),
    .B(_11127_),
    .C(_11126_),
    .Y(_11129_)
);

NAND2X1 _21069_ (
    .A(_11125_),
    .B(_11129_),
    .Y(_11130_)
);

NOR2X1 _21070_ (
    .A(_10950_),
    .B(_10605_),
    .Y(_11131_)
);

AND2X2 _21071_ (
    .A(_10889_),
    .B(_10882_),
    .Y(_11133_)
);

NAND2X1 _21072_ (
    .A(areg_18_bF$buf0),
    .B(breg_23_bF$buf1),
    .Y(_11134_)
);

NAND2X1 _21073_ (
    .A(areg_20_bF$buf2),
    .B(breg_22_bF$buf4),
    .Y(_11135_)
);

OAI21X1 _21074_ (
    .A(_3958__bF$buf1),
    .B(_3781__bF$buf1),
    .C(_11072_),
    .Y(_11136_)
);

OAI21X1 _21075_ (
    .A(_10818_),
    .B(_11135_),
    .C(_11136_),
    .Y(_11137_)
);

XNOR2X1 _21076_ (
    .A(_11137_),
    .B(_11134_),
    .Y(_11138_)
);

AOI21X1 _21077_ (
    .A(_10829_),
    .B(_10832_),
    .C(_10839_),
    .Y(_11139_)
);

NAND2X1 _21078_ (
    .A(breg_20_bF$buf1),
    .B(areg_21_bF$buf4),
    .Y(_11140_)
);

AND2X2 _21079_ (
    .A(breg_18_bF$buf3),
    .B(areg_23_bF$buf3),
    .Y(_11141_)
);

OAI21X1 _21080_ (
    .A(_3253__bF$buf1),
    .B(_4551__bF$buf0),
    .C(_11141_),
    .Y(_11142_)
);

AND2X2 _21081_ (
    .A(breg_19_bF$buf4),
    .B(areg_22_bF$buf4),
    .Y(_11144_)
);

OAI21X1 _21082_ (
    .A(_3529__bF$buf3),
    .B(_4541__bF$buf3),
    .C(_11144_),
    .Y(_11145_)
);

AOI21X1 _21083_ (
    .A(_11142_),
    .B(_11145_),
    .C(_11140_),
    .Y(_11146_)
);

INVX2 _21084_ (
    .A(_11140_),
    .Y(_11147_)
);

NAND2X1 _21085_ (
    .A(_11144_),
    .B(_11141_),
    .Y(_11148_)
);

OAI22X1 _21086_ (
    .A(_3529__bF$buf2),
    .B(_4541__bF$buf2),
    .C(_3253__bF$buf0),
    .D(_4551__bF$buf4),
    .Y(_11149_)
);

AOI21X1 _21087_ (
    .A(_11149_),
    .B(_11148_),
    .C(_11147_),
    .Y(_11150_)
);

NOR3X1 _21088_ (
    .A(_11150_),
    .B(_11139_),
    .C(_11146_),
    .Y(_11151_)
);

OAI21X1 _21089_ (
    .A(_10840_),
    .B(_10822_),
    .C(_10830_),
    .Y(_11152_)
);

NAND3X1 _21090_ (
    .A(_11147_),
    .B(_11149_),
    .C(_11148_),
    .Y(_11153_)
);

NAND2X1 _21091_ (
    .A(breg_19_bF$buf3),
    .B(areg_23_bF$buf2),
    .Y(_11155_)
);

NOR2X1 _21092_ (
    .A(_10838_),
    .B(_11155_),
    .Y(_11156_)
);

NOR2X1 _21093_ (
    .A(_11144_),
    .B(_11141_),
    .Y(_11157_)
);

OAI21X1 _21094_ (
    .A(_11157_),
    .B(_11156_),
    .C(_11140_),
    .Y(_11158_)
);

AOI21X1 _21095_ (
    .A(_11153_),
    .B(_11158_),
    .C(_11152_),
    .Y(_11159_)
);

NOR3X1 _21096_ (
    .A(_11138_),
    .B(_11159_),
    .C(_11151_),
    .Y(_11160_)
);

INVX2 _21097_ (
    .A(_11134_),
    .Y(_11161_)
);

XNOR2X1 _21098_ (
    .A(_11137_),
    .B(_11161_),
    .Y(_11162_)
);

NAND3X1 _21099_ (
    .A(_11153_),
    .B(_11152_),
    .C(_11158_),
    .Y(_11163_)
);

OAI21X1 _21100_ (
    .A(_11146_),
    .B(_11150_),
    .C(_11139_),
    .Y(_11164_)
);

AOI21X1 _21101_ (
    .A(_11164_),
    .B(_11163_),
    .C(_11162_),
    .Y(_11166_)
);

NOR2X1 _21102_ (
    .A(_11166_),
    .B(_11160_),
    .Y(_11167_)
);

OAI21X1 _21103_ (
    .A(_10879_),
    .B(_10877_),
    .C(_10868_),
    .Y(_11168_)
);

OAI21X1 _21104_ (
    .A(_10863_),
    .B(_10853_),
    .C(_10857_),
    .Y(_11169_)
);

NAND2X1 _21105_ (
    .A(breg_17_bF$buf4),
    .B(areg_24_bF$buf1),
    .Y(_11170_)
);

INVX1 _21106_ (
    .A(_11170_),
    .Y(_11171_)
);

AND2X2 _21107_ (
    .A(breg_16_bF$buf4),
    .B(areg_25_bF$buf3),
    .Y(_11172_)
);

AND2X2 _21108_ (
    .A(breg_15_bF$buf0),
    .B(areg_26_bF$buf4),
    .Y(_11173_)
);

NAND2X1 _21109_ (
    .A(_11172_),
    .B(_11173_),
    .Y(_11174_)
);

OAI22X1 _21110_ (
    .A(_2362__bF$buf5),
    .B(_6686__bF$buf0),
    .C(_2560__bF$buf3),
    .D(_6300__bF$buf1),
    .Y(_11175_)
);

NAND3X1 _21111_ (
    .A(_11171_),
    .B(_11175_),
    .C(_11174_),
    .Y(_11177_)
);

OAI21X1 _21112_ (
    .A(_2560__bF$buf2),
    .B(_6300__bF$buf0),
    .C(_11173_),
    .Y(_11178_)
);

OAI21X1 _21113_ (
    .A(_2362__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_11172_),
    .Y(_11179_)
);

NAND3X1 _21114_ (
    .A(_11170_),
    .B(_11178_),
    .C(_11179_),
    .Y(_11180_)
);

NAND2X1 _21115_ (
    .A(breg_13_bF$buf1),
    .B(areg_28_bF$buf3),
    .Y(_11181_)
);

AND2X2 _21116_ (
    .A(_10865_),
    .B(_10912_),
    .Y(_11182_)
);

OAI22X1 _21117_ (
    .A(_10558_),
    .B(_11181_),
    .C(_11182_),
    .D(_10911_),
    .Y(_11183_)
);

NAND3X1 _21118_ (
    .A(_11177_),
    .B(_11180_),
    .C(_11183_),
    .Y(_11184_)
);

AOI21X1 _21119_ (
    .A(_11178_),
    .B(_11179_),
    .C(_11170_),
    .Y(_11185_)
);

AOI21X1 _21120_ (
    .A(_11175_),
    .B(_11174_),
    .C(_11171_),
    .Y(_11186_)
);

NOR2X1 _21121_ (
    .A(_10865_),
    .B(_10912_),
    .Y(_11188_)
);

OAI21X1 _21122_ (
    .A(_2586__bF$buf0),
    .B(_7520__bF$buf2),
    .C(_10865_),
    .Y(_11189_)
);

AOI21X1 _21123_ (
    .A(_10933_),
    .B(_11189_),
    .C(_11188_),
    .Y(_11190_)
);

OAI21X1 _21124_ (
    .A(_11185_),
    .B(_11186_),
    .C(_11190_),
    .Y(_11191_)
);

NAND3X1 _21125_ (
    .A(_11169_),
    .B(_11184_),
    .C(_11191_),
    .Y(_11192_)
);

INVX2 _21126_ (
    .A(_11169_),
    .Y(_11193_)
);

NOR3X1 _21127_ (
    .A(_11186_),
    .B(_11190_),
    .C(_11185_),
    .Y(_11194_)
);

AOI21X1 _21128_ (
    .A(_11177_),
    .B(_11180_),
    .C(_11183_),
    .Y(_11195_)
);

OAI21X1 _21129_ (
    .A(_11194_),
    .B(_11195_),
    .C(_11193_),
    .Y(_11196_)
);

NAND3X1 _21130_ (
    .A(_11168_),
    .B(_11192_),
    .C(_11196_),
    .Y(_11197_)
);

AOI21X1 _21131_ (
    .A(_10852_),
    .B(_10875_),
    .C(_10878_),
    .Y(_11199_)
);

NAND3X1 _21132_ (
    .A(_11190_),
    .B(_11177_),
    .C(_11180_),
    .Y(_11200_)
);

OAI21X1 _21133_ (
    .A(_11185_),
    .B(_11186_),
    .C(_11183_),
    .Y(_11201_)
);

AOI21X1 _21134_ (
    .A(_11200_),
    .B(_11201_),
    .C(_11193_),
    .Y(_11202_)
);

AOI21X1 _21135_ (
    .A(_11184_),
    .B(_11191_),
    .C(_11169_),
    .Y(_11203_)
);

OAI21X1 _21136_ (
    .A(_11202_),
    .B(_11203_),
    .C(_11199_),
    .Y(_11204_)
);

NAND3X1 _21137_ (
    .A(_11197_),
    .B(_11204_),
    .C(_11167_),
    .Y(_11205_)
);

OR2X2 _21138_ (
    .A(_11160_),
    .B(_11166_),
    .Y(_11206_)
);

OAI21X1 _21139_ (
    .A(_11202_),
    .B(_11203_),
    .C(_11168_),
    .Y(_11207_)
);

NAND3X1 _21140_ (
    .A(_11192_),
    .B(_11196_),
    .C(_11199_),
    .Y(_11208_)
);

NAND3X1 _21141_ (
    .A(_11207_),
    .B(_11208_),
    .C(_11206_),
    .Y(_11210_)
);

NOR3X1 _21142_ (
    .A(_10942_),
    .B(_10940_),
    .C(_10941_),
    .Y(_11211_)
);

AOI21X1 _21143_ (
    .A(_10910_),
    .B(_10943_),
    .C(_11211_),
    .Y(_11212_)
);

NAND3X1 _21144_ (
    .A(_11205_),
    .B(_11212_),
    .C(_11210_),
    .Y(_11213_)
);

AOI21X1 _21145_ (
    .A(_11207_),
    .B(_11208_),
    .C(_11206_),
    .Y(_11214_)
);

AOI21X1 _21146_ (
    .A(_11204_),
    .B(_11197_),
    .C(_11167_),
    .Y(_11215_)
);

AOI21X1 _21147_ (
    .A(_10932_),
    .B(_10938_),
    .C(_10258_),
    .Y(_11216_)
);

OAI21X1 _21148_ (
    .A(_11216_),
    .B(_10945_),
    .C(_10939_),
    .Y(_11217_)
);

OAI21X1 _21149_ (
    .A(_11214_),
    .B(_11215_),
    .C(_11217_),
    .Y(_11218_)
);

AOI21X1 _21150_ (
    .A(_11213_),
    .B(_11218_),
    .C(_11133_),
    .Y(_11219_)
);

NAND2X1 _21151_ (
    .A(_10882_),
    .B(_10889_),
    .Y(_11221_)
);

NAND3X1 _21152_ (
    .A(_11205_),
    .B(_11217_),
    .C(_11210_),
    .Y(_11222_)
);

OAI21X1 _21153_ (
    .A(_11214_),
    .B(_11215_),
    .C(_11212_),
    .Y(_11223_)
);

AOI21X1 _21154_ (
    .A(_11222_),
    .B(_11223_),
    .C(_11221_),
    .Y(_11224_)
);

AND2X2 _21155_ (
    .A(_10932_),
    .B(_10927_),
    .Y(_11225_)
);

NAND2X1 _21156_ (
    .A(breg_14_bF$buf2),
    .B(areg_27_bF$buf2),
    .Y(_11226_)
);

INVX2 _21157_ (
    .A(_11226_),
    .Y(_11227_)
);

NAND2X1 _21158_ (
    .A(breg_13_bF$buf0),
    .B(areg_29_bF$buf0),
    .Y(_11228_)
);

INVX1 _21159_ (
    .A(breg_13_bF$buf4),
    .Y(_11229_)
);

NAND2X1 _21160_ (
    .A(breg_12_bF$buf4),
    .B(areg_29_bF$buf5),
    .Y(_11230_)
);

OAI21X1 _21161_ (
    .A(_11229_),
    .B(_7520__bF$buf1),
    .C(_11230_),
    .Y(_11232_)
);

OAI21X1 _21162_ (
    .A(_10912_),
    .B(_11228_),
    .C(_11232_),
    .Y(_11233_)
);

XNOR2X1 _21163_ (
    .A(_11233_),
    .B(_11227_),
    .Y(_11234_)
);

INVX2 _21164_ (
    .A(_11234_),
    .Y(_11235_)
);

NAND2X1 _21165_ (
    .A(_10920_),
    .B(_10922_),
    .Y(_11236_)
);

NAND2X1 _21166_ (
    .A(breg_11_bF$buf1),
    .B(areg_31_bF$buf4),
    .Y(_11237_)
);

NOR2X1 _21167_ (
    .A(_10570_),
    .B(_11237_),
    .Y(_11238_)
);

AOI22X1 _21168_ (
    .A(breg_10_bF$buf3),
    .B(areg_31_bF$buf3),
    .C(breg_11_bF$buf0),
    .D(areg_30_bF$buf4),
    .Y(_11239_)
);

NOR2X1 _21169_ (
    .A(_11239_),
    .B(_11238_),
    .Y(_11240_)
);

NOR2X1 _21170_ (
    .A(_11240_),
    .B(_11236_),
    .Y(_11241_)
);

AND2X2 _21171_ (
    .A(_11236_),
    .B(_11240_),
    .Y(_11243_)
);

OAI21X1 _21172_ (
    .A(_11243_),
    .B(_11241_),
    .C(_11235_),
    .Y(_11244_)
);

INVX1 _21173_ (
    .A(_11244_),
    .Y(_11245_)
);

XNOR2X1 _21174_ (
    .A(_11236_),
    .B(_11240_),
    .Y(_11246_)
);

NOR2X1 _21175_ (
    .A(_11235_),
    .B(_11246_),
    .Y(_11247_)
);

OAI21X1 _21176_ (
    .A(_11245_),
    .B(_11247_),
    .C(_11225_),
    .Y(_11248_)
);

NAND2X1 _21177_ (
    .A(_10927_),
    .B(_10932_),
    .Y(_11249_)
);

OR2X2 _21178_ (
    .A(_11246_),
    .B(_11235_),
    .Y(_11250_)
);

NAND3X1 _21179_ (
    .A(_11249_),
    .B(_11244_),
    .C(_11250_),
    .Y(_11251_)
);

NAND2X1 _21180_ (
    .A(_11251_),
    .B(_11248_),
    .Y(_11252_)
);

OAI21X1 _21181_ (
    .A(_11219_),
    .B(_11224_),
    .C(_11252_),
    .Y(_11254_)
);

NAND3X1 _21182_ (
    .A(_11221_),
    .B(_11222_),
    .C(_11223_),
    .Y(_11255_)
);

NAND3X1 _21183_ (
    .A(_11133_),
    .B(_11213_),
    .C(_11218_),
    .Y(_11256_)
);

INVX1 _21184_ (
    .A(_11252_),
    .Y(_11257_)
);

NAND3X1 _21185_ (
    .A(_11257_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11258_)
);

NAND2X1 _21186_ (
    .A(_11258_),
    .B(_11254_),
    .Y(_11259_)
);

OAI21X1 _21187_ (
    .A(_10952_),
    .B(_11131_),
    .C(_11259_),
    .Y(_11260_)
);

NOR2X1 _21188_ (
    .A(_10953_),
    .B(_10954_),
    .Y(_11261_)
);

AOI21X1 _21189_ (
    .A(_10961_),
    .B(_11261_),
    .C(_11131_),
    .Y(_11262_)
);

AND2X2 _21190_ (
    .A(_11254_),
    .B(_11258_),
    .Y(_11263_)
);

NAND2X1 _21191_ (
    .A(_11262_),
    .B(_11263_),
    .Y(_11265_)
);

AOI21X1 _21192_ (
    .A(_11260_),
    .B(_11265_),
    .C(_11130_),
    .Y(_11266_)
);

NAND3X1 _21193_ (
    .A(_11118_),
    .B(_11124_),
    .C(_11126_),
    .Y(_11267_)
);

NAND3X1 _21194_ (
    .A(_11015_),
    .B(_11128_),
    .C(_11127_),
    .Y(_11268_)
);

NAND2X1 _21195_ (
    .A(_11268_),
    .B(_11267_),
    .Y(_11269_)
);

INVX1 _21196_ (
    .A(_11131_),
    .Y(_11270_)
);

OAI21X1 _21197_ (
    .A(_10909_),
    .B(_10951_),
    .C(_11270_),
    .Y(_11271_)
);

NAND3X1 _21198_ (
    .A(_11254_),
    .B(_11258_),
    .C(_11271_),
    .Y(_11272_)
);

NAND2X1 _21199_ (
    .A(_11259_),
    .B(_11262_),
    .Y(_11273_)
);

AOI21X1 _21200_ (
    .A(_11272_),
    .B(_11273_),
    .C(_11269_),
    .Y(_11274_)
);

OAI21X1 _21201_ (
    .A(_11266_),
    .B(_11274_),
    .C(_11014_),
    .Y(_11276_)
);

NAND2X1 _21202_ (
    .A(_10955_),
    .B(_10962_),
    .Y(_11277_)
);

NOR2X1 _21203_ (
    .A(_10960_),
    .B(_11277_),
    .Y(_11278_)
);

AOI21X1 _21204_ (
    .A(_10967_),
    .B(_10970_),
    .C(_11278_),
    .Y(_11279_)
);

NAND3X1 _21205_ (
    .A(_11272_),
    .B(_11273_),
    .C(_11269_),
    .Y(_11280_)
);

NOR2X1 _21206_ (
    .A(_11259_),
    .B(_11262_),
    .Y(_11281_)
);

AOI21X1 _21207_ (
    .A(_11254_),
    .B(_11258_),
    .C(_11271_),
    .Y(_11282_)
);

OAI21X1 _21208_ (
    .A(_11281_),
    .B(_11282_),
    .C(_11130_),
    .Y(_11283_)
);

NAND3X1 _21209_ (
    .A(_11280_),
    .B(_11283_),
    .C(_11279_),
    .Y(_11284_)
);

AOI21X1 _21210_ (
    .A(_11284_),
    .B(_11276_),
    .C(_11012_),
    .Y(_11285_)
);

NAND3X1 _21211_ (
    .A(_11280_),
    .B(_11014_),
    .C(_11283_),
    .Y(_11287_)
);

OAI21X1 _21212_ (
    .A(_11266_),
    .B(_11274_),
    .C(_11279_),
    .Y(_11288_)
);

AOI21X1 _21213_ (
    .A(_11287_),
    .B(_11288_),
    .C(_11010_),
    .Y(_11289_)
);

OAI21X1 _21214_ (
    .A(_11285_),
    .B(_11289_),
    .C(_11009_),
    .Y(_11290_)
);

NOR3X1 _21215_ (
    .A(_10964_),
    .B(_10971_),
    .C(_10974_),
    .Y(_11291_)
);

AOI21X1 _21216_ (
    .A(_10981_),
    .B(_10694_),
    .C(_11291_),
    .Y(_11292_)
);

NAND3X1 _21217_ (
    .A(_11010_),
    .B(_11287_),
    .C(_11288_),
    .Y(_11293_)
);

NAND3X1 _21218_ (
    .A(_11012_),
    .B(_11284_),
    .C(_11276_),
    .Y(_11294_)
);

NAND3X1 _21219_ (
    .A(_11293_),
    .B(_11294_),
    .C(_11292_),
    .Y(_11295_)
);

AOI21X1 _21220_ (
    .A(_11295_),
    .B(_11290_),
    .C(_11007_),
    .Y(_11296_)
);

NAND3X1 _21221_ (
    .A(_11293_),
    .B(_11294_),
    .C(_11009_),
    .Y(_11298_)
);

OAI21X1 _21222_ (
    .A(_11285_),
    .B(_11289_),
    .C(_11292_),
    .Y(_11299_)
);

AOI21X1 _21223_ (
    .A(_11298_),
    .B(_11299_),
    .C(_11006_),
    .Y(_11300_)
);

OAI21X1 _21224_ (
    .A(_11296_),
    .B(_11300_),
    .C(_11005_),
    .Y(_11301_)
);

NOR3X1 _21225_ (
    .A(_10982_),
    .B(_10978_),
    .C(_10984_),
    .Y(_11302_)
);

AOI21X1 _21226_ (
    .A(_10690_),
    .B(_10991_),
    .C(_11302_),
    .Y(_11303_)
);

NAND3X1 _21227_ (
    .A(_11006_),
    .B(_11298_),
    .C(_11299_),
    .Y(_11304_)
);

NAND3X1 _21228_ (
    .A(_11007_),
    .B(_11295_),
    .C(_11290_),
    .Y(_11305_)
);

NAND3X1 _21229_ (
    .A(_11304_),
    .B(_11305_),
    .C(_11303_),
    .Y(_11306_)
);

NAND2X1 _21230_ (
    .A(_11306_),
    .B(_11301_),
    .Y(_11307_)
);

XNOR2X1 _21231_ (
    .A(_11003_),
    .B(_11307_),
    .Y(_0_[41])
);

OAI21X1 _21232_ (
    .A(_11296_),
    .B(_11300_),
    .C(_11303_),
    .Y(_11309_)
);

NAND3X1 _21233_ (
    .A(_11005_),
    .B(_11304_),
    .C(_11305_),
    .Y(_11310_)
);

OAI21X1 _21234_ (
    .A(_11001_),
    .B(_10994_),
    .C(_11310_),
    .Y(_11311_)
);

AND2X2 _21235_ (
    .A(_11311_),
    .B(_11309_),
    .Y(_11312_)
);

AOI22X1 _21236_ (
    .A(_11301_),
    .B(_11306_),
    .C(_10993_),
    .D(_10997_),
    .Y(_11313_)
);

AND2X2 _21237_ (
    .A(_10688_),
    .B(_11313_),
    .Y(_11314_)
);

NOR2X1 _21238_ (
    .A(_11312_),
    .B(_11314_),
    .Y(_11315_)
);

AOI21X1 _21239_ (
    .A(_11293_),
    .B(_11294_),
    .C(_11009_),
    .Y(_11316_)
);

OAI21X1 _21240_ (
    .A(_11316_),
    .B(_11007_),
    .C(_11298_),
    .Y(_11317_)
);

OAI21X1 _21241_ (
    .A(_11047_),
    .B(_11017_),
    .C(_11054_),
    .Y(_11319_)
);

INVX2 _21242_ (
    .A(_11319_),
    .Y(_11320_)
);

AOI21X1 _21243_ (
    .A(_11280_),
    .B(_11283_),
    .C(_11014_),
    .Y(_11321_)
);

OAI21X1 _21244_ (
    .A(_11321_),
    .B(_11012_),
    .C(_11287_),
    .Y(_11322_)
);

NAND2X1 _21245_ (
    .A(_11118_),
    .B(_11125_),
    .Y(_11323_)
);

INVX2 _21246_ (
    .A(_11323_),
    .Y(_11324_)
);

OAI21X1 _21247_ (
    .A(_11130_),
    .B(_11282_),
    .C(_11272_),
    .Y(_11325_)
);

NAND2X1 _21248_ (
    .A(_11103_),
    .B(_11111_),
    .Y(_11326_)
);

NOR2X1 _21249_ (
    .A(_9104__bF$buf0),
    .B(_7225__bF$buf3),
    .Y(_11327_)
);

INVX1 _21250_ (
    .A(_11327_),
    .Y(_11328_)
);

OAI21X1 _21251_ (
    .A(_11034_),
    .B(_11020_),
    .C(_11045_),
    .Y(_11330_)
);

NOR2X1 _21252_ (
    .A(_10869__bF$buf2),
    .B(_6815__bF$buf2),
    .Y(_11331_)
);

INVX2 _21253_ (
    .A(_11331_),
    .Y(_11332_)
);

OAI21X1 _21254_ (
    .A(_11032_),
    .B(_11023_),
    .C(_11027_),
    .Y(_11333_)
);

NAND2X1 _21255_ (
    .A(areg_13_bF$buf3),
    .B(breg_29_bF$buf1),
    .Y(_11334_)
);

INVX2 _21256_ (
    .A(_11334_),
    .Y(_11335_)
);

AND2X2 _21257_ (
    .A(areg_14_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_11336_)
);

AND2X2 _21258_ (
    .A(areg_15_bF$buf1),
    .B(breg_27_bF$buf3),
    .Y(_11337_)
);

NAND2X1 _21259_ (
    .A(_11336_),
    .B(_11337_),
    .Y(_11338_)
);

OAI21X1 _21260_ (
    .A(_2465__bF$buf3),
    .B(_5668__bF$buf5),
    .C(_11030_),
    .Y(_11339_)
);

NAND3X1 _21261_ (
    .A(_11335_),
    .B(_11339_),
    .C(_11338_),
    .Y(_11340_)
);

NAND2X1 _21262_ (
    .A(areg_15_bF$buf0),
    .B(breg_27_bF$buf2),
    .Y(_11341_)
);

NOR2X1 _21263_ (
    .A(_11030_),
    .B(_11341_),
    .Y(_11342_)
);

NOR2X1 _21264_ (
    .A(_11336_),
    .B(_11337_),
    .Y(_11343_)
);

OAI21X1 _21265_ (
    .A(_11343_),
    .B(_11342_),
    .C(_11334_),
    .Y(_11344_)
);

AOI21X1 _21266_ (
    .A(_11340_),
    .B(_11344_),
    .C(_11333_),
    .Y(_11345_)
);

AOI21X1 _21267_ (
    .A(_11024_),
    .B(_11028_),
    .C(_11031_),
    .Y(_11346_)
);

OAI21X1 _21268_ (
    .A(_2287__bF$buf0),
    .B(_6050__bF$buf2),
    .C(_11337_),
    .Y(_11347_)
);

OAI21X1 _21269_ (
    .A(_2465__bF$buf2),
    .B(_5668__bF$buf4),
    .C(_11336_),
    .Y(_11348_)
);

AOI21X1 _21270_ (
    .A(_11347_),
    .B(_11348_),
    .C(_11334_),
    .Y(_11349_)
);

AOI21X1 _21271_ (
    .A(_11339_),
    .B(_11338_),
    .C(_11335_),
    .Y(_11351_)
);

NOR3X1 _21272_ (
    .A(_11351_),
    .B(_11346_),
    .C(_11349_),
    .Y(_11352_)
);

OAI21X1 _21273_ (
    .A(_11352_),
    .B(_11345_),
    .C(_11332_),
    .Y(_11353_)
);

OAI21X1 _21274_ (
    .A(_11349_),
    .B(_11351_),
    .C(_11346_),
    .Y(_11354_)
);

NAND3X1 _21275_ (
    .A(_11340_),
    .B(_11344_),
    .C(_11333_),
    .Y(_11355_)
);

NAND3X1 _21276_ (
    .A(_11331_),
    .B(_11354_),
    .C(_11355_),
    .Y(_11356_)
);

AOI21X1 _21277_ (
    .A(_11356_),
    .B(_11353_),
    .C(_11330_),
    .Y(_11357_)
);

AOI21X1 _21278_ (
    .A(_11019_),
    .B(_11042_),
    .C(_11040_),
    .Y(_11358_)
);

AOI21X1 _21279_ (
    .A(_11354_),
    .B(_11355_),
    .C(_11331_),
    .Y(_11359_)
);

NOR3X1 _21280_ (
    .A(_11345_),
    .B(_11332_),
    .C(_11352_),
    .Y(_11360_)
);

NOR3X1 _21281_ (
    .A(_11358_),
    .B(_11359_),
    .C(_11360_),
    .Y(_11363_)
);

OAI21X1 _21282_ (
    .A(_11363_),
    .B(_11357_),
    .C(_11328_),
    .Y(_11364_)
);

OAI21X1 _21283_ (
    .A(_11360_),
    .B(_11359_),
    .C(_11358_),
    .Y(_11365_)
);

NAND3X1 _21284_ (
    .A(_11330_),
    .B(_11356_),
    .C(_11353_),
    .Y(_11366_)
);

NAND3X1 _21285_ (
    .A(_11327_),
    .B(_11366_),
    .C(_11365_),
    .Y(_11367_)
);

AND2X2 _21286_ (
    .A(_11364_),
    .B(_11367_),
    .Y(_11368_)
);

OAI21X1 _21287_ (
    .A(_11101_),
    .B(_11098_),
    .C(_11091_),
    .Y(_11369_)
);

NAND2X1 _21288_ (
    .A(_11075_),
    .B(_11083_),
    .Y(_11370_)
);

OAI21X1 _21289_ (
    .A(_11065_),
    .B(_11061_),
    .C(_11069_),
    .Y(_11371_)
);

NAND2X1 _21290_ (
    .A(areg_16_bF$buf5),
    .B(breg_26_bF$buf3),
    .Y(_11372_)
);

NAND2X1 _21291_ (
    .A(areg_17_bF$buf5),
    .B(breg_25_bF$buf1),
    .Y(_11374_)
);

NAND2X1 _21292_ (
    .A(areg_18_bF$buf5),
    .B(breg_24_bF$buf2),
    .Y(_11375_)
);

NOR2X1 _21293_ (
    .A(_11374_),
    .B(_11375_),
    .Y(_11376_)
);

AOI22X1 _21294_ (
    .A(areg_17_bF$buf4),
    .B(breg_25_bF$buf0),
    .C(areg_18_bF$buf4),
    .D(breg_24_bF$buf1),
    .Y(_11377_)
);

OAI21X1 _21295_ (
    .A(_11376_),
    .B(_11377_),
    .C(_11372_),
    .Y(_11378_)
);

INVX1 _21296_ (
    .A(_11372_),
    .Y(_11379_)
);

OR2X2 _21297_ (
    .A(_11374_),
    .B(_11375_),
    .Y(_11380_)
);

INVX1 _21298_ (
    .A(_11377_),
    .Y(_11381_)
);

NAND3X1 _21299_ (
    .A(_11379_),
    .B(_11381_),
    .C(_11380_),
    .Y(_11382_)
);

NAND2X1 _21300_ (
    .A(areg_20_bF$buf1),
    .B(breg_21_bF$buf0),
    .Y(_11383_)
);

AND2X2 _21301_ (
    .A(_11072_),
    .B(_11383_),
    .Y(_11385_)
);

OAI22X1 _21302_ (
    .A(_10818_),
    .B(_11135_),
    .C(_11385_),
    .D(_11134_),
    .Y(_11386_)
);

NAND3X1 _21303_ (
    .A(_11378_),
    .B(_11382_),
    .C(_11386_),
    .Y(_11387_)
);

AOI21X1 _21304_ (
    .A(_11381_),
    .B(_11380_),
    .C(_11379_),
    .Y(_11388_)
);

NOR3X1 _21305_ (
    .A(_11372_),
    .B(_11377_),
    .C(_11376_),
    .Y(_11389_)
);

NOR2X1 _21306_ (
    .A(_11072_),
    .B(_11383_),
    .Y(_11390_)
);

AOI21X1 _21307_ (
    .A(_11161_),
    .B(_11136_),
    .C(_11390_),
    .Y(_11391_)
);

OAI21X1 _21308_ (
    .A(_11388_),
    .B(_11389_),
    .C(_11391_),
    .Y(_11392_)
);

NAND3X1 _21309_ (
    .A(_11371_),
    .B(_11387_),
    .C(_11392_),
    .Y(_11393_)
);

INVX1 _21310_ (
    .A(_11371_),
    .Y(_11394_)
);

NAND3X1 _21311_ (
    .A(_11391_),
    .B(_11378_),
    .C(_11382_),
    .Y(_11396_)
);

OAI21X1 _21312_ (
    .A(_11388_),
    .B(_11389_),
    .C(_11386_),
    .Y(_11397_)
);

NAND3X1 _21313_ (
    .A(_11396_),
    .B(_11394_),
    .C(_11397_),
    .Y(_11398_)
);

OAI21X1 _21314_ (
    .A(_11138_),
    .B(_11159_),
    .C(_11163_),
    .Y(_11399_)
);

NAND3X1 _21315_ (
    .A(_11393_),
    .B(_11398_),
    .C(_11399_),
    .Y(_11400_)
);

AOI21X1 _21316_ (
    .A(_11396_),
    .B(_11397_),
    .C(_11394_),
    .Y(_11401_)
);

AOI21X1 _21317_ (
    .A(_11387_),
    .B(_11392_),
    .C(_11371_),
    .Y(_11402_)
);

AOI21X1 _21318_ (
    .A(_11164_),
    .B(_11162_),
    .C(_11151_),
    .Y(_11403_)
);

OAI21X1 _21319_ (
    .A(_11402_),
    .B(_11401_),
    .C(_11403_),
    .Y(_11404_)
);

NAND3X1 _21320_ (
    .A(_11370_),
    .B(_11400_),
    .C(_11404_),
    .Y(_11405_)
);

AND2X2 _21321_ (
    .A(_11083_),
    .B(_11075_),
    .Y(_11407_)
);

NOR3X1 _21322_ (
    .A(_11401_),
    .B(_11402_),
    .C(_11403_),
    .Y(_11408_)
);

AOI21X1 _21323_ (
    .A(_11393_),
    .B(_11398_),
    .C(_11399_),
    .Y(_11409_)
);

OAI21X1 _21324_ (
    .A(_11408_),
    .B(_11409_),
    .C(_11407_),
    .Y(_11410_)
);

NAND3X1 _21325_ (
    .A(_11369_),
    .B(_11405_),
    .C(_11410_),
    .Y(_11411_)
);

AOI21X1 _21326_ (
    .A(_11059_),
    .B(_11096_),
    .C(_11100_),
    .Y(_11412_)
);

NAND3X1 _21327_ (
    .A(_11398_),
    .B(_11393_),
    .C(_11403_),
    .Y(_11413_)
);

OAI21X1 _21328_ (
    .A(_11402_),
    .B(_11401_),
    .C(_11399_),
    .Y(_11414_)
);

AOI21X1 _21329_ (
    .A(_11413_),
    .B(_11414_),
    .C(_11407_),
    .Y(_11415_)
);

AOI21X1 _21330_ (
    .A(_11400_),
    .B(_11404_),
    .C(_11370_),
    .Y(_11416_)
);

OAI21X1 _21331_ (
    .A(_11416_),
    .B(_11415_),
    .C(_11412_),
    .Y(_11418_)
);

NAND3X1 _21332_ (
    .A(_11411_),
    .B(_11418_),
    .C(_11368_),
    .Y(_11419_)
);

NAND2X1 _21333_ (
    .A(_11367_),
    .B(_11364_),
    .Y(_11420_)
);

OAI21X1 _21334_ (
    .A(_11416_),
    .B(_11415_),
    .C(_11369_),
    .Y(_11421_)
);

NAND3X1 _21335_ (
    .A(_11405_),
    .B(_11412_),
    .C(_11410_),
    .Y(_11422_)
);

NAND3X1 _21336_ (
    .A(_11421_),
    .B(_11420_),
    .C(_11422_),
    .Y(_11423_)
);

AOI21X1 _21337_ (
    .A(_11205_),
    .B(_11210_),
    .C(_11217_),
    .Y(_11424_)
);

OAI21X1 _21338_ (
    .A(_11424_),
    .B(_11133_),
    .C(_11222_),
    .Y(_11425_)
);

NAND3X1 _21339_ (
    .A(_11423_),
    .B(_11425_),
    .C(_11419_),
    .Y(_11426_)
);

AOI21X1 _21340_ (
    .A(_11421_),
    .B(_11422_),
    .C(_11420_),
    .Y(_11427_)
);

AOI21X1 _21341_ (
    .A(_11411_),
    .B(_11418_),
    .C(_11368_),
    .Y(_11429_)
);

NOR3X1 _21342_ (
    .A(_11212_),
    .B(_11215_),
    .C(_11214_),
    .Y(_11430_)
);

AOI21X1 _21343_ (
    .A(_11221_),
    .B(_11223_),
    .C(_11430_),
    .Y(_11431_)
);

OAI21X1 _21344_ (
    .A(_11429_),
    .B(_11427_),
    .C(_11431_),
    .Y(_11432_)
);

NAND3X1 _21345_ (
    .A(_11326_),
    .B(_11426_),
    .C(_11432_),
    .Y(_11433_)
);

AND2X2 _21346_ (
    .A(_11111_),
    .B(_11103_),
    .Y(_11434_)
);

NAND3X1 _21347_ (
    .A(_11423_),
    .B(_11419_),
    .C(_11431_),
    .Y(_11435_)
);

OAI21X1 _21348_ (
    .A(_11429_),
    .B(_11427_),
    .C(_11425_),
    .Y(_11436_)
);

NAND3X1 _21349_ (
    .A(_11436_),
    .B(_11435_),
    .C(_11434_),
    .Y(_11437_)
);

NAND2X1 _21350_ (
    .A(_11433_),
    .B(_11437_),
    .Y(_11438_)
);

AND2X2 _21351_ (
    .A(_11205_),
    .B(_11197_),
    .Y(_11440_)
);

NAND2X1 _21352_ (
    .A(areg_19_bF$buf1),
    .B(breg_23_bF$buf0),
    .Y(_11441_)
);

NAND2X1 _21353_ (
    .A(areg_21_bF$buf3),
    .B(breg_22_bF$buf3),
    .Y(_11442_)
);

OAI21X1 _21354_ (
    .A(_3961__bF$buf1),
    .B(_3781__bF$buf0),
    .C(_11135_),
    .Y(_11443_)
);

OAI21X1 _21355_ (
    .A(_11383_),
    .B(_11442_),
    .C(_11443_),
    .Y(_11444_)
);

XNOR2X1 _21356_ (
    .A(_11444_),
    .B(_11441_),
    .Y(_11445_)
);

OAI21X1 _21357_ (
    .A(_11157_),
    .B(_11140_),
    .C(_11148_),
    .Y(_11446_)
);

NAND2X1 _21358_ (
    .A(breg_20_bF$buf0),
    .B(areg_22_bF$buf3),
    .Y(_11447_)
);

NAND2X1 _21359_ (
    .A(breg_18_bF$buf2),
    .B(areg_24_bF$buf0),
    .Y(_11448_)
);

NOR2X1 _21360_ (
    .A(_11155_),
    .B(_11448_),
    .Y(_11449_)
);

AND2X2 _21361_ (
    .A(breg_19_bF$buf2),
    .B(areg_23_bF$buf1),
    .Y(_11451_)
);

AND2X2 _21362_ (
    .A(breg_18_bF$buf1),
    .B(areg_24_bF$buf4),
    .Y(_11452_)
);

NOR2X1 _21363_ (
    .A(_11451_),
    .B(_11452_),
    .Y(_11453_)
);

NOR3X1 _21364_ (
    .A(_11447_),
    .B(_11449_),
    .C(_11453_),
    .Y(_11454_)
);

INVX2 _21365_ (
    .A(_11447_),
    .Y(_11455_)
);

NAND2X1 _21366_ (
    .A(_11451_),
    .B(_11452_),
    .Y(_11456_)
);

OAI21X1 _21367_ (
    .A(_3529__bF$buf1),
    .B(_5921__bF$buf1),
    .C(_11155_),
    .Y(_11457_)
);

AOI21X1 _21368_ (
    .A(_11457_),
    .B(_11456_),
    .C(_11455_),
    .Y(_11458_)
);

OAI21X1 _21369_ (
    .A(_11454_),
    .B(_11458_),
    .C(_11446_),
    .Y(_11459_)
);

AOI21X1 _21370_ (
    .A(_11147_),
    .B(_11149_),
    .C(_11156_),
    .Y(_11460_)
);

NAND3X1 _21371_ (
    .A(_11455_),
    .B(_11457_),
    .C(_11456_),
    .Y(_11462_)
);

OAI21X1 _21372_ (
    .A(_11453_),
    .B(_11449_),
    .C(_11447_),
    .Y(_11463_)
);

NAND3X1 _21373_ (
    .A(_11460_),
    .B(_11462_),
    .C(_11463_),
    .Y(_11464_)
);

AOI21X1 _21374_ (
    .A(_11464_),
    .B(_11459_),
    .C(_11445_),
    .Y(_11465_)
);

INVX2 _21375_ (
    .A(_11441_),
    .Y(_11466_)
);

XNOR2X1 _21376_ (
    .A(_11444_),
    .B(_11466_),
    .Y(_11467_)
);

NAND3X1 _21377_ (
    .A(_11462_),
    .B(_11446_),
    .C(_11463_),
    .Y(_11468_)
);

OAI21X1 _21378_ (
    .A(_11454_),
    .B(_11458_),
    .C(_11460_),
    .Y(_11469_)
);

AOI21X1 _21379_ (
    .A(_11468_),
    .B(_11469_),
    .C(_11467_),
    .Y(_11470_)
);

OR2X2 _21380_ (
    .A(_11470_),
    .B(_11465_),
    .Y(_11471_)
);

OAI21X1 _21381_ (
    .A(_11195_),
    .B(_11193_),
    .C(_11184_),
    .Y(_11473_)
);

AND2X2 _21382_ (
    .A(breg_16_bF$buf3),
    .B(areg_26_bF$buf3),
    .Y(_11474_)
);

AOI21X1 _21383_ (
    .A(_10856_),
    .B(_11474_),
    .C(_11185_),
    .Y(_11475_)
);

NAND2X1 _21384_ (
    .A(breg_17_bF$buf3),
    .B(areg_25_bF$buf2),
    .Y(_11476_)
);

INVX1 _21385_ (
    .A(_11476_),
    .Y(_11477_)
);

AND2X2 _21386_ (
    .A(breg_15_bF$buf5),
    .B(areg_27_bF$buf1),
    .Y(_11478_)
);

NAND2X1 _21387_ (
    .A(_11474_),
    .B(_11478_),
    .Y(_11479_)
);

NAND2X1 _21388_ (
    .A(breg_16_bF$buf2),
    .B(areg_26_bF$buf2),
    .Y(_11480_)
);

OAI21X1 _21389_ (
    .A(_2362__bF$buf3),
    .B(_7100__bF$buf2),
    .C(_11480_),
    .Y(_11481_)
);

NAND3X1 _21390_ (
    .A(_11477_),
    .B(_11481_),
    .C(_11479_),
    .Y(_11482_)
);

OAI21X1 _21391_ (
    .A(_2560__bF$buf1),
    .B(_6686__bF$buf2),
    .C(_11478_),
    .Y(_11484_)
);

OAI21X1 _21392_ (
    .A(_2362__bF$buf2),
    .B(_7100__bF$buf1),
    .C(_11474_),
    .Y(_11485_)
);

NAND3X1 _21393_ (
    .A(_11476_),
    .B(_11484_),
    .C(_11485_),
    .Y(_11486_)
);

NOR2X1 _21394_ (
    .A(_11181_),
    .B(_11230_),
    .Y(_11487_)
);

AOI21X1 _21395_ (
    .A(_11227_),
    .B(_11232_),
    .C(_11487_),
    .Y(_11488_)
);

NAND3X1 _21396_ (
    .A(_11488_),
    .B(_11482_),
    .C(_11486_),
    .Y(_11489_)
);

AOI21X1 _21397_ (
    .A(_11484_),
    .B(_11485_),
    .C(_11476_),
    .Y(_11490_)
);

AOI21X1 _21398_ (
    .A(_11481_),
    .B(_11479_),
    .C(_11477_),
    .Y(_11491_)
);

AND2X2 _21399_ (
    .A(_11181_),
    .B(_11230_),
    .Y(_11492_)
);

OAI22X1 _21400_ (
    .A(_10912_),
    .B(_11228_),
    .C(_11492_),
    .D(_11226_),
    .Y(_11493_)
);

OAI21X1 _21401_ (
    .A(_11490_),
    .B(_11491_),
    .C(_11493_),
    .Y(_11495_)
);

AOI21X1 _21402_ (
    .A(_11489_),
    .B(_11495_),
    .C(_11475_),
    .Y(_11496_)
);

OAI21X1 _21403_ (
    .A(_10861_),
    .B(_11480_),
    .C(_11177_),
    .Y(_11497_)
);

NAND3X1 _21404_ (
    .A(_11482_),
    .B(_11486_),
    .C(_11493_),
    .Y(_11498_)
);

OAI21X1 _21405_ (
    .A(_11490_),
    .B(_11491_),
    .C(_11488_),
    .Y(_11499_)
);

AOI21X1 _21406_ (
    .A(_11498_),
    .B(_11499_),
    .C(_11497_),
    .Y(_11500_)
);

OAI21X1 _21407_ (
    .A(_11496_),
    .B(_11500_),
    .C(_11473_),
    .Y(_11501_)
);

AOI21X1 _21408_ (
    .A(_11169_),
    .B(_11191_),
    .C(_11194_),
    .Y(_11502_)
);

NAND3X1 _21409_ (
    .A(_11497_),
    .B(_11498_),
    .C(_11499_),
    .Y(_11503_)
);

NAND3X1 _21410_ (
    .A(_11475_),
    .B(_11489_),
    .C(_11495_),
    .Y(_11504_)
);

NAND3X1 _21411_ (
    .A(_11503_),
    .B(_11504_),
    .C(_11502_),
    .Y(_11506_)
);

AOI21X1 _21412_ (
    .A(_11501_),
    .B(_11506_),
    .C(_11471_),
    .Y(_11507_)
);

NOR2X1 _21413_ (
    .A(_11465_),
    .B(_11470_),
    .Y(_11508_)
);

NAND3X1 _21414_ (
    .A(_11503_),
    .B(_11504_),
    .C(_11473_),
    .Y(_11509_)
);

OAI21X1 _21415_ (
    .A(_11496_),
    .B(_11500_),
    .C(_11502_),
    .Y(_11510_)
);

AOI21X1 _21416_ (
    .A(_11509_),
    .B(_11510_),
    .C(_11508_),
    .Y(_11511_)
);

NOR3X1 _21417_ (
    .A(_11251_),
    .B(_11511_),
    .C(_11507_),
    .Y(_11512_)
);

NOR3X1 _21418_ (
    .A(_11225_),
    .B(_11247_),
    .C(_11245_),
    .Y(_11513_)
);

NAND3X1 _21419_ (
    .A(_11509_),
    .B(_11510_),
    .C(_11508_),
    .Y(_11514_)
);

NAND3X1 _21420_ (
    .A(_11501_),
    .B(_11506_),
    .C(_11471_),
    .Y(_11515_)
);

AOI21X1 _21421_ (
    .A(_11514_),
    .B(_11515_),
    .C(_11513_),
    .Y(_11517_)
);

OAI21X1 _21422_ (
    .A(_11512_),
    .B(_11517_),
    .C(_11440_),
    .Y(_11518_)
);

NAND2X1 _21423_ (
    .A(_11197_),
    .B(_11205_),
    .Y(_11519_)
);

NAND3X1 _21424_ (
    .A(_11514_),
    .B(_11515_),
    .C(_11513_),
    .Y(_11520_)
);

OAI21X1 _21425_ (
    .A(_11507_),
    .B(_11511_),
    .C(_11251_),
    .Y(_11521_)
);

NAND3X1 _21426_ (
    .A(_11519_),
    .B(_11521_),
    .C(_11520_),
    .Y(_11522_)
);

INVX1 _21427_ (
    .A(_11241_),
    .Y(_11523_)
);

AOI21X1 _21428_ (
    .A(_11234_),
    .B(_11523_),
    .C(_11243_),
    .Y(_11524_)
);

NOR2X1 _21429_ (
    .A(_2379_),
    .B(_7520__bF$buf0),
    .Y(_11525_)
);

INVX2 _21430_ (
    .A(_11525_),
    .Y(_11526_)
);

NAND2X1 _21431_ (
    .A(breg_13_bF$buf3),
    .B(areg_30_bF$buf3),
    .Y(_11528_)
);

OAI21X1 _21432_ (
    .A(_2586__bF$buf4),
    .B(_8759_),
    .C(_11228_),
    .Y(_11529_)
);

OAI21X1 _21433_ (
    .A(_11230_),
    .B(_11528_),
    .C(_11529_),
    .Y(_11530_)
);

XNOR2X1 _21434_ (
    .A(_11530_),
    .B(_11526_),
    .Y(_11531_)
);

OAI21X1 _21435_ (
    .A(_10565_),
    .B(_11237_),
    .C(_11531_),
    .Y(_11532_)
);

OR2X2 _21436_ (
    .A(_10565_),
    .B(_11237_),
    .Y(_11533_)
);

OR2X2 _21437_ (
    .A(_11531_),
    .B(_11533_),
    .Y(_11534_)
);

NAND2X1 _21438_ (
    .A(_11532_),
    .B(_11534_),
    .Y(_11535_)
);

NAND2X1 _21439_ (
    .A(_11535_),
    .B(_11524_),
    .Y(_11536_)
);

OR2X2 _21440_ (
    .A(_11524_),
    .B(_11535_),
    .Y(_11537_)
);

NAND2X1 _21441_ (
    .A(_11536_),
    .B(_11537_),
    .Y(_11539_)
);

INVX1 _21442_ (
    .A(_11539_),
    .Y(_11540_)
);

NAND3X1 _21443_ (
    .A(_11522_),
    .B(_11540_),
    .C(_11518_),
    .Y(_11541_)
);

AOI21X1 _21444_ (
    .A(_11521_),
    .B(_11520_),
    .C(_11519_),
    .Y(_11542_)
);

INVX1 _21445_ (
    .A(_11522_),
    .Y(_11543_)
);

OAI21X1 _21446_ (
    .A(_11543_),
    .B(_11542_),
    .C(_11539_),
    .Y(_11544_)
);

NAND3X1 _21447_ (
    .A(_11258_),
    .B(_11541_),
    .C(_11544_),
    .Y(_11545_)
);

INVX2 _21448_ (
    .A(_11258_),
    .Y(_11546_)
);

NAND3X1 _21449_ (
    .A(_11522_),
    .B(_11539_),
    .C(_11518_),
    .Y(_11547_)
);

OAI21X1 _21450_ (
    .A(_11543_),
    .B(_11542_),
    .C(_11540_),
    .Y(_11548_)
);

NAND3X1 _21451_ (
    .A(_11547_),
    .B(_11546_),
    .C(_11548_),
    .Y(_11550_)
);

AOI21X1 _21452_ (
    .A(_11545_),
    .B(_11550_),
    .C(_11438_),
    .Y(_11551_)
);

NAND3X1 _21453_ (
    .A(_11426_),
    .B(_11432_),
    .C(_11434_),
    .Y(_11552_)
);

NAND3X1 _21454_ (
    .A(_11326_),
    .B(_11436_),
    .C(_11435_),
    .Y(_11553_)
);

NAND2X1 _21455_ (
    .A(_11553_),
    .B(_11552_),
    .Y(_11554_)
);

NAND3X1 _21456_ (
    .A(_11541_),
    .B(_11546_),
    .C(_11544_),
    .Y(_11555_)
);

NAND3X1 _21457_ (
    .A(_11258_),
    .B(_11547_),
    .C(_11548_),
    .Y(_11556_)
);

AOI21X1 _21458_ (
    .A(_11555_),
    .B(_11556_),
    .C(_11554_),
    .Y(_11557_)
);

OAI21X1 _21459_ (
    .A(_11551_),
    .B(_11557_),
    .C(_11325_),
    .Y(_11558_)
);

AOI21X1 _21460_ (
    .A(_11273_),
    .B(_11269_),
    .C(_11281_),
    .Y(_11559_)
);

NAND3X1 _21461_ (
    .A(_11555_),
    .B(_11556_),
    .C(_11554_),
    .Y(_11561_)
);

AOI21X1 _21462_ (
    .A(_11547_),
    .B(_11548_),
    .C(_11258_),
    .Y(_11562_)
);

AOI21X1 _21463_ (
    .A(_11541_),
    .B(_11544_),
    .C(_11546_),
    .Y(_11563_)
);

OAI21X1 _21464_ (
    .A(_11562_),
    .B(_11563_),
    .C(_11438_),
    .Y(_11564_)
);

NAND3X1 _21465_ (
    .A(_11564_),
    .B(_11561_),
    .C(_11559_),
    .Y(_11565_)
);

AOI21X1 _21466_ (
    .A(_11565_),
    .B(_11558_),
    .C(_11324_),
    .Y(_11566_)
);

NAND3X1 _21467_ (
    .A(_11564_),
    .B(_11561_),
    .C(_11325_),
    .Y(_11567_)
);

OAI21X1 _21468_ (
    .A(_11551_),
    .B(_11557_),
    .C(_11559_),
    .Y(_11568_)
);

AOI21X1 _21469_ (
    .A(_11567_),
    .B(_11568_),
    .C(_11323_),
    .Y(_11569_)
);

OAI21X1 _21470_ (
    .A(_11566_),
    .B(_11569_),
    .C(_11322_),
    .Y(_11570_)
);

NOR3X1 _21471_ (
    .A(_11279_),
    .B(_11274_),
    .C(_11266_),
    .Y(_11572_)
);

AOI21X1 _21472_ (
    .A(_11010_),
    .B(_11288_),
    .C(_11572_),
    .Y(_11573_)
);

NAND3X1 _21473_ (
    .A(_11323_),
    .B(_11567_),
    .C(_11568_),
    .Y(_11574_)
);

NOR3X1 _21474_ (
    .A(_11551_),
    .B(_11557_),
    .C(_11559_),
    .Y(_11575_)
);

AOI21X1 _21475_ (
    .A(_11564_),
    .B(_11561_),
    .C(_11325_),
    .Y(_11576_)
);

OAI21X1 _21476_ (
    .A(_11575_),
    .B(_11576_),
    .C(_11324_),
    .Y(_11577_)
);

NAND3X1 _21477_ (
    .A(_11574_),
    .B(_11577_),
    .C(_11573_),
    .Y(_11578_)
);

AOI21X1 _21478_ (
    .A(_11570_),
    .B(_11578_),
    .C(_11320_),
    .Y(_11579_)
);

NAND3X1 _21479_ (
    .A(_11322_),
    .B(_11574_),
    .C(_11577_),
    .Y(_11580_)
);

OAI21X1 _21480_ (
    .A(_11566_),
    .B(_11569_),
    .C(_11573_),
    .Y(_11581_)
);

AOI21X1 _21481_ (
    .A(_11581_),
    .B(_11580_),
    .C(_11319_),
    .Y(_11583_)
);

OAI21X1 _21482_ (
    .A(_11579_),
    .B(_11583_),
    .C(_11317_),
    .Y(_11584_)
);

NOR3X1 _21483_ (
    .A(_11285_),
    .B(_11289_),
    .C(_11292_),
    .Y(_11585_)
);

AOI21X1 _21484_ (
    .A(_11006_),
    .B(_11299_),
    .C(_11585_),
    .Y(_11586_)
);

NAND3X1 _21485_ (
    .A(_11319_),
    .B(_11581_),
    .C(_11580_),
    .Y(_11587_)
);

NAND3X1 _21486_ (
    .A(_11320_),
    .B(_11570_),
    .C(_11578_),
    .Y(_11588_)
);

NAND3X1 _21487_ (
    .A(_11587_),
    .B(_11588_),
    .C(_11586_),
    .Y(_11589_)
);

NAND2X1 _21488_ (
    .A(_11589_),
    .B(_11584_),
    .Y(_11590_)
);

XNOR2X1 _21489_ (
    .A(_11315_),
    .B(_11590_),
    .Y(_0_[42])
);

NAND3X1 _21490_ (
    .A(_11317_),
    .B(_11587_),
    .C(_11588_),
    .Y(_11591_)
);

INVX1 _21491_ (
    .A(_11590_),
    .Y(_11593_)
);

OAI21X1 _21492_ (
    .A(_11315_),
    .B(_11593_),
    .C(_11591_),
    .Y(_11594_)
);

AOI21X1 _21493_ (
    .A(_11574_),
    .B(_11577_),
    .C(_11322_),
    .Y(_11595_)
);

OAI21X1 _21494_ (
    .A(_11595_),
    .B(_11320_),
    .C(_11580_),
    .Y(_11596_)
);

OAI21X1 _21495_ (
    .A(_11357_),
    .B(_11328_),
    .C(_11366_),
    .Y(_11597_)
);

INVX1 _21496_ (
    .A(_11597_),
    .Y(_11598_)
);

OAI21X1 _21497_ (
    .A(_11576_),
    .B(_11324_),
    .C(_11567_),
    .Y(_11599_)
);

NAND2X1 _21498_ (
    .A(_11426_),
    .B(_11433_),
    .Y(_11600_)
);

INVX2 _21499_ (
    .A(_11600_),
    .Y(_11601_)
);

OAI21X1 _21500_ (
    .A(_11438_),
    .B(_11563_),
    .C(_11555_),
    .Y(_11602_)
);

NAND2X1 _21501_ (
    .A(_11411_),
    .B(_11419_),
    .Y(_11604_)
);

NOR2X1 _21502_ (
    .A(_10869__bF$buf1),
    .B(_7225__bF$buf2),
    .Y(_11605_)
);

INVX1 _21503_ (
    .A(_11605_),
    .Y(_11606_)
);

OAI21X1 _21504_ (
    .A(_11345_),
    .B(_11332_),
    .C(_11355_),
    .Y(_11607_)
);

NOR2X1 _21505_ (
    .A(_549__bF$buf0),
    .B(_6815__bF$buf1),
    .Y(_11608_)
);

INVX2 _21506_ (
    .A(_11608_),
    .Y(_11609_)
);

OAI21X1 _21507_ (
    .A(_11343_),
    .B(_11334_),
    .C(_11338_),
    .Y(_11610_)
);

NAND2X1 _21508_ (
    .A(areg_14_bF$buf1),
    .B(breg_29_bF$buf0),
    .Y(_11611_)
);

INVX2 _21509_ (
    .A(_11611_),
    .Y(_11612_)
);

AND2X2 _21510_ (
    .A(areg_15_bF$buf4),
    .B(breg_28_bF$buf1),
    .Y(_11613_)
);

AND2X2 _21511_ (
    .A(areg_16_bF$buf4),
    .B(breg_27_bF$buf1),
    .Y(_11615_)
);

NAND2X1 _21512_ (
    .A(_11613_),
    .B(_11615_),
    .Y(_11616_)
);

NAND2X1 _21513_ (
    .A(areg_15_bF$buf3),
    .B(breg_28_bF$buf0),
    .Y(_11617_)
);

OAI21X1 _21514_ (
    .A(_2669__bF$buf3),
    .B(_5668__bF$buf3),
    .C(_11617_),
    .Y(_11618_)
);

NAND3X1 _21515_ (
    .A(_11612_),
    .B(_11618_),
    .C(_11616_),
    .Y(_11619_)
);

NAND2X1 _21516_ (
    .A(areg_16_bF$buf3),
    .B(breg_27_bF$buf0),
    .Y(_11620_)
);

NOR2X1 _21517_ (
    .A(_11617_),
    .B(_11620_),
    .Y(_11621_)
);

NOR2X1 _21518_ (
    .A(_11613_),
    .B(_11615_),
    .Y(_11622_)
);

OAI21X1 _21519_ (
    .A(_11622_),
    .B(_11621_),
    .C(_11611_),
    .Y(_11623_)
);

AOI21X1 _21520_ (
    .A(_11619_),
    .B(_11623_),
    .C(_11610_),
    .Y(_11624_)
);

AOI21X1 _21521_ (
    .A(_11335_),
    .B(_11339_),
    .C(_11342_),
    .Y(_11626_)
);

OAI21X1 _21522_ (
    .A(_2465__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_11615_),
    .Y(_11627_)
);

OAI21X1 _21523_ (
    .A(_2669__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_11613_),
    .Y(_11628_)
);

AOI21X1 _21524_ (
    .A(_11627_),
    .B(_11628_),
    .C(_11611_),
    .Y(_11629_)
);

AOI21X1 _21525_ (
    .A(_11618_),
    .B(_11616_),
    .C(_11612_),
    .Y(_11630_)
);

NOR3X1 _21526_ (
    .A(_11630_),
    .B(_11626_),
    .C(_11629_),
    .Y(_11631_)
);

OAI21X1 _21527_ (
    .A(_11631_),
    .B(_11624_),
    .C(_11609_),
    .Y(_11632_)
);

OAI21X1 _21528_ (
    .A(_11629_),
    .B(_11630_),
    .C(_11626_),
    .Y(_11633_)
);

NAND3X1 _21529_ (
    .A(_11619_),
    .B(_11610_),
    .C(_11623_),
    .Y(_11634_)
);

NAND3X1 _21530_ (
    .A(_11608_),
    .B(_11633_),
    .C(_11634_),
    .Y(_11635_)
);

AOI21X1 _21531_ (
    .A(_11635_),
    .B(_11632_),
    .C(_11607_),
    .Y(_11637_)
);

AOI21X1 _21532_ (
    .A(_11331_),
    .B(_11354_),
    .C(_11352_),
    .Y(_11638_)
);

AOI21X1 _21533_ (
    .A(_11633_),
    .B(_11634_),
    .C(_11608_),
    .Y(_11639_)
);

NOR3X1 _21534_ (
    .A(_11624_),
    .B(_11609_),
    .C(_11631_),
    .Y(_11640_)
);

NOR3X1 _21535_ (
    .A(_11638_),
    .B(_11639_),
    .C(_11640_),
    .Y(_11641_)
);

OAI21X1 _21536_ (
    .A(_11641_),
    .B(_11637_),
    .C(_11606_),
    .Y(_11642_)
);

OAI21X1 _21537_ (
    .A(_11640_),
    .B(_11639_),
    .C(_11638_),
    .Y(_11643_)
);

NAND3X1 _21538_ (
    .A(_11607_),
    .B(_11635_),
    .C(_11632_),
    .Y(_11644_)
);

NAND3X1 _21539_ (
    .A(_11605_),
    .B(_11644_),
    .C(_11643_),
    .Y(_11645_)
);

AND2X2 _21540_ (
    .A(_11642_),
    .B(_11645_),
    .Y(_11646_)
);

OAI21X1 _21541_ (
    .A(_11409_),
    .B(_11407_),
    .C(_11400_),
    .Y(_11647_)
);

NAND2X1 _21542_ (
    .A(_11387_),
    .B(_11393_),
    .Y(_11648_)
);

OAI21X1 _21543_ (
    .A(_11372_),
    .B(_11377_),
    .C(_11380_),
    .Y(_11649_)
);

NAND2X1 _21544_ (
    .A(areg_17_bF$buf3),
    .B(breg_26_bF$buf2),
    .Y(_11650_)
);

NAND2X1 _21545_ (
    .A(areg_18_bF$buf3),
    .B(breg_25_bF$buf5),
    .Y(_11651_)
);

NAND2X1 _21546_ (
    .A(areg_19_bF$buf0),
    .B(breg_24_bF$buf0),
    .Y(_11652_)
);

NOR2X1 _21547_ (
    .A(_11651_),
    .B(_11652_),
    .Y(_11653_)
);

AOI22X1 _21548_ (
    .A(areg_18_bF$buf2),
    .B(breg_25_bF$buf4),
    .C(areg_19_bF$buf5),
    .D(breg_24_bF$buf5),
    .Y(_11654_)
);

OAI21X1 _21549_ (
    .A(_11653_),
    .B(_11654_),
    .C(_11650_),
    .Y(_11655_)
);

INVX1 _21550_ (
    .A(_11650_),
    .Y(_11656_)
);

OR2X2 _21551_ (
    .A(_11651_),
    .B(_11652_),
    .Y(_11658_)
);

INVX1 _21552_ (
    .A(_11654_),
    .Y(_11659_)
);

NAND3X1 _21553_ (
    .A(_11656_),
    .B(_11659_),
    .C(_11658_),
    .Y(_11660_)
);

NAND2X1 _21554_ (
    .A(areg_21_bF$buf2),
    .B(breg_21_bF$buf4),
    .Y(_11661_)
);

AND2X2 _21555_ (
    .A(_11135_),
    .B(_11661_),
    .Y(_11662_)
);

OAI22X1 _21556_ (
    .A(_11383_),
    .B(_11442_),
    .C(_11662_),
    .D(_11441_),
    .Y(_11663_)
);

NAND3X1 _21557_ (
    .A(_11655_),
    .B(_11660_),
    .C(_11663_),
    .Y(_11664_)
);

AOI21X1 _21558_ (
    .A(_11659_),
    .B(_11658_),
    .C(_11656_),
    .Y(_11665_)
);

NOR3X1 _21559_ (
    .A(_11650_),
    .B(_11654_),
    .C(_11653_),
    .Y(_11666_)
);

NOR2X1 _21560_ (
    .A(_11135_),
    .B(_11661_),
    .Y(_11667_)
);

AOI21X1 _21561_ (
    .A(_11466_),
    .B(_11443_),
    .C(_11667_),
    .Y(_11669_)
);

OAI21X1 _21562_ (
    .A(_11665_),
    .B(_11666_),
    .C(_11669_),
    .Y(_11670_)
);

NAND3X1 _21563_ (
    .A(_11649_),
    .B(_11664_),
    .C(_11670_),
    .Y(_11671_)
);

INVX1 _21564_ (
    .A(_11649_),
    .Y(_11672_)
);

NAND3X1 _21565_ (
    .A(_11669_),
    .B(_11655_),
    .C(_11660_),
    .Y(_11673_)
);

OAI21X1 _21566_ (
    .A(_11665_),
    .B(_11666_),
    .C(_11663_),
    .Y(_11674_)
);

NAND3X1 _21567_ (
    .A(_11672_),
    .B(_11673_),
    .C(_11674_),
    .Y(_11675_)
);

AOI21X1 _21568_ (
    .A(_11462_),
    .B(_11463_),
    .C(_11446_),
    .Y(_11676_)
);

OAI21X1 _21569_ (
    .A(_11445_),
    .B(_11676_),
    .C(_11468_),
    .Y(_11677_)
);

NAND3X1 _21570_ (
    .A(_11671_),
    .B(_11675_),
    .C(_11677_),
    .Y(_11678_)
);

AOI21X1 _21571_ (
    .A(_11673_),
    .B(_11674_),
    .C(_11672_),
    .Y(_11680_)
);

AOI21X1 _21572_ (
    .A(_11664_),
    .B(_11670_),
    .C(_11649_),
    .Y(_11681_)
);

NOR3X1 _21573_ (
    .A(_11460_),
    .B(_11458_),
    .C(_11454_),
    .Y(_11682_)
);

AOI21X1 _21574_ (
    .A(_11469_),
    .B(_11467_),
    .C(_11682_),
    .Y(_11683_)
);

OAI21X1 _21575_ (
    .A(_11680_),
    .B(_11681_),
    .C(_11683_),
    .Y(_11684_)
);

NAND3X1 _21576_ (
    .A(_11648_),
    .B(_11678_),
    .C(_11684_),
    .Y(_11685_)
);

INVX2 _21577_ (
    .A(_11648_),
    .Y(_11686_)
);

NAND3X1 _21578_ (
    .A(_11671_),
    .B(_11675_),
    .C(_11683_),
    .Y(_11687_)
);

OAI21X1 _21579_ (
    .A(_11680_),
    .B(_11681_),
    .C(_11677_),
    .Y(_11688_)
);

NAND3X1 _21580_ (
    .A(_11687_),
    .B(_11688_),
    .C(_11686_),
    .Y(_11689_)
);

NAND3X1 _21581_ (
    .A(_11685_),
    .B(_11647_),
    .C(_11689_),
    .Y(_11691_)
);

AOI21X1 _21582_ (
    .A(_11370_),
    .B(_11404_),
    .C(_11408_),
    .Y(_11692_)
);

AOI21X1 _21583_ (
    .A(_11688_),
    .B(_11687_),
    .C(_11686_),
    .Y(_11693_)
);

AOI21X1 _21584_ (
    .A(_11678_),
    .B(_11684_),
    .C(_11648_),
    .Y(_11694_)
);

OAI21X1 _21585_ (
    .A(_11693_),
    .B(_11694_),
    .C(_11692_),
    .Y(_11695_)
);

NAND3X1 _21586_ (
    .A(_11691_),
    .B(_11695_),
    .C(_11646_),
    .Y(_11696_)
);

NAND2X1 _21587_ (
    .A(_11645_),
    .B(_11642_),
    .Y(_11697_)
);

OAI21X1 _21588_ (
    .A(_11693_),
    .B(_11694_),
    .C(_11647_),
    .Y(_11698_)
);

NAND3X1 _21589_ (
    .A(_11685_),
    .B(_11692_),
    .C(_11689_),
    .Y(_11699_)
);

NAND3X1 _21590_ (
    .A(_11699_),
    .B(_11698_),
    .C(_11697_),
    .Y(_11700_)
);

OAI21X1 _21591_ (
    .A(_11517_),
    .B(_11440_),
    .C(_11520_),
    .Y(_11702_)
);

NAND3X1 _21592_ (
    .A(_11700_),
    .B(_11702_),
    .C(_11696_),
    .Y(_11703_)
);

AOI21X1 _21593_ (
    .A(_11699_),
    .B(_11698_),
    .C(_11697_),
    .Y(_11704_)
);

AOI21X1 _21594_ (
    .A(_11691_),
    .B(_11695_),
    .C(_11646_),
    .Y(_11705_)
);

AOI21X1 _21595_ (
    .A(_11519_),
    .B(_11521_),
    .C(_11512_),
    .Y(_11706_)
);

OAI21X1 _21596_ (
    .A(_11705_),
    .B(_11704_),
    .C(_11706_),
    .Y(_11707_)
);

NAND3X1 _21597_ (
    .A(_11604_),
    .B(_11703_),
    .C(_11707_),
    .Y(_11708_)
);

INVX1 _21598_ (
    .A(_11411_),
    .Y(_11709_)
);

NOR2X1 _21599_ (
    .A(_11709_),
    .B(_11427_),
    .Y(_11710_)
);

NAND3X1 _21600_ (
    .A(_11700_),
    .B(_11706_),
    .C(_11696_),
    .Y(_11711_)
);

OAI21X1 _21601_ (
    .A(_11705_),
    .B(_11704_),
    .C(_11702_),
    .Y(_11713_)
);

NAND3X1 _21602_ (
    .A(_11710_),
    .B(_11711_),
    .C(_11713_),
    .Y(_11714_)
);

NAND2X1 _21603_ (
    .A(_11714_),
    .B(_11708_),
    .Y(_11715_)
);

INVX1 _21604_ (
    .A(_11541_),
    .Y(_11716_)
);

NAND2X1 _21605_ (
    .A(_11509_),
    .B(_11514_),
    .Y(_11717_)
);

NOR2X1 _21606_ (
    .A(_11535_),
    .B(_11524_),
    .Y(_11718_)
);

NAND2X1 _21607_ (
    .A(areg_20_bF$buf0),
    .B(breg_23_bF$buf3),
    .Y(_11719_)
);

INVX2 _21608_ (
    .A(_11719_),
    .Y(_11720_)
);

NAND2X1 _21609_ (
    .A(breg_21_bF$buf3),
    .B(areg_22_bF$buf2),
    .Y(_11721_)
);

NOR2X1 _21610_ (
    .A(_11442_),
    .B(_11721_),
    .Y(_11722_)
);

AND2X2 _21611_ (
    .A(_11442_),
    .B(_11721_),
    .Y(_11724_)
);

NOR2X1 _21612_ (
    .A(_11722_),
    .B(_11724_),
    .Y(_11725_)
);

XNOR2X1 _21613_ (
    .A(_11725_),
    .B(_11720_),
    .Y(_11726_)
);

OAI21X1 _21614_ (
    .A(_11453_),
    .B(_11447_),
    .C(_11456_),
    .Y(_11727_)
);

NAND2X1 _21615_ (
    .A(breg_20_bF$buf4),
    .B(areg_23_bF$buf0),
    .Y(_11728_)
);

NAND2X1 _21616_ (
    .A(breg_19_bF$buf1),
    .B(areg_25_bF$buf1),
    .Y(_11729_)
);

NOR2X1 _21617_ (
    .A(_11448_),
    .B(_11729_),
    .Y(_11730_)
);

AND2X2 _21618_ (
    .A(breg_19_bF$buf0),
    .B(areg_24_bF$buf3),
    .Y(_11731_)
);

AND2X2 _21619_ (
    .A(breg_18_bF$buf0),
    .B(areg_25_bF$buf0),
    .Y(_11732_)
);

NOR2X1 _21620_ (
    .A(_11731_),
    .B(_11732_),
    .Y(_11733_)
);

NOR3X1 _21621_ (
    .A(_11728_),
    .B(_11730_),
    .C(_11733_),
    .Y(_11735_)
);

INVX2 _21622_ (
    .A(_11728_),
    .Y(_11736_)
);

NAND2X1 _21623_ (
    .A(_11731_),
    .B(_11732_),
    .Y(_11737_)
);

OAI22X1 _21624_ (
    .A(_3529__bF$buf0),
    .B(_6300__bF$buf3),
    .C(_3253__bF$buf3),
    .D(_5921__bF$buf0),
    .Y(_11738_)
);

AOI21X1 _21625_ (
    .A(_11738_),
    .B(_11737_),
    .C(_11736_),
    .Y(_11739_)
);

OAI21X1 _21626_ (
    .A(_11735_),
    .B(_11739_),
    .C(_11727_),
    .Y(_11740_)
);

AOI21X1 _21627_ (
    .A(_11455_),
    .B(_11457_),
    .C(_11449_),
    .Y(_11741_)
);

NAND3X1 _21628_ (
    .A(_11736_),
    .B(_11738_),
    .C(_11737_),
    .Y(_11742_)
);

OAI21X1 _21629_ (
    .A(_11733_),
    .B(_11730_),
    .C(_11728_),
    .Y(_11743_)
);

NAND3X1 _21630_ (
    .A(_11741_),
    .B(_11742_),
    .C(_11743_),
    .Y(_11744_)
);

AOI21X1 _21631_ (
    .A(_11740_),
    .B(_11744_),
    .C(_11726_),
    .Y(_11746_)
);

XNOR2X1 _21632_ (
    .A(_11725_),
    .B(_11719_),
    .Y(_11747_)
);

NAND3X1 _21633_ (
    .A(_11742_),
    .B(_11727_),
    .C(_11743_),
    .Y(_11748_)
);

OAI21X1 _21634_ (
    .A(_11735_),
    .B(_11739_),
    .C(_11741_),
    .Y(_11749_)
);

AOI21X1 _21635_ (
    .A(_11749_),
    .B(_11748_),
    .C(_11747_),
    .Y(_11750_)
);

NOR2X1 _21636_ (
    .A(_11746_),
    .B(_11750_),
    .Y(_11751_)
);

AOI21X1 _21637_ (
    .A(_11482_),
    .B(_11486_),
    .C(_11493_),
    .Y(_11752_)
);

OAI21X1 _21638_ (
    .A(_11752_),
    .B(_11475_),
    .C(_11498_),
    .Y(_11753_)
);

NAND2X1 _21639_ (
    .A(breg_15_bF$buf4),
    .B(areg_27_bF$buf0),
    .Y(_11754_)
);

OAI21X1 _21640_ (
    .A(_11480_),
    .B(_11754_),
    .C(_11482_),
    .Y(_11755_)
);

NOR2X1 _21641_ (
    .A(_2763_),
    .B(_6686__bF$buf1),
    .Y(_11757_)
);

AND2X2 _21642_ (
    .A(breg_16_bF$buf1),
    .B(areg_27_bF$buf5),
    .Y(_11758_)
);

AND2X2 _21643_ (
    .A(breg_15_bF$buf3),
    .B(areg_28_bF$buf2),
    .Y(_11759_)
);

NAND2X1 _21644_ (
    .A(_11758_),
    .B(_11759_),
    .Y(_11760_)
);

NAND2X1 _21645_ (
    .A(breg_15_bF$buf2),
    .B(areg_28_bF$buf1),
    .Y(_11761_)
);

OAI21X1 _21646_ (
    .A(_2560__bF$buf0),
    .B(_7100__bF$buf0),
    .C(_11761_),
    .Y(_11762_)
);

NAND3X1 _21647_ (
    .A(_11757_),
    .B(_11762_),
    .C(_11760_),
    .Y(_11763_)
);

NAND2X1 _21648_ (
    .A(breg_16_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_11764_)
);

OAI21X1 _21649_ (
    .A(_11754_),
    .B(_11764_),
    .C(_11762_),
    .Y(_11765_)
);

OAI21X1 _21650_ (
    .A(_2763_),
    .B(_6686__bF$buf0),
    .C(_11765_),
    .Y(_11766_)
);

AOI22X1 _21651_ (
    .A(breg_12_bF$buf3),
    .B(areg_30_bF$buf2),
    .C(breg_13_bF$buf2),
    .D(areg_29_bF$buf4),
    .Y(_11768_)
);

OAI22X1 _21652_ (
    .A(_11230_),
    .B(_11528_),
    .C(_11526_),
    .D(_11768_),
    .Y(_11769_)
);

NAND3X1 _21653_ (
    .A(_11763_),
    .B(_11769_),
    .C(_11766_),
    .Y(_11770_)
);

INVX1 _21654_ (
    .A(_11757_),
    .Y(_11771_)
);

OAI21X1 _21655_ (
    .A(_2560__bF$buf4),
    .B(_7100__bF$buf3),
    .C(_11759_),
    .Y(_11772_)
);

OAI21X1 _21656_ (
    .A(_2362__bF$buf1),
    .B(_7520__bF$buf3),
    .C(_11758_),
    .Y(_11773_)
);

AOI21X1 _21657_ (
    .A(_11772_),
    .B(_11773_),
    .C(_11771_),
    .Y(_11774_)
);

AOI21X1 _21658_ (
    .A(_11762_),
    .B(_11760_),
    .C(_11757_),
    .Y(_11775_)
);

NOR2X1 _21659_ (
    .A(_11230_),
    .B(_11528_),
    .Y(_11776_)
);

AOI21X1 _21660_ (
    .A(_11525_),
    .B(_11529_),
    .C(_11776_),
    .Y(_11777_)
);

OAI21X1 _21661_ (
    .A(_11774_),
    .B(_11775_),
    .C(_11777_),
    .Y(_11779_)
);

NAND3X1 _21662_ (
    .A(_11755_),
    .B(_11779_),
    .C(_11770_),
    .Y(_11780_)
);

INVX2 _21663_ (
    .A(_11755_),
    .Y(_11781_)
);

NOR3X1 _21664_ (
    .A(_11775_),
    .B(_11777_),
    .C(_11774_),
    .Y(_11782_)
);

AOI21X1 _21665_ (
    .A(_11763_),
    .B(_11766_),
    .C(_11769_),
    .Y(_11783_)
);

OAI21X1 _21666_ (
    .A(_11783_),
    .B(_11782_),
    .C(_11781_),
    .Y(_11784_)
);

NAND3X1 _21667_ (
    .A(_11753_),
    .B(_11780_),
    .C(_11784_),
    .Y(_11785_)
);

INVX1 _21668_ (
    .A(_11498_),
    .Y(_11786_)
);

AOI21X1 _21669_ (
    .A(_11497_),
    .B(_11499_),
    .C(_11786_),
    .Y(_11787_)
);

NAND3X1 _21670_ (
    .A(_11763_),
    .B(_11777_),
    .C(_11766_),
    .Y(_11788_)
);

OAI21X1 _21671_ (
    .A(_11774_),
    .B(_11775_),
    .C(_11769_),
    .Y(_11790_)
);

AOI21X1 _21672_ (
    .A(_11790_),
    .B(_11788_),
    .C(_11781_),
    .Y(_11791_)
);

AOI21X1 _21673_ (
    .A(_11779_),
    .B(_11770_),
    .C(_11755_),
    .Y(_11792_)
);

OAI21X1 _21674_ (
    .A(_11791_),
    .B(_11792_),
    .C(_11787_),
    .Y(_11793_)
);

NAND3X1 _21675_ (
    .A(_11751_),
    .B(_11785_),
    .C(_11793_),
    .Y(_11794_)
);

OR2X2 _21676_ (
    .A(_11746_),
    .B(_11750_),
    .Y(_11795_)
);

OAI21X1 _21677_ (
    .A(_11791_),
    .B(_11792_),
    .C(_11753_),
    .Y(_11796_)
);

NAND3X1 _21678_ (
    .A(_11780_),
    .B(_11784_),
    .C(_11787_),
    .Y(_11797_)
);

NAND3X1 _21679_ (
    .A(_11796_),
    .B(_11797_),
    .C(_11795_),
    .Y(_11798_)
);

NAND3X1 _21680_ (
    .A(_11718_),
    .B(_11794_),
    .C(_11798_),
    .Y(_11799_)
);

AOI21X1 _21681_ (
    .A(_11796_),
    .B(_11797_),
    .C(_11795_),
    .Y(_11801_)
);

AOI21X1 _21682_ (
    .A(_11785_),
    .B(_11793_),
    .C(_11751_),
    .Y(_11802_)
);

OAI21X1 _21683_ (
    .A(_11801_),
    .B(_11802_),
    .C(_11537_),
    .Y(_11803_)
);

AOI21X1 _21684_ (
    .A(_11799_),
    .B(_11803_),
    .C(_11717_),
    .Y(_11804_)
);

AND2X2 _21685_ (
    .A(_11514_),
    .B(_11509_),
    .Y(_11805_)
);

NOR3X1 _21686_ (
    .A(_11802_),
    .B(_11537_),
    .C(_11801_),
    .Y(_11806_)
);

AOI21X1 _21687_ (
    .A(_11794_),
    .B(_11798_),
    .C(_11718_),
    .Y(_11807_)
);

NOR3X1 _21688_ (
    .A(_11805_),
    .B(_11807_),
    .C(_11806_),
    .Y(_11808_)
);

NOR2X1 _21689_ (
    .A(_11533_),
    .B(_11531_),
    .Y(_11809_)
);

NOR2X1 _21690_ (
    .A(_11238_),
    .B(_11809_),
    .Y(_11810_)
);

NOR2X1 _21691_ (
    .A(_2379_),
    .B(_9153_),
    .Y(_11812_)
);

NAND2X1 _21692_ (
    .A(breg_12_bF$buf2),
    .B(areg_31_bF$buf2),
    .Y(_11813_)
);

NOR2X1 _21693_ (
    .A(_11528_),
    .B(_11813_),
    .Y(_11814_)
);

AND2X2 _21694_ (
    .A(_11528_),
    .B(_11813_),
    .Y(_11815_)
);

NOR2X1 _21695_ (
    .A(_11814_),
    .B(_11815_),
    .Y(_11816_)
);

XNOR2X1 _21696_ (
    .A(_11816_),
    .B(_11812_),
    .Y(_11817_)
);

OR2X2 _21697_ (
    .A(_11810_),
    .B(_11817_),
    .Y(_11818_)
);

NAND2X1 _21698_ (
    .A(_11817_),
    .B(_11810_),
    .Y(_11819_)
);

NAND2X1 _21699_ (
    .A(_11819_),
    .B(_11818_),
    .Y(_11820_)
);

OAI21X1 _21700_ (
    .A(_11808_),
    .B(_11804_),
    .C(_11820_),
    .Y(_11821_)
);

OAI21X1 _21701_ (
    .A(_11806_),
    .B(_11807_),
    .C(_11805_),
    .Y(_11823_)
);

NAND3X1 _21702_ (
    .A(_11717_),
    .B(_11799_),
    .C(_11803_),
    .Y(_11824_)
);

INVX1 _21703_ (
    .A(_11820_),
    .Y(_11825_)
);

NAND3X1 _21704_ (
    .A(_11824_),
    .B(_11825_),
    .C(_11823_),
    .Y(_11826_)
);

AOI21X1 _21705_ (
    .A(_11826_),
    .B(_11821_),
    .C(_11716_),
    .Y(_11827_)
);

AOI21X1 _21706_ (
    .A(_11824_),
    .B(_11823_),
    .C(_11825_),
    .Y(_11828_)
);

NOR3X1 _21707_ (
    .A(_11804_),
    .B(_11820_),
    .C(_11808_),
    .Y(_11829_)
);

NOR3X1 _21708_ (
    .A(_11541_),
    .B(_11828_),
    .C(_11829_),
    .Y(_11830_)
);

NOR3X1 _21709_ (
    .A(_11830_),
    .B(_11827_),
    .C(_11715_),
    .Y(_11831_)
);

AOI21X1 _21710_ (
    .A(_11711_),
    .B(_11713_),
    .C(_11710_),
    .Y(_11832_)
);

AOI21X1 _21711_ (
    .A(_11703_),
    .B(_11707_),
    .C(_11604_),
    .Y(_11834_)
);

NOR2X1 _21712_ (
    .A(_11832_),
    .B(_11834_),
    .Y(_11835_)
);

OAI21X1 _21713_ (
    .A(_11829_),
    .B(_11828_),
    .C(_11541_),
    .Y(_11836_)
);

NAND3X1 _21714_ (
    .A(_11826_),
    .B(_11821_),
    .C(_11716_),
    .Y(_11837_)
);

AOI21X1 _21715_ (
    .A(_11836_),
    .B(_11837_),
    .C(_11835_),
    .Y(_11838_)
);

OAI21X1 _21716_ (
    .A(_11831_),
    .B(_11838_),
    .C(_11602_),
    .Y(_11839_)
);

AOI21X1 _21717_ (
    .A(_11556_),
    .B(_11554_),
    .C(_11562_),
    .Y(_11840_)
);

NAND3X1 _21718_ (
    .A(_11836_),
    .B(_11837_),
    .C(_11835_),
    .Y(_11841_)
);

OAI21X1 _21719_ (
    .A(_11830_),
    .B(_11827_),
    .C(_11715_),
    .Y(_11842_)
);

NAND3X1 _21720_ (
    .A(_11842_),
    .B(_11840_),
    .C(_11841_),
    .Y(_11843_)
);

AOI21X1 _21721_ (
    .A(_11843_),
    .B(_11839_),
    .C(_11601_),
    .Y(_11845_)
);

NAND3X1 _21722_ (
    .A(_11842_),
    .B(_11602_),
    .C(_11841_),
    .Y(_11846_)
);

OAI21X1 _21723_ (
    .A(_11831_),
    .B(_11838_),
    .C(_11840_),
    .Y(_11847_)
);

AOI21X1 _21724_ (
    .A(_11846_),
    .B(_11847_),
    .C(_11600_),
    .Y(_11848_)
);

OAI21X1 _21725_ (
    .A(_11845_),
    .B(_11848_),
    .C(_11599_),
    .Y(_11849_)
);

AOI21X1 _21726_ (
    .A(_11323_),
    .B(_11568_),
    .C(_11575_),
    .Y(_11850_)
);

NAND3X1 _21727_ (
    .A(_11600_),
    .B(_11846_),
    .C(_11847_),
    .Y(_11851_)
);

NAND3X1 _21728_ (
    .A(_11601_),
    .B(_11843_),
    .C(_11839_),
    .Y(_11852_)
);

NAND3X1 _21729_ (
    .A(_11850_),
    .B(_11851_),
    .C(_11852_),
    .Y(_11853_)
);

AOI21X1 _21730_ (
    .A(_11853_),
    .B(_11849_),
    .C(_11598_),
    .Y(_11854_)
);

NAND3X1 _21731_ (
    .A(_11599_),
    .B(_11852_),
    .C(_11851_),
    .Y(_11856_)
);

OAI21X1 _21732_ (
    .A(_11845_),
    .B(_11848_),
    .C(_11850_),
    .Y(_11857_)
);

AOI21X1 _21733_ (
    .A(_11856_),
    .B(_11857_),
    .C(_11597_),
    .Y(_11858_)
);

OAI21X1 _21734_ (
    .A(_11854_),
    .B(_11858_),
    .C(_11596_),
    .Y(_11859_)
);

NOR3X1 _21735_ (
    .A(_11566_),
    .B(_11569_),
    .C(_11573_),
    .Y(_11860_)
);

AOI21X1 _21736_ (
    .A(_11319_),
    .B(_11581_),
    .C(_11860_),
    .Y(_11861_)
);

NAND3X1 _21737_ (
    .A(_11597_),
    .B(_11856_),
    .C(_11857_),
    .Y(_11862_)
);

NAND3X1 _21738_ (
    .A(_11598_),
    .B(_11853_),
    .C(_11849_),
    .Y(_11863_)
);

NAND3X1 _21739_ (
    .A(_11862_),
    .B(_11863_),
    .C(_11861_),
    .Y(_11864_)
);

NAND2X1 _21740_ (
    .A(_11864_),
    .B(_11859_),
    .Y(_11865_)
);

XOR2X1 _21741_ (
    .A(_11594_),
    .B(_11865_),
    .Y(_0_[43])
);

NAND2X1 _21742_ (
    .A(_11309_),
    .B(_11311_),
    .Y(_11867_)
);

NAND2X1 _21743_ (
    .A(_11590_),
    .B(_11865_),
    .Y(_11868_)
);

OAI21X1 _21744_ (
    .A(_11854_),
    .B(_11858_),
    .C(_11861_),
    .Y(_11869_)
);

NAND3X1 _21745_ (
    .A(_11862_),
    .B(_11863_),
    .C(_11596_),
    .Y(_11870_)
);

NAND2X1 _21746_ (
    .A(_11591_),
    .B(_11870_),
    .Y(_11871_)
);

NAND2X1 _21747_ (
    .A(_11869_),
    .B(_11871_),
    .Y(_11872_)
);

OAI21X1 _21748_ (
    .A(_11868_),
    .B(_11867_),
    .C(_11872_),
    .Y(_11873_)
);

AOI22X1 _21749_ (
    .A(_11584_),
    .B(_11589_),
    .C(_11859_),
    .D(_11864_),
    .Y(_11874_)
);

NAND2X1 _21750_ (
    .A(_11313_),
    .B(_11874_),
    .Y(_11875_)
);

INVX1 _21751_ (
    .A(_11875_),
    .Y(_11877_)
);

AND2X2 _21752_ (
    .A(_10688_),
    .B(_11877_),
    .Y(_11878_)
);

NOR2X1 _21753_ (
    .A(_11873_),
    .B(_11878_),
    .Y(_11879_)
);

NOR3X1 _21754_ (
    .A(_11845_),
    .B(_11850_),
    .C(_11848_),
    .Y(_11880_)
);

OAI21X1 _21755_ (
    .A(_11637_),
    .B(_11606_),
    .C(_11644_),
    .Y(_11881_)
);

INVX2 _21756_ (
    .A(_11881_),
    .Y(_11882_)
);

AOI21X1 _21757_ (
    .A(_11842_),
    .B(_11841_),
    .C(_11602_),
    .Y(_11883_)
);

OAI21X1 _21758_ (
    .A(_11883_),
    .B(_11601_),
    .C(_11846_),
    .Y(_11884_)
);

NAND2X1 _21759_ (
    .A(_11703_),
    .B(_11708_),
    .Y(_11885_)
);

INVX2 _21760_ (
    .A(_11885_),
    .Y(_11886_)
);

OAI21X1 _21761_ (
    .A(_11715_),
    .B(_11827_),
    .C(_11837_),
    .Y(_11888_)
);

NAND2X1 _21762_ (
    .A(_11691_),
    .B(_11696_),
    .Y(_11889_)
);

NOR2X1 _21763_ (
    .A(_549__bF$buf4),
    .B(_7225__bF$buf1),
    .Y(_11890_)
);

INVX1 _21764_ (
    .A(_11890_),
    .Y(_11891_)
);

OAI21X1 _21765_ (
    .A(_11624_),
    .B(_11609_),
    .C(_11634_),
    .Y(_11892_)
);

NOR2X1 _21766_ (
    .A(_2287__bF$buf3),
    .B(_6815__bF$buf0),
    .Y(_11893_)
);

INVX2 _21767_ (
    .A(_11893_),
    .Y(_11894_)
);

OAI21X1 _21768_ (
    .A(_11622_),
    .B(_11611_),
    .C(_11616_),
    .Y(_11895_)
);

NAND2X1 _21769_ (
    .A(areg_15_bF$buf2),
    .B(breg_29_bF$buf4),
    .Y(_11896_)
);

INVX2 _21770_ (
    .A(_11896_),
    .Y(_11897_)
);

AND2X2 _21771_ (
    .A(areg_16_bF$buf2),
    .B(breg_28_bF$buf5),
    .Y(_11899_)
);

AND2X2 _21772_ (
    .A(areg_17_bF$buf2),
    .B(breg_27_bF$buf5),
    .Y(_11900_)
);

NAND2X1 _21773_ (
    .A(_11899_),
    .B(_11900_),
    .Y(_11901_)
);

NAND2X1 _21774_ (
    .A(areg_16_bF$buf1),
    .B(breg_28_bF$buf4),
    .Y(_11902_)
);

OAI21X1 _21775_ (
    .A(_2884__bF$buf1),
    .B(_5668__bF$buf1),
    .C(_11902_),
    .Y(_11903_)
);

NAND3X1 _21776_ (
    .A(_11897_),
    .B(_11903_),
    .C(_11901_),
    .Y(_11904_)
);

NAND2X1 _21777_ (
    .A(areg_17_bF$buf1),
    .B(breg_27_bF$buf4),
    .Y(_11905_)
);

NOR2X1 _21778_ (
    .A(_11902_),
    .B(_11905_),
    .Y(_11906_)
);

NOR2X1 _21779_ (
    .A(_11899_),
    .B(_11900_),
    .Y(_11907_)
);

OAI21X1 _21780_ (
    .A(_11907_),
    .B(_11906_),
    .C(_11896_),
    .Y(_11908_)
);

AOI21X1 _21781_ (
    .A(_11904_),
    .B(_11908_),
    .C(_11895_),
    .Y(_2_)
);

AOI21X1 _21782_ (
    .A(_11612_),
    .B(_11618_),
    .C(_11621_),
    .Y(_3_)
);

OAI21X1 _21783_ (
    .A(_2669__bF$buf1),
    .B(_6050__bF$buf0),
    .C(_11900_),
    .Y(_4_)
);

OAI21X1 _21784_ (
    .A(_2884__bF$buf0),
    .B(_5668__bF$buf0),
    .C(_11899_),
    .Y(_5_)
);

AOI21X1 _21785_ (
    .A(_4_),
    .B(_5_),
    .C(_11896_),
    .Y(_6_)
);

AOI21X1 _21786_ (
    .A(_11903_),
    .B(_11901_),
    .C(_11897_),
    .Y(_7_)
);

NOR3X1 _21787_ (
    .A(_7_),
    .B(_3_),
    .C(_6_),
    .Y(_8_)
);

OAI21X1 _21788_ (
    .A(_8_),
    .B(_2_),
    .C(_11894_),
    .Y(_9_)
);

OAI21X1 _21789_ (
    .A(_6_),
    .B(_7_),
    .C(_3_),
    .Y(_10_)
);

NAND3X1 _21790_ (
    .A(_11904_),
    .B(_11895_),
    .C(_11908_),
    .Y(_11_)
);

NAND3X1 _21791_ (
    .A(_11893_),
    .B(_10_),
    .C(_11_),
    .Y(_13_)
);

AOI21X1 _21792_ (
    .A(_13_),
    .B(_9_),
    .C(_11892_),
    .Y(_14_)
);

AOI21X1 _21793_ (
    .A(_11608_),
    .B(_11633_),
    .C(_11631_),
    .Y(_15_)
);

AOI21X1 _21794_ (
    .A(_10_),
    .B(_11_),
    .C(_11893_),
    .Y(_16_)
);

NOR3X1 _21795_ (
    .A(_2_),
    .B(_11894_),
    .C(_8_),
    .Y(_17_)
);

NOR3X1 _21796_ (
    .A(_15_),
    .B(_16_),
    .C(_17_),
    .Y(_18_)
);

OAI21X1 _21797_ (
    .A(_18_),
    .B(_14_),
    .C(_11891_),
    .Y(_19_)
);

OAI21X1 _21798_ (
    .A(_17_),
    .B(_16_),
    .C(_15_),
    .Y(_20_)
);

NAND3X1 _21799_ (
    .A(_11892_),
    .B(_13_),
    .C(_9_),
    .Y(_21_)
);

NAND3X1 _21800_ (
    .A(_11890_),
    .B(_21_),
    .C(_20_),
    .Y(_22_)
);

AND2X2 _21801_ (
    .A(_19_),
    .B(_22_),
    .Y(_24_)
);

AOI21X1 _21802_ (
    .A(_11671_),
    .B(_11675_),
    .C(_11677_),
    .Y(_25_)
);

OAI21X1 _21803_ (
    .A(_11686_),
    .B(_25_),
    .C(_11678_),
    .Y(_26_)
);

NAND2X1 _21804_ (
    .A(_11664_),
    .B(_11671_),
    .Y(_27_)
);

OAI21X1 _21805_ (
    .A(_11650_),
    .B(_11654_),
    .C(_11658_),
    .Y(_28_)
);

NAND2X1 _21806_ (
    .A(areg_18_bF$buf1),
    .B(breg_26_bF$buf1),
    .Y(_29_)
);

NAND2X1 _21807_ (
    .A(areg_19_bF$buf4),
    .B(breg_25_bF$buf3),
    .Y(_30_)
);

NAND2X1 _21808_ (
    .A(areg_20_bF$buf4),
    .B(breg_24_bF$buf4),
    .Y(_31_)
);

NOR2X1 _21809_ (
    .A(_30_),
    .B(_31_),
    .Y(_32_)
);

AOI22X1 _21810_ (
    .A(areg_19_bF$buf3),
    .B(breg_25_bF$buf2),
    .C(areg_20_bF$buf3),
    .D(breg_24_bF$buf3),
    .Y(_33_)
);

OAI21X1 _21811_ (
    .A(_32_),
    .B(_33_),
    .C(_29_),
    .Y(_35_)
);

INVX1 _21812_ (
    .A(_29_),
    .Y(_36_)
);

OR2X2 _21813_ (
    .A(_30_),
    .B(_31_),
    .Y(_37_)
);

INVX1 _21814_ (
    .A(_33_),
    .Y(_38_)
);

NAND3X1 _21815_ (
    .A(_36_),
    .B(_38_),
    .C(_37_),
    .Y(_39_)
);

NAND2X1 _21816_ (
    .A(areg_22_bF$buf1),
    .B(breg_22_bF$buf2),
    .Y(_40_)
);

OAI22X1 _21817_ (
    .A(_11661_),
    .B(_40_),
    .C(_11724_),
    .D(_11719_),
    .Y(_41_)
);

NAND3X1 _21818_ (
    .A(_35_),
    .B(_39_),
    .C(_41_),
    .Y(_42_)
);

AOI21X1 _21819_ (
    .A(_38_),
    .B(_37_),
    .C(_36_),
    .Y(_43_)
);

NOR3X1 _21820_ (
    .A(_29_),
    .B(_33_),
    .C(_32_),
    .Y(_44_)
);

OAI21X1 _21821_ (
    .A(_3781__bF$buf3),
    .B(_4551__bF$buf3),
    .C(_11442_),
    .Y(_46_)
);

AOI21X1 _21822_ (
    .A(_11720_),
    .B(_46_),
    .C(_11722_),
    .Y(_47_)
);

OAI21X1 _21823_ (
    .A(_43_),
    .B(_44_),
    .C(_47_),
    .Y(_48_)
);

NAND3X1 _21824_ (
    .A(_28_),
    .B(_42_),
    .C(_48_),
    .Y(_49_)
);

INVX1 _21825_ (
    .A(_28_),
    .Y(_50_)
);

NAND3X1 _21826_ (
    .A(_47_),
    .B(_35_),
    .C(_39_),
    .Y(_51_)
);

OAI21X1 _21827_ (
    .A(_43_),
    .B(_44_),
    .C(_41_),
    .Y(_52_)
);

NAND3X1 _21828_ (
    .A(_50_),
    .B(_51_),
    .C(_52_),
    .Y(_53_)
);

AOI21X1 _21829_ (
    .A(_11742_),
    .B(_11743_),
    .C(_11727_),
    .Y(_54_)
);

OAI21X1 _21830_ (
    .A(_11726_),
    .B(_54_),
    .C(_11748_),
    .Y(_55_)
);

NAND3X1 _21831_ (
    .A(_49_),
    .B(_53_),
    .C(_55_),
    .Y(_57_)
);

AOI21X1 _21832_ (
    .A(_51_),
    .B(_52_),
    .C(_50_),
    .Y(_58_)
);

AOI21X1 _21833_ (
    .A(_42_),
    .B(_48_),
    .C(_28_),
    .Y(_59_)
);

NOR3X1 _21834_ (
    .A(_11741_),
    .B(_11739_),
    .C(_11735_),
    .Y(_60_)
);

AOI21X1 _21835_ (
    .A(_11749_),
    .B(_11747_),
    .C(_60_),
    .Y(_61_)
);

OAI21X1 _21836_ (
    .A(_58_),
    .B(_59_),
    .C(_61_),
    .Y(_62_)
);

NAND3X1 _21837_ (
    .A(_27_),
    .B(_62_),
    .C(_57_),
    .Y(_63_)
);

INVX2 _21838_ (
    .A(_27_),
    .Y(_64_)
);

NAND3X1 _21839_ (
    .A(_49_),
    .B(_53_),
    .C(_61_),
    .Y(_65_)
);

OAI21X1 _21840_ (
    .A(_58_),
    .B(_59_),
    .C(_55_),
    .Y(_66_)
);

NAND3X1 _21841_ (
    .A(_66_),
    .B(_65_),
    .C(_64_),
    .Y(_68_)
);

NAND3X1 _21842_ (
    .A(_63_),
    .B(_68_),
    .C(_26_),
    .Y(_69_)
);

NOR3X1 _21843_ (
    .A(_11680_),
    .B(_11681_),
    .C(_11683_),
    .Y(_70_)
);

AOI21X1 _21844_ (
    .A(_11648_),
    .B(_11684_),
    .C(_70_),
    .Y(_71_)
);

AOI21X1 _21845_ (
    .A(_66_),
    .B(_65_),
    .C(_64_),
    .Y(_72_)
);

AOI21X1 _21846_ (
    .A(_62_),
    .B(_57_),
    .C(_27_),
    .Y(_73_)
);

OAI21X1 _21847_ (
    .A(_72_),
    .B(_73_),
    .C(_71_),
    .Y(_74_)
);

NAND3X1 _21848_ (
    .A(_69_),
    .B(_74_),
    .C(_24_),
    .Y(_75_)
);

NAND2X1 _21849_ (
    .A(_22_),
    .B(_19_),
    .Y(_76_)
);

OAI21X1 _21850_ (
    .A(_72_),
    .B(_73_),
    .C(_26_),
    .Y(_77_)
);

NAND3X1 _21851_ (
    .A(_63_),
    .B(_71_),
    .C(_68_),
    .Y(_79_)
);

NAND3X1 _21852_ (
    .A(_76_),
    .B(_79_),
    .C(_77_),
    .Y(_80_)
);

OAI21X1 _21853_ (
    .A(_11807_),
    .B(_11805_),
    .C(_11799_),
    .Y(_81_)
);

NAND3X1 _21854_ (
    .A(_80_),
    .B(_81_),
    .C(_75_),
    .Y(_82_)
);

AOI21X1 _21855_ (
    .A(_79_),
    .B(_77_),
    .C(_76_),
    .Y(_83_)
);

AOI21X1 _21856_ (
    .A(_69_),
    .B(_74_),
    .C(_24_),
    .Y(_84_)
);

AOI21X1 _21857_ (
    .A(_11717_),
    .B(_11803_),
    .C(_11806_),
    .Y(_85_)
);

OAI21X1 _21858_ (
    .A(_84_),
    .B(_83_),
    .C(_85_),
    .Y(_86_)
);

NAND3X1 _21859_ (
    .A(_11889_),
    .B(_82_),
    .C(_86_),
    .Y(_87_)
);

AND2X2 _21860_ (
    .A(_11696_),
    .B(_11691_),
    .Y(_88_)
);

NAND3X1 _21861_ (
    .A(_75_),
    .B(_80_),
    .C(_85_),
    .Y(_90_)
);

OAI21X1 _21862_ (
    .A(_84_),
    .B(_83_),
    .C(_81_),
    .Y(_91_)
);

NAND3X1 _21863_ (
    .A(_91_),
    .B(_88_),
    .C(_90_),
    .Y(_92_)
);

NAND2X1 _21864_ (
    .A(_87_),
    .B(_92_),
    .Y(_93_)
);

AND2X2 _21865_ (
    .A(_11794_),
    .B(_11785_),
    .Y(_94_)
);

NAND2X1 _21866_ (
    .A(areg_21_bF$buf1),
    .B(breg_23_bF$buf2),
    .Y(_95_)
);

INVX2 _21867_ (
    .A(_95_),
    .Y(_96_)
);

NAND2X1 _21868_ (
    .A(breg_21_bF$buf2),
    .B(areg_23_bF$buf4),
    .Y(_97_)
);

NOR2X1 _21869_ (
    .A(_40_),
    .B(_97_),
    .Y(_98_)
);

AND2X2 _21870_ (
    .A(_40_),
    .B(_97_),
    .Y(_99_)
);

NOR2X1 _21871_ (
    .A(_98_),
    .B(_99_),
    .Y(_101_)
);

XNOR2X1 _21872_ (
    .A(_101_),
    .B(_96_),
    .Y(_102_)
);

OAI21X1 _21873_ (
    .A(_11733_),
    .B(_11728_),
    .C(_11737_),
    .Y(_103_)
);

NAND2X1 _21874_ (
    .A(breg_20_bF$buf3),
    .B(areg_24_bF$buf2),
    .Y(_104_)
);

NAND2X1 _21875_ (
    .A(breg_18_bF$buf5),
    .B(areg_26_bF$buf1),
    .Y(_105_)
);

NOR2X1 _21876_ (
    .A(_11729_),
    .B(_105_),
    .Y(_106_)
);

AND2X2 _21877_ (
    .A(_11729_),
    .B(_105_),
    .Y(_107_)
);

NOR3X1 _21878_ (
    .A(_104_),
    .B(_106_),
    .C(_107_),
    .Y(_108_)
);

INVX2 _21879_ (
    .A(_104_),
    .Y(_109_)
);

AND2X2 _21880_ (
    .A(breg_19_bF$buf5),
    .B(areg_26_bF$buf0),
    .Y(_110_)
);

NAND2X1 _21881_ (
    .A(_11732_),
    .B(_110_),
    .Y(_112_)
);

OAI21X1 _21882_ (
    .A(_3529__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_11729_),
    .Y(_113_)
);

AOI21X1 _21883_ (
    .A(_113_),
    .B(_112_),
    .C(_109_),
    .Y(_114_)
);

OAI21X1 _21884_ (
    .A(_108_),
    .B(_114_),
    .C(_103_),
    .Y(_115_)
);

AOI21X1 _21885_ (
    .A(_11736_),
    .B(_11738_),
    .C(_11730_),
    .Y(_116_)
);

NAND3X1 _21886_ (
    .A(_109_),
    .B(_113_),
    .C(_112_),
    .Y(_117_)
);

OAI21X1 _21887_ (
    .A(_107_),
    .B(_106_),
    .C(_104_),
    .Y(_118_)
);

NAND3X1 _21888_ (
    .A(_116_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

AOI21X1 _21889_ (
    .A(_119_),
    .B(_115_),
    .C(_102_),
    .Y(_120_)
);

XNOR2X1 _21890_ (
    .A(_101_),
    .B(_95_),
    .Y(_121_)
);

NAND3X1 _21891_ (
    .A(_117_),
    .B(_118_),
    .C(_103_),
    .Y(_123_)
);

OAI21X1 _21892_ (
    .A(_108_),
    .B(_114_),
    .C(_116_),
    .Y(_124_)
);

AOI21X1 _21893_ (
    .A(_123_),
    .B(_124_),
    .C(_121_),
    .Y(_125_)
);

OR2X2 _21894_ (
    .A(_120_),
    .B(_125_),
    .Y(_126_)
);

OAI21X1 _21895_ (
    .A(_11783_),
    .B(_11781_),
    .C(_11770_),
    .Y(_127_)
);

OAI21X1 _21896_ (
    .A(_11765_),
    .B(_11771_),
    .C(_11760_),
    .Y(_128_)
);

INVX1 _21897_ (
    .A(_128_),
    .Y(_129_)
);

NAND2X1 _21898_ (
    .A(breg_17_bF$buf2),
    .B(areg_27_bF$buf4),
    .Y(_130_)
);

NAND2X1 _21899_ (
    .A(breg_15_bF$buf1),
    .B(areg_29_bF$buf3),
    .Y(_131_)
);

AND2X2 _21900_ (
    .A(_11764_),
    .B(_131_),
    .Y(_132_)
);

NOR2X1 _21901_ (
    .A(_11764_),
    .B(_131_),
    .Y(_134_)
);

OAI21X1 _21902_ (
    .A(_132_),
    .B(_134_),
    .C(_130_),
    .Y(_135_)
);

INVX1 _21903_ (
    .A(_130_),
    .Y(_136_)
);

OAI21X1 _21904_ (
    .A(_2560__bF$buf3),
    .B(_7520__bF$buf2),
    .C(_131_),
    .Y(_137_)
);

OR2X2 _21905_ (
    .A(_11764_),
    .B(_131_),
    .Y(_138_)
);

NAND3X1 _21906_ (
    .A(_136_),
    .B(_137_),
    .C(_138_),
    .Y(_139_)
);

OAI21X1 _21907_ (
    .A(_2586__bF$buf3),
    .B(_8773_),
    .C(_11528_),
    .Y(_140_)
);

AOI21X1 _21908_ (
    .A(_11812_),
    .B(_140_),
    .C(_11814_),
    .Y(_141_)
);

NAND3X1 _21909_ (
    .A(_141_),
    .B(_135_),
    .C(_139_),
    .Y(_142_)
);

AOI21X1 _21910_ (
    .A(_137_),
    .B(_138_),
    .C(_136_),
    .Y(_143_)
);

NOR3X1 _21911_ (
    .A(_130_),
    .B(_134_),
    .C(_132_),
    .Y(_145_)
);

INVX1 _21912_ (
    .A(_11812_),
    .Y(_146_)
);

INVX1 _21913_ (
    .A(_11814_),
    .Y(_147_)
);

OAI21X1 _21914_ (
    .A(_146_),
    .B(_11815_),
    .C(_147_),
    .Y(_148_)
);

OAI21X1 _21915_ (
    .A(_145_),
    .B(_143_),
    .C(_148_),
    .Y(_149_)
);

AOI21X1 _21916_ (
    .A(_142_),
    .B(_149_),
    .C(_129_),
    .Y(_150_)
);

NAND3X1 _21917_ (
    .A(_135_),
    .B(_139_),
    .C(_148_),
    .Y(_151_)
);

OAI21X1 _21918_ (
    .A(_145_),
    .B(_143_),
    .C(_141_),
    .Y(_152_)
);

AOI21X1 _21919_ (
    .A(_152_),
    .B(_151_),
    .C(_128_),
    .Y(_153_)
);

OAI21X1 _21920_ (
    .A(_153_),
    .B(_150_),
    .C(_127_),
    .Y(_154_)
);

AOI21X1 _21921_ (
    .A(_11755_),
    .B(_11779_),
    .C(_11782_),
    .Y(_156_)
);

NAND3X1 _21922_ (
    .A(_128_),
    .B(_152_),
    .C(_151_),
    .Y(_157_)
);

NAND3X1 _21923_ (
    .A(_142_),
    .B(_149_),
    .C(_129_),
    .Y(_158_)
);

NAND3X1 _21924_ (
    .A(_157_),
    .B(_158_),
    .C(_156_),
    .Y(_159_)
);

AOI21X1 _21925_ (
    .A(_159_),
    .B(_154_),
    .C(_126_),
    .Y(_160_)
);

NOR2X1 _21926_ (
    .A(_120_),
    .B(_125_),
    .Y(_161_)
);

NAND3X1 _21927_ (
    .A(_157_),
    .B(_158_),
    .C(_127_),
    .Y(_162_)
);

OAI21X1 _21928_ (
    .A(_153_),
    .B(_150_),
    .C(_156_),
    .Y(_163_)
);

AOI21X1 _21929_ (
    .A(_163_),
    .B(_162_),
    .C(_161_),
    .Y(_164_)
);

NOR3X1 _21930_ (
    .A(_160_),
    .B(_11818_),
    .C(_164_),
    .Y(_165_)
);

NOR2X1 _21931_ (
    .A(_11817_),
    .B(_11810_),
    .Y(_167_)
);

NAND3X1 _21932_ (
    .A(_161_),
    .B(_163_),
    .C(_162_),
    .Y(_168_)
);

NAND3X1 _21933_ (
    .A(_159_),
    .B(_154_),
    .C(_126_),
    .Y(_169_)
);

AOI21X1 _21934_ (
    .A(_168_),
    .B(_169_),
    .C(_167_),
    .Y(_170_)
);

OAI21X1 _21935_ (
    .A(_165_),
    .B(_170_),
    .C(_94_),
    .Y(_171_)
);

NAND2X1 _21936_ (
    .A(_11785_),
    .B(_11794_),
    .Y(_172_)
);

NAND3X1 _21937_ (
    .A(_167_),
    .B(_168_),
    .C(_169_),
    .Y(_173_)
);

OAI21X1 _21938_ (
    .A(_164_),
    .B(_160_),
    .C(_11818_),
    .Y(_174_)
);

NAND3X1 _21939_ (
    .A(_172_),
    .B(_173_),
    .C(_174_),
    .Y(_175_)
);

NOR2X1 _21940_ (
    .A(_2379_),
    .B(_8773_),
    .Y(_176_)
);

INVX2 _21941_ (
    .A(_176_),
    .Y(_178_)
);

OAI22X1 _21942_ (
    .A(_11229_),
    .B(_8773_),
    .C(_2379_),
    .D(_8759_),
    .Y(_179_)
);

OAI21X1 _21943_ (
    .A(_178_),
    .B(_11528_),
    .C(_179_),
    .Y(_180_)
);

NAND3X1 _21944_ (
    .A(_175_),
    .B(_180_),
    .C(_171_),
    .Y(_181_)
);

AOI21X1 _21945_ (
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_182_)
);

NOR3X1 _21946_ (
    .A(_94_),
    .B(_170_),
    .C(_165_),
    .Y(_183_)
);

INVX1 _21947_ (
    .A(_180_),
    .Y(_184_)
);

OAI21X1 _21948_ (
    .A(_183_),
    .B(_182_),
    .C(_184_),
    .Y(_185_)
);

NAND2X1 _21949_ (
    .A(_181_),
    .B(_185_),
    .Y(_186_)
);

NAND2X1 _21950_ (
    .A(_11826_),
    .B(_186_),
    .Y(_187_)
);

NAND3X1 _21951_ (
    .A(_181_),
    .B(_185_),
    .C(_11829_),
    .Y(_189_)
);

AOI21X1 _21952_ (
    .A(_189_),
    .B(_187_),
    .C(_93_),
    .Y(_190_)
);

NAND3X1 _21953_ (
    .A(_82_),
    .B(_86_),
    .C(_88_),
    .Y(_191_)
);

NAND3X1 _21954_ (
    .A(_11889_),
    .B(_91_),
    .C(_90_),
    .Y(_192_)
);

NAND2X1 _21955_ (
    .A(_191_),
    .B(_192_),
    .Y(_193_)
);

NAND2X1 _21956_ (
    .A(_11829_),
    .B(_186_),
    .Y(_194_)
);

NAND3X1 _21957_ (
    .A(_181_),
    .B(_11826_),
    .C(_185_),
    .Y(_195_)
);

AOI21X1 _21958_ (
    .A(_195_),
    .B(_194_),
    .C(_193_),
    .Y(_196_)
);

OAI21X1 _21959_ (
    .A(_190_),
    .B(_196_),
    .C(_11888_),
    .Y(_197_)
);

AOI21X1 _21960_ (
    .A(_11836_),
    .B(_11835_),
    .C(_11830_),
    .Y(_198_)
);

AOI21X1 _21961_ (
    .A(_91_),
    .B(_90_),
    .C(_11889_),
    .Y(_200_)
);

AOI21X1 _21962_ (
    .A(_82_),
    .B(_86_),
    .C(_88_),
    .Y(_201_)
);

AOI21X1 _21963_ (
    .A(_181_),
    .B(_185_),
    .C(_11829_),
    .Y(_202_)
);

NAND3X1 _21964_ (
    .A(_175_),
    .B(_184_),
    .C(_171_),
    .Y(_203_)
);

OAI21X1 _21965_ (
    .A(_183_),
    .B(_182_),
    .C(_180_),
    .Y(_204_)
);

AOI21X1 _21966_ (
    .A(_203_),
    .B(_204_),
    .C(_11826_),
    .Y(_205_)
);

OAI22X1 _21967_ (
    .A(_200_),
    .B(_201_),
    .C(_202_),
    .D(_205_),
    .Y(_206_)
);

AOI21X1 _21968_ (
    .A(_91_),
    .B(_90_),
    .C(_88_),
    .Y(_207_)
);

AOI21X1 _21969_ (
    .A(_82_),
    .B(_86_),
    .C(_11889_),
    .Y(_208_)
);

AOI21X1 _21970_ (
    .A(_181_),
    .B(_185_),
    .C(_11826_),
    .Y(_209_)
);

AOI21X1 _21971_ (
    .A(_203_),
    .B(_204_),
    .C(_11829_),
    .Y(_211_)
);

OAI22X1 _21972_ (
    .A(_207_),
    .B(_208_),
    .C(_211_),
    .D(_209_),
    .Y(_212_)
);

NAND3X1 _21973_ (
    .A(_206_),
    .B(_212_),
    .C(_198_),
    .Y(_213_)
);

AOI21X1 _21974_ (
    .A(_197_),
    .B(_213_),
    .C(_11886_),
    .Y(_214_)
);

NAND3X1 _21975_ (
    .A(_206_),
    .B(_212_),
    .C(_11888_),
    .Y(_215_)
);

OAI21X1 _21976_ (
    .A(_190_),
    .B(_196_),
    .C(_198_),
    .Y(_216_)
);

AOI21X1 _21977_ (
    .A(_215_),
    .B(_216_),
    .C(_11885_),
    .Y(_217_)
);

OAI21X1 _21978_ (
    .A(_214_),
    .B(_217_),
    .C(_11884_),
    .Y(_218_)
);

NOR3X1 _21979_ (
    .A(_11838_),
    .B(_11840_),
    .C(_11831_),
    .Y(_219_)
);

AOI21X1 _21980_ (
    .A(_11600_),
    .B(_11847_),
    .C(_219_),
    .Y(_220_)
);

NAND3X1 _21981_ (
    .A(_11885_),
    .B(_215_),
    .C(_216_),
    .Y(_222_)
);

NAND3X1 _21982_ (
    .A(_11886_),
    .B(_197_),
    .C(_213_),
    .Y(_223_)
);

NAND3X1 _21983_ (
    .A(_222_),
    .B(_223_),
    .C(_220_),
    .Y(_224_)
);

AOI21X1 _21984_ (
    .A(_224_),
    .B(_218_),
    .C(_11882_),
    .Y(_225_)
);

NAND3X1 _21985_ (
    .A(_222_),
    .B(_223_),
    .C(_11884_),
    .Y(_226_)
);

OAI21X1 _21986_ (
    .A(_214_),
    .B(_217_),
    .C(_220_),
    .Y(_227_)
);

AOI21X1 _21987_ (
    .A(_226_),
    .B(_227_),
    .C(_11881_),
    .Y(_228_)
);

OAI22X1 _21988_ (
    .A(_225_),
    .B(_228_),
    .C(_11854_),
    .D(_11880_),
    .Y(_229_)
);

AOI21X1 _21989_ (
    .A(_11597_),
    .B(_11857_),
    .C(_11880_),
    .Y(_230_)
);

NAND3X1 _21990_ (
    .A(_11881_),
    .B(_226_),
    .C(_227_),
    .Y(_231_)
);

NAND3X1 _21991_ (
    .A(_11882_),
    .B(_224_),
    .C(_218_),
    .Y(_233_)
);

NAND3X1 _21992_ (
    .A(_231_),
    .B(_233_),
    .C(_230_),
    .Y(_234_)
);

NAND2X1 _21993_ (
    .A(_234_),
    .B(_229_),
    .Y(_235_)
);

XNOR2X1 _21994_ (
    .A(_11879_),
    .B(_235_),
    .Y(_0_[44])
);

NAND2X1 _21995_ (
    .A(_231_),
    .B(_233_),
    .Y(_236_)
);

OR2X2 _21996_ (
    .A(_236_),
    .B(_230_),
    .Y(_237_)
);

INVX1 _21997_ (
    .A(_235_),
    .Y(_238_)
);

OAI21X1 _21998_ (
    .A(_11879_),
    .B(_238_),
    .C(_237_),
    .Y(_239_)
);

AOI21X1 _21999_ (
    .A(_222_),
    .B(_223_),
    .C(_11884_),
    .Y(_240_)
);

OAI21X1 _22000_ (
    .A(_240_),
    .B(_11882_),
    .C(_226_),
    .Y(_241_)
);

OAI21X1 _22001_ (
    .A(_14_),
    .B(_11891_),
    .C(_21_),
    .Y(_243_)
);

INVX2 _22002_ (
    .A(_243_),
    .Y(_244_)
);

AOI21X1 _22003_ (
    .A(_206_),
    .B(_212_),
    .C(_11888_),
    .Y(_245_)
);

OAI21X1 _22004_ (
    .A(_245_),
    .B(_11886_),
    .C(_215_),
    .Y(_246_)
);

NAND2X1 _22005_ (
    .A(_82_),
    .B(_87_),
    .Y(_247_)
);

INVX2 _22006_ (
    .A(_247_),
    .Y(_248_)
);

OAI21X1 _22007_ (
    .A(_93_),
    .B(_211_),
    .C(_194_),
    .Y(_249_)
);

NAND2X1 _22008_ (
    .A(_69_),
    .B(_75_),
    .Y(_250_)
);

NOR2X1 _22009_ (
    .A(_2287__bF$buf2),
    .B(_7225__bF$buf0),
    .Y(_251_)
);

INVX1 _22010_ (
    .A(_251_),
    .Y(_252_)
);

OAI21X1 _22011_ (
    .A(_2_),
    .B(_11894_),
    .C(_11_),
    .Y(_254_)
);

NOR2X1 _22012_ (
    .A(_2465__bF$buf0),
    .B(_6815__bF$buf4),
    .Y(_255_)
);

INVX2 _22013_ (
    .A(_255_),
    .Y(_256_)
);

OAI21X1 _22014_ (
    .A(_11907_),
    .B(_11896_),
    .C(_11901_),
    .Y(_257_)
);

NAND2X1 _22015_ (
    .A(areg_16_bF$buf0),
    .B(breg_29_bF$buf3),
    .Y(_258_)
);

INVX2 _22016_ (
    .A(_258_),
    .Y(_259_)
);

AND2X2 _22017_ (
    .A(areg_17_bF$buf0),
    .B(breg_28_bF$buf3),
    .Y(_260_)
);

AND2X2 _22018_ (
    .A(areg_18_bF$buf0),
    .B(breg_27_bF$buf3),
    .Y(_261_)
);

NAND2X1 _22019_ (
    .A(_260_),
    .B(_261_),
    .Y(_262_)
);

NAND2X1 _22020_ (
    .A(areg_18_bF$buf5),
    .B(breg_27_bF$buf2),
    .Y(_263_)
);

OAI21X1 _22021_ (
    .A(_2884__bF$buf3),
    .B(_6050__bF$buf3),
    .C(_263_),
    .Y(_265_)
);

NAND3X1 _22022_ (
    .A(_259_),
    .B(_265_),
    .C(_262_),
    .Y(_266_)
);

NAND2X1 _22023_ (
    .A(areg_18_bF$buf4),
    .B(breg_28_bF$buf2),
    .Y(_267_)
);

NOR2X1 _22024_ (
    .A(_11905_),
    .B(_267_),
    .Y(_268_)
);

NOR2X1 _22025_ (
    .A(_260_),
    .B(_261_),
    .Y(_269_)
);

OAI21X1 _22026_ (
    .A(_269_),
    .B(_268_),
    .C(_258_),
    .Y(_270_)
);

AOI21X1 _22027_ (
    .A(_266_),
    .B(_270_),
    .C(_257_),
    .Y(_271_)
);

AOI21X1 _22028_ (
    .A(_11897_),
    .B(_11903_),
    .C(_11906_),
    .Y(_272_)
);

OAI21X1 _22029_ (
    .A(_2884__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_261_),
    .Y(_273_)
);

OAI21X1 _22030_ (
    .A(_3146__bF$buf3),
    .B(_5668__bF$buf5),
    .C(_260_),
    .Y(_274_)
);

AOI21X1 _22031_ (
    .A(_273_),
    .B(_274_),
    .C(_258_),
    .Y(_276_)
);

AOI21X1 _22032_ (
    .A(_265_),
    .B(_262_),
    .C(_259_),
    .Y(_277_)
);

NOR3X1 _22033_ (
    .A(_277_),
    .B(_272_),
    .C(_276_),
    .Y(_278_)
);

OAI21X1 _22034_ (
    .A(_278_),
    .B(_271_),
    .C(_256_),
    .Y(_279_)
);

OAI21X1 _22035_ (
    .A(_276_),
    .B(_277_),
    .C(_272_),
    .Y(_280_)
);

NAND3X1 _22036_ (
    .A(_266_),
    .B(_257_),
    .C(_270_),
    .Y(_281_)
);

NAND3X1 _22037_ (
    .A(_255_),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

AOI21X1 _22038_ (
    .A(_282_),
    .B(_279_),
    .C(_254_),
    .Y(_283_)
);

AOI21X1 _22039_ (
    .A(_11893_),
    .B(_10_),
    .C(_8_),
    .Y(_284_)
);

AOI21X1 _22040_ (
    .A(_280_),
    .B(_281_),
    .C(_255_),
    .Y(_285_)
);

NOR3X1 _22041_ (
    .A(_271_),
    .B(_256_),
    .C(_278_),
    .Y(_287_)
);

NOR3X1 _22042_ (
    .A(_284_),
    .B(_285_),
    .C(_287_),
    .Y(_288_)
);

OAI21X1 _22043_ (
    .A(_288_),
    .B(_283_),
    .C(_252_),
    .Y(_289_)
);

OAI21X1 _22044_ (
    .A(_287_),
    .B(_285_),
    .C(_284_),
    .Y(_290_)
);

NAND3X1 _22045_ (
    .A(_254_),
    .B(_282_),
    .C(_279_),
    .Y(_291_)
);

NAND3X1 _22046_ (
    .A(_251_),
    .B(_291_),
    .C(_290_),
    .Y(_292_)
);

AND2X2 _22047_ (
    .A(_289_),
    .B(_292_),
    .Y(_293_)
);

AOI21X1 _22048_ (
    .A(_49_),
    .B(_53_),
    .C(_55_),
    .Y(_294_)
);

OAI21X1 _22049_ (
    .A(_64_),
    .B(_294_),
    .C(_57_),
    .Y(_295_)
);

NAND2X1 _22050_ (
    .A(_42_),
    .B(_49_),
    .Y(_296_)
);

OAI21X1 _22051_ (
    .A(_29_),
    .B(_33_),
    .C(_37_),
    .Y(_298_)
);

NAND2X1 _22052_ (
    .A(areg_19_bF$buf2),
    .B(breg_26_bF$buf0),
    .Y(_299_)
);

NAND2X1 _22053_ (
    .A(areg_21_bF$buf0),
    .B(breg_25_bF$buf1),
    .Y(_300_)
);

NOR2X1 _22054_ (
    .A(_31_),
    .B(_300_),
    .Y(_301_)
);

NAND2X1 _22055_ (
    .A(areg_20_bF$buf2),
    .B(breg_25_bF$buf0),
    .Y(_302_)
);

NAND2X1 _22056_ (
    .A(areg_21_bF$buf4),
    .B(breg_24_bF$buf2),
    .Y(_303_)
);

AND2X2 _22057_ (
    .A(_302_),
    .B(_303_),
    .Y(_304_)
);

OAI21X1 _22058_ (
    .A(_304_),
    .B(_301_),
    .C(_299_),
    .Y(_305_)
);

INVX1 _22059_ (
    .A(_299_),
    .Y(_306_)
);

OR2X2 _22060_ (
    .A(_302_),
    .B(_303_),
    .Y(_307_)
);

OAI21X1 _22061_ (
    .A(_3961__bF$buf0),
    .B(_5315__bF$buf1),
    .C(_302_),
    .Y(_309_)
);

NAND3X1 _22062_ (
    .A(_306_),
    .B(_309_),
    .C(_307_),
    .Y(_310_)
);

NAND2X1 _22063_ (
    .A(breg_22_bF$buf1),
    .B(areg_23_bF$buf3),
    .Y(_311_)
);

OAI22X1 _22064_ (
    .A(_11721_),
    .B(_311_),
    .C(_99_),
    .D(_95_),
    .Y(_312_)
);

NAND3X1 _22065_ (
    .A(_305_),
    .B(_310_),
    .C(_312_),
    .Y(_313_)
);

AOI21X1 _22066_ (
    .A(_309_),
    .B(_307_),
    .C(_306_),
    .Y(_314_)
);

NOR3X1 _22067_ (
    .A(_299_),
    .B(_301_),
    .C(_304_),
    .Y(_315_)
);

OAI21X1 _22068_ (
    .A(_3781__bF$buf2),
    .B(_4541__bF$buf1),
    .C(_40_),
    .Y(_316_)
);

AOI21X1 _22069_ (
    .A(_96_),
    .B(_316_),
    .C(_98_),
    .Y(_317_)
);

OAI21X1 _22070_ (
    .A(_315_),
    .B(_314_),
    .C(_317_),
    .Y(_318_)
);

NAND3X1 _22071_ (
    .A(_298_),
    .B(_313_),
    .C(_318_),
    .Y(_320_)
);

INVX1 _22072_ (
    .A(_298_),
    .Y(_321_)
);

NAND3X1 _22073_ (
    .A(_317_),
    .B(_305_),
    .C(_310_),
    .Y(_322_)
);

OAI21X1 _22074_ (
    .A(_315_),
    .B(_314_),
    .C(_312_),
    .Y(_323_)
);

NAND3X1 _22075_ (
    .A(_321_),
    .B(_322_),
    .C(_323_),
    .Y(_324_)
);

AOI21X1 _22076_ (
    .A(_117_),
    .B(_118_),
    .C(_103_),
    .Y(_325_)
);

OAI21X1 _22077_ (
    .A(_102_),
    .B(_325_),
    .C(_123_),
    .Y(_326_)
);

NAND3X1 _22078_ (
    .A(_320_),
    .B(_324_),
    .C(_326_),
    .Y(_327_)
);

AOI21X1 _22079_ (
    .A(_322_),
    .B(_323_),
    .C(_321_),
    .Y(_328_)
);

AOI21X1 _22080_ (
    .A(_313_),
    .B(_318_),
    .C(_298_),
    .Y(_329_)
);

NAND2X1 _22081_ (
    .A(_117_),
    .B(_118_),
    .Y(_331_)
);

NOR2X1 _22082_ (
    .A(_116_),
    .B(_331_),
    .Y(_332_)
);

AOI21X1 _22083_ (
    .A(_121_),
    .B(_124_),
    .C(_332_),
    .Y(_333_)
);

OAI21X1 _22084_ (
    .A(_328_),
    .B(_329_),
    .C(_333_),
    .Y(_334_)
);

NAND3X1 _22085_ (
    .A(_296_),
    .B(_334_),
    .C(_327_),
    .Y(_335_)
);

INVX2 _22086_ (
    .A(_296_),
    .Y(_336_)
);

NAND3X1 _22087_ (
    .A(_320_),
    .B(_324_),
    .C(_333_),
    .Y(_337_)
);

OAI21X1 _22088_ (
    .A(_328_),
    .B(_329_),
    .C(_326_),
    .Y(_338_)
);

NAND3X1 _22089_ (
    .A(_338_),
    .B(_336_),
    .C(_337_),
    .Y(_339_)
);

NAND3X1 _22090_ (
    .A(_335_),
    .B(_295_),
    .C(_339_),
    .Y(_340_)
);

NAND2X1 _22091_ (
    .A(_49_),
    .B(_53_),
    .Y(_342_)
);

NOR2X1 _22092_ (
    .A(_61_),
    .B(_342_),
    .Y(_343_)
);

AOI21X1 _22093_ (
    .A(_27_),
    .B(_62_),
    .C(_343_),
    .Y(_344_)
);

AOI21X1 _22094_ (
    .A(_338_),
    .B(_337_),
    .C(_336_),
    .Y(_345_)
);

AOI21X1 _22095_ (
    .A(_334_),
    .B(_327_),
    .C(_296_),
    .Y(_346_)
);

OAI21X1 _22096_ (
    .A(_345_),
    .B(_346_),
    .C(_344_),
    .Y(_347_)
);

NAND3X1 _22097_ (
    .A(_340_),
    .B(_347_),
    .C(_293_),
    .Y(_348_)
);

NAND2X1 _22098_ (
    .A(_292_),
    .B(_289_),
    .Y(_349_)
);

OAI21X1 _22099_ (
    .A(_345_),
    .B(_346_),
    .C(_295_),
    .Y(_350_)
);

NAND3X1 _22100_ (
    .A(_335_),
    .B(_339_),
    .C(_344_),
    .Y(_351_)
);

NAND3X1 _22101_ (
    .A(_349_),
    .B(_350_),
    .C(_351_),
    .Y(_353_)
);

OAI21X1 _22102_ (
    .A(_170_),
    .B(_94_),
    .C(_173_),
    .Y(_354_)
);

NAND3X1 _22103_ (
    .A(_354_),
    .B(_348_),
    .C(_353_),
    .Y(_355_)
);

AOI21X1 _22104_ (
    .A(_350_),
    .B(_351_),
    .C(_349_),
    .Y(_356_)
);

AOI21X1 _22105_ (
    .A(_340_),
    .B(_347_),
    .C(_293_),
    .Y(_357_)
);

AOI21X1 _22106_ (
    .A(_172_),
    .B(_174_),
    .C(_165_),
    .Y(_358_)
);

OAI21X1 _22107_ (
    .A(_356_),
    .B(_357_),
    .C(_358_),
    .Y(_359_)
);

NAND3X1 _22108_ (
    .A(_250_),
    .B(_355_),
    .C(_359_),
    .Y(_360_)
);

AND2X2 _22109_ (
    .A(_75_),
    .B(_69_),
    .Y(_361_)
);

NAND3X1 _22110_ (
    .A(_348_),
    .B(_353_),
    .C(_358_),
    .Y(_362_)
);

OAI21X1 _22111_ (
    .A(_356_),
    .B(_357_),
    .C(_354_),
    .Y(_363_)
);

NAND3X1 _22112_ (
    .A(_361_),
    .B(_362_),
    .C(_363_),
    .Y(_364_)
);

NAND2X1 _22113_ (
    .A(_360_),
    .B(_364_),
    .Y(_365_)
);

NAND2X1 _22114_ (
    .A(_162_),
    .B(_168_),
    .Y(_366_)
);

NOR2X1 _22115_ (
    .A(_4551__bF$buf2),
    .B(_5369_),
    .Y(_367_)
);

NAND2X1 _22116_ (
    .A(breg_21_bF$buf1),
    .B(areg_24_bF$buf1),
    .Y(_368_)
);

NOR2X1 _22117_ (
    .A(_311_),
    .B(_368_),
    .Y(_369_)
);

AND2X2 _22118_ (
    .A(_311_),
    .B(_368_),
    .Y(_370_)
);

NOR2X1 _22119_ (
    .A(_369_),
    .B(_370_),
    .Y(_371_)
);

XNOR2X1 _22120_ (
    .A(_371_),
    .B(_367_),
    .Y(_372_)
);

AOI21X1 _22121_ (
    .A(_109_),
    .B(_113_),
    .C(_106_),
    .Y(_375_)
);

NOR2X1 _22122_ (
    .A(_3526_),
    .B(_6300__bF$buf2),
    .Y(_376_)
);

INVX1 _22123_ (
    .A(_376_),
    .Y(_377_)
);

NAND2X1 _22124_ (
    .A(breg_19_bF$buf4),
    .B(areg_27_bF$buf3),
    .Y(_378_)
);

NAND2X1 _22125_ (
    .A(breg_19_bF$buf3),
    .B(areg_26_bF$buf4),
    .Y(_379_)
);

OAI21X1 _22126_ (
    .A(_3529__bF$buf3),
    .B(_7100__bF$buf2),
    .C(_379_),
    .Y(_380_)
);

OAI21X1 _22127_ (
    .A(_105_),
    .B(_378_),
    .C(_380_),
    .Y(_381_)
);

NOR2X1 _22128_ (
    .A(_377_),
    .B(_381_),
    .Y(_382_)
);

NAND2X1 _22129_ (
    .A(breg_18_bF$buf4),
    .B(areg_27_bF$buf2),
    .Y(_383_)
);

OR2X2 _22130_ (
    .A(_379_),
    .B(_383_),
    .Y(_384_)
);

AOI21X1 _22131_ (
    .A(_380_),
    .B(_384_),
    .C(_376_),
    .Y(_386_)
);

NOR3X1 _22132_ (
    .A(_375_),
    .B(_386_),
    .C(_382_),
    .Y(_387_)
);

INVX1 _22133_ (
    .A(_375_),
    .Y(_388_)
);

NAND3X1 _22134_ (
    .A(_376_),
    .B(_380_),
    .C(_384_),
    .Y(_389_)
);

OAI21X1 _22135_ (
    .A(_3526_),
    .B(_6300__bF$buf1),
    .C(_381_),
    .Y(_390_)
);

AOI21X1 _22136_ (
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_391_)
);

NOR3X1 _22137_ (
    .A(_391_),
    .B(_372_),
    .C(_387_),
    .Y(_392_)
);

INVX1 _22138_ (
    .A(_367_),
    .Y(_393_)
);

XNOR2X1 _22139_ (
    .A(_371_),
    .B(_393_),
    .Y(_394_)
);

NAND3X1 _22140_ (
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_395_)
);

OAI21X1 _22141_ (
    .A(_382_),
    .B(_386_),
    .C(_375_),
    .Y(_397_)
);

AOI21X1 _22142_ (
    .A(_395_),
    .B(_397_),
    .C(_394_),
    .Y(_398_)
);

NOR2X1 _22143_ (
    .A(_398_),
    .B(_392_),
    .Y(_399_)
);

INVX1 _22144_ (
    .A(_151_),
    .Y(_400_)
);

AOI21X1 _22145_ (
    .A(_128_),
    .B(_152_),
    .C(_400_),
    .Y(_401_)
);

OAI21X1 _22146_ (
    .A(_132_),
    .B(_130_),
    .C(_138_),
    .Y(_402_)
);

NOR2X1 _22147_ (
    .A(_11528_),
    .B(_178_),
    .Y(_403_)
);

NAND2X1 _22148_ (
    .A(breg_17_bF$buf1),
    .B(areg_28_bF$buf5),
    .Y(_404_)
);

NAND2X1 _22149_ (
    .A(breg_16_bF$buf5),
    .B(areg_30_bF$buf1),
    .Y(_405_)
);

NOR2X1 _22150_ (
    .A(_131_),
    .B(_405_),
    .Y(_406_)
);

AOI22X1 _22151_ (
    .A(breg_15_bF$buf0),
    .B(areg_30_bF$buf0),
    .C(breg_16_bF$buf4),
    .D(areg_29_bF$buf2),
    .Y(_408_)
);

OAI21X1 _22152_ (
    .A(_406_),
    .B(_408_),
    .C(_404_),
    .Y(_409_)
);

NOR3X1 _22153_ (
    .A(_404_),
    .B(_408_),
    .C(_406_),
    .Y(_410_)
);

INVX1 _22154_ (
    .A(_410_),
    .Y(_411_)
);

NAND3X1 _22155_ (
    .A(_403_),
    .B(_409_),
    .C(_411_),
    .Y(_412_)
);

OR2X2 _22156_ (
    .A(_178_),
    .B(_11528_),
    .Y(_413_)
);

INVX1 _22157_ (
    .A(_409_),
    .Y(_414_)
);

OAI21X1 _22158_ (
    .A(_414_),
    .B(_410_),
    .C(_413_),
    .Y(_415_)
);

AOI21X1 _22159_ (
    .A(_415_),
    .B(_412_),
    .C(_402_),
    .Y(_416_)
);

INVX2 _22160_ (
    .A(_402_),
    .Y(_417_)
);

NOR3X1 _22161_ (
    .A(_413_),
    .B(_410_),
    .C(_414_),
    .Y(_419_)
);

AOI21X1 _22162_ (
    .A(_409_),
    .B(_411_),
    .C(_403_),
    .Y(_420_)
);

NOR3X1 _22163_ (
    .A(_420_),
    .B(_417_),
    .C(_419_),
    .Y(_421_)
);

OAI21X1 _22164_ (
    .A(_421_),
    .B(_416_),
    .C(_401_),
    .Y(_422_)
);

NAND2X1 _22165_ (
    .A(_151_),
    .B(_157_),
    .Y(_423_)
);

OAI21X1 _22166_ (
    .A(_419_),
    .B(_420_),
    .C(_417_),
    .Y(_424_)
);

NAND3X1 _22167_ (
    .A(_402_),
    .B(_415_),
    .C(_412_),
    .Y(_425_)
);

NAND3X1 _22168_ (
    .A(_424_),
    .B(_425_),
    .C(_423_),
    .Y(_426_)
);

NAND3X1 _22169_ (
    .A(_399_),
    .B(_426_),
    .C(_422_),
    .Y(_427_)
);

OR2X2 _22170_ (
    .A(_392_),
    .B(_398_),
    .Y(_428_)
);

AOI21X1 _22171_ (
    .A(_425_),
    .B(_424_),
    .C(_423_),
    .Y(_430_)
);

NOR3X1 _22172_ (
    .A(_401_),
    .B(_416_),
    .C(_421_),
    .Y(_431_)
);

OAI21X1 _22173_ (
    .A(_431_),
    .B(_430_),
    .C(_428_),
    .Y(_432_)
);

NAND3X1 _22174_ (
    .A(_427_),
    .B(_432_),
    .C(_366_),
    .Y(_433_)
);

INVX1 _22175_ (
    .A(_162_),
    .Y(_434_)
);

AOI21X1 _22176_ (
    .A(_163_),
    .B(_161_),
    .C(_434_),
    .Y(_435_)
);

OAI21X1 _22177_ (
    .A(_431_),
    .B(_430_),
    .C(_399_),
    .Y(_436_)
);

NAND3X1 _22178_ (
    .A(_426_),
    .B(_428_),
    .C(_422_),
    .Y(_437_)
);

NAND3X1 _22179_ (
    .A(_437_),
    .B(_435_),
    .C(_436_),
    .Y(_438_)
);

NAND3X1 _22180_ (
    .A(_176_),
    .B(_438_),
    .C(_433_),
    .Y(_439_)
);

AOI21X1 _22181_ (
    .A(_437_),
    .B(_436_),
    .C(_435_),
    .Y(_441_)
);

AOI21X1 _22182_ (
    .A(_427_),
    .B(_432_),
    .C(_366_),
    .Y(_442_)
);

OAI21X1 _22183_ (
    .A(_441_),
    .B(_442_),
    .C(_178_),
    .Y(_443_)
);

NAND2X1 _22184_ (
    .A(_439_),
    .B(_443_),
    .Y(_444_)
);

XNOR2X1 _22185_ (
    .A(_444_),
    .B(_203_),
    .Y(_445_)
);

NOR2X1 _22186_ (
    .A(_365_),
    .B(_445_),
    .Y(_446_)
);

NAND2X1 _22187_ (
    .A(_203_),
    .B(_444_),
    .Y(_447_)
);

OR2X2 _22188_ (
    .A(_444_),
    .B(_203_),
    .Y(_448_)
);

AOI22X1 _22189_ (
    .A(_360_),
    .B(_364_),
    .C(_448_),
    .D(_447_),
    .Y(_449_)
);

OAI21X1 _22190_ (
    .A(_446_),
    .B(_449_),
    .C(_249_),
    .Y(_450_)
);

AOI21X1 _22191_ (
    .A(_195_),
    .B(_193_),
    .C(_209_),
    .Y(_452_)
);

AOI21X1 _22192_ (
    .A(_362_),
    .B(_363_),
    .C(_361_),
    .Y(_453_)
);

AOI21X1 _22193_ (
    .A(_355_),
    .B(_359_),
    .C(_250_),
    .Y(_454_)
);

NOR2X1 _22194_ (
    .A(_453_),
    .B(_454_),
    .Y(_455_)
);

XOR2X1 _22195_ (
    .A(_444_),
    .B(_203_),
    .Y(_456_)
);

NAND2X1 _22196_ (
    .A(_456_),
    .B(_455_),
    .Y(_457_)
);

OAI21X1 _22197_ (
    .A(_453_),
    .B(_454_),
    .C(_445_),
    .Y(_458_)
);

NAND3X1 _22198_ (
    .A(_458_),
    .B(_457_),
    .C(_452_),
    .Y(_459_)
);

AOI21X1 _22199_ (
    .A(_459_),
    .B(_450_),
    .C(_248_),
    .Y(_460_)
);

NAND3X1 _22200_ (
    .A(_458_),
    .B(_457_),
    .C(_249_),
    .Y(_461_)
);

OAI21X1 _22201_ (
    .A(_446_),
    .B(_449_),
    .C(_452_),
    .Y(_463_)
);

AOI21X1 _22202_ (
    .A(_461_),
    .B(_463_),
    .C(_247_),
    .Y(_464_)
);

OAI21X1 _22203_ (
    .A(_460_),
    .B(_464_),
    .C(_246_),
    .Y(_465_)
);

NAND2X1 _22204_ (
    .A(_206_),
    .B(_212_),
    .Y(_466_)
);

NOR2X1 _22205_ (
    .A(_198_),
    .B(_466_),
    .Y(_467_)
);

AOI21X1 _22206_ (
    .A(_11885_),
    .B(_216_),
    .C(_467_),
    .Y(_468_)
);

NAND3X1 _22207_ (
    .A(_247_),
    .B(_461_),
    .C(_463_),
    .Y(_469_)
);

NAND3X1 _22208_ (
    .A(_248_),
    .B(_459_),
    .C(_450_),
    .Y(_470_)
);

NAND3X1 _22209_ (
    .A(_469_),
    .B(_470_),
    .C(_468_),
    .Y(_471_)
);

AOI21X1 _22210_ (
    .A(_465_),
    .B(_471_),
    .C(_244_),
    .Y(_472_)
);

NAND3X1 _22211_ (
    .A(_246_),
    .B(_469_),
    .C(_470_),
    .Y(_474_)
);

OAI21X1 _22212_ (
    .A(_460_),
    .B(_464_),
    .C(_468_),
    .Y(_475_)
);

AOI21X1 _22213_ (
    .A(_474_),
    .B(_475_),
    .C(_243_),
    .Y(_476_)
);

OAI21X1 _22214_ (
    .A(_472_),
    .B(_476_),
    .C(_241_),
    .Y(_477_)
);

NOR3X1 _22215_ (
    .A(_214_),
    .B(_217_),
    .C(_220_),
    .Y(_478_)
);

AOI21X1 _22216_ (
    .A(_11881_),
    .B(_227_),
    .C(_478_),
    .Y(_479_)
);

NAND3X1 _22217_ (
    .A(_243_),
    .B(_474_),
    .C(_475_),
    .Y(_480_)
);

NAND3X1 _22218_ (
    .A(_244_),
    .B(_465_),
    .C(_471_),
    .Y(_481_)
);

NAND3X1 _22219_ (
    .A(_480_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

NAND2X1 _22220_ (
    .A(_482_),
    .B(_477_),
    .Y(_483_)
);

XOR2X1 _22221_ (
    .A(_239_),
    .B(_483_),
    .Y(_0_[45])
);

NOR2X1 _22222_ (
    .A(_230_),
    .B(_236_),
    .Y(_485_)
);

NOR3X1 _22223_ (
    .A(_472_),
    .B(_476_),
    .C(_479_),
    .Y(_486_)
);

OAI21X1 _22224_ (
    .A(_472_),
    .B(_476_),
    .C(_479_),
    .Y(_487_)
);

AOI21X1 _22225_ (
    .A(_487_),
    .B(_485_),
    .C(_486_),
    .Y(_488_)
);

AOI22X1 _22226_ (
    .A(_477_),
    .B(_482_),
    .C(_229_),
    .D(_234_),
    .Y(_489_)
);

OAI21X1 _22227_ (
    .A(_11878_),
    .B(_11873_),
    .C(_489_),
    .Y(_490_)
);

AOI21X1 _22228_ (
    .A(_469_),
    .B(_470_),
    .C(_246_),
    .Y(_491_)
);

OAI21X1 _22229_ (
    .A(_491_),
    .B(_244_),
    .C(_474_),
    .Y(_492_)
);

OAI21X1 _22230_ (
    .A(_283_),
    .B(_252_),
    .C(_291_),
    .Y(_493_)
);

INVX2 _22231_ (
    .A(_493_),
    .Y(_495_)
);

AOI21X1 _22232_ (
    .A(_458_),
    .B(_457_),
    .C(_249_),
    .Y(_496_)
);

OAI21X1 _22233_ (
    .A(_496_),
    .B(_248_),
    .C(_461_),
    .Y(_497_)
);

NAND2X1 _22234_ (
    .A(_355_),
    .B(_360_),
    .Y(_498_)
);

INVX2 _22235_ (
    .A(_498_),
    .Y(_499_)
);

OAI21X1 _22236_ (
    .A(_445_),
    .B(_365_),
    .C(_448_),
    .Y(_500_)
);

AND2X2 _22237_ (
    .A(_348_),
    .B(_340_),
    .Y(_501_)
);

NOR2X1 _22238_ (
    .A(_2465__bF$buf4),
    .B(_7225__bF$buf4),
    .Y(_502_)
);

INVX1 _22239_ (
    .A(_502_),
    .Y(_503_)
);

OAI21X1 _22240_ (
    .A(_271_),
    .B(_256_),
    .C(_281_),
    .Y(_504_)
);

NOR2X1 _22241_ (
    .A(_2669__bF$buf0),
    .B(_6815__bF$buf3),
    .Y(_506_)
);

INVX2 _22242_ (
    .A(_506_),
    .Y(_507_)
);

OAI21X1 _22243_ (
    .A(_269_),
    .B(_258_),
    .C(_262_),
    .Y(_508_)
);

NAND2X1 _22244_ (
    .A(areg_17_bF$buf5),
    .B(breg_29_bF$buf2),
    .Y(_509_)
);

NAND2X1 _22245_ (
    .A(areg_19_bF$buf1),
    .B(breg_28_bF$buf1),
    .Y(_510_)
);

NOR2X1 _22246_ (
    .A(_263_),
    .B(_510_),
    .Y(_511_)
);

NAND2X1 _22247_ (
    .A(areg_19_bF$buf0),
    .B(breg_27_bF$buf1),
    .Y(_512_)
);

AND2X2 _22248_ (
    .A(_267_),
    .B(_512_),
    .Y(_513_)
);

OAI21X1 _22249_ (
    .A(_513_),
    .B(_511_),
    .C(_509_),
    .Y(_514_)
);

INVX1 _22250_ (
    .A(_509_),
    .Y(_515_)
);

OR2X2 _22251_ (
    .A(_267_),
    .B(_512_),
    .Y(_517_)
);

OAI21X1 _22252_ (
    .A(_3402__bF$buf2),
    .B(_5668__bF$buf4),
    .C(_267_),
    .Y(_518_)
);

NAND3X1 _22253_ (
    .A(_515_),
    .B(_518_),
    .C(_517_),
    .Y(_519_)
);

AOI21X1 _22254_ (
    .A(_514_),
    .B(_519_),
    .C(_508_),
    .Y(_520_)
);

AOI21X1 _22255_ (
    .A(_259_),
    .B(_265_),
    .C(_268_),
    .Y(_521_)
);

AOI21X1 _22256_ (
    .A(_518_),
    .B(_517_),
    .C(_515_),
    .Y(_522_)
);

NOR3X1 _22257_ (
    .A(_509_),
    .B(_511_),
    .C(_513_),
    .Y(_523_)
);

NOR3X1 _22258_ (
    .A(_522_),
    .B(_521_),
    .C(_523_),
    .Y(_524_)
);

OAI21X1 _22259_ (
    .A(_524_),
    .B(_520_),
    .C(_507_),
    .Y(_525_)
);

OAI21X1 _22260_ (
    .A(_523_),
    .B(_522_),
    .C(_521_),
    .Y(_526_)
);

NAND3X1 _22261_ (
    .A(_514_),
    .B(_519_),
    .C(_508_),
    .Y(_528_)
);

NAND3X1 _22262_ (
    .A(_506_),
    .B(_528_),
    .C(_526_),
    .Y(_529_)
);

AOI21X1 _22263_ (
    .A(_529_),
    .B(_525_),
    .C(_504_),
    .Y(_530_)
);

AOI21X1 _22264_ (
    .A(_255_),
    .B(_280_),
    .C(_278_),
    .Y(_531_)
);

AOI21X1 _22265_ (
    .A(_528_),
    .B(_526_),
    .C(_506_),
    .Y(_532_)
);

NOR3X1 _22266_ (
    .A(_507_),
    .B(_520_),
    .C(_524_),
    .Y(_533_)
);

NOR3X1 _22267_ (
    .A(_531_),
    .B(_532_),
    .C(_533_),
    .Y(_534_)
);

OAI21X1 _22268_ (
    .A(_534_),
    .B(_530_),
    .C(_503_),
    .Y(_535_)
);

OAI21X1 _22269_ (
    .A(_533_),
    .B(_532_),
    .C(_531_),
    .Y(_536_)
);

NAND3X1 _22270_ (
    .A(_504_),
    .B(_529_),
    .C(_525_),
    .Y(_537_)
);

NAND3X1 _22271_ (
    .A(_502_),
    .B(_537_),
    .C(_536_),
    .Y(_539_)
);

AND2X2 _22272_ (
    .A(_535_),
    .B(_539_),
    .Y(_540_)
);

AOI21X1 _22273_ (
    .A(_320_),
    .B(_324_),
    .C(_326_),
    .Y(_541_)
);

OAI21X1 _22274_ (
    .A(_336_),
    .B(_541_),
    .C(_327_),
    .Y(_542_)
);

NAND2X1 _22275_ (
    .A(_313_),
    .B(_320_),
    .Y(_543_)
);

OAI21X1 _22276_ (
    .A(_304_),
    .B(_299_),
    .C(_307_),
    .Y(_544_)
);

NOR2X1 _22277_ (
    .A(_3958__bF$buf0),
    .B(_5676_),
    .Y(_545_)
);

INVX1 _22278_ (
    .A(_300_),
    .Y(_546_)
);

NAND2X1 _22279_ (
    .A(areg_22_bF$buf0),
    .B(breg_24_bF$buf1),
    .Y(_547_)
);

INVX1 _22280_ (
    .A(_547_),
    .Y(_548_)
);

NAND2X1 _22281_ (
    .A(_546_),
    .B(_548_),
    .Y(_550_)
);

OAI21X1 _22282_ (
    .A(_4551__bF$buf1),
    .B(_5315__bF$buf0),
    .C(_300_),
    .Y(_551_)
);

NAND3X1 _22283_ (
    .A(_545_),
    .B(_551_),
    .C(_550_),
    .Y(_552_)
);

NAND2X1 _22284_ (
    .A(areg_22_bF$buf4),
    .B(breg_25_bF$buf5),
    .Y(_553_)
);

OAI21X1 _22285_ (
    .A(_303_),
    .B(_553_),
    .C(_551_),
    .Y(_554_)
);

OAI21X1 _22286_ (
    .A(_3958__bF$buf3),
    .B(_5676_),
    .C(_554_),
    .Y(_555_)
);

OAI21X1 _22287_ (
    .A(_3781__bF$buf1),
    .B(_5921__bF$buf3),
    .C(_311_),
    .Y(_556_)
);

AOI21X1 _22288_ (
    .A(_367_),
    .B(_556_),
    .C(_369_),
    .Y(_557_)
);

INVX1 _22289_ (
    .A(_557_),
    .Y(_558_)
);

NAND3X1 _22290_ (
    .A(_552_),
    .B(_555_),
    .C(_558_),
    .Y(_559_)
);

INVX1 _22291_ (
    .A(_545_),
    .Y(_561_)
);

OAI21X1 _22292_ (
    .A(_3961__bF$buf4),
    .B(_5318_),
    .C(_548_),
    .Y(_562_)
);

OAI21X1 _22293_ (
    .A(_4551__bF$buf0),
    .B(_5315__bF$buf4),
    .C(_546_),
    .Y(_563_)
);

AOI21X1 _22294_ (
    .A(_562_),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

AOI21X1 _22295_ (
    .A(_551_),
    .B(_550_),
    .C(_545_),
    .Y(_565_)
);

OAI21X1 _22296_ (
    .A(_564_),
    .B(_565_),
    .C(_557_),
    .Y(_566_)
);

NAND3X1 _22297_ (
    .A(_544_),
    .B(_559_),
    .C(_566_),
    .Y(_567_)
);

INVX1 _22298_ (
    .A(_544_),
    .Y(_568_)
);

NAND3X1 _22299_ (
    .A(_552_),
    .B(_557_),
    .C(_555_),
    .Y(_569_)
);

OAI21X1 _22300_ (
    .A(_564_),
    .B(_565_),
    .C(_558_),
    .Y(_570_)
);

NAND3X1 _22301_ (
    .A(_568_),
    .B(_569_),
    .C(_570_),
    .Y(_572_)
);

OAI21X1 _22302_ (
    .A(_391_),
    .B(_372_),
    .C(_395_),
    .Y(_573_)
);

NAND3X1 _22303_ (
    .A(_567_),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

AOI21X1 _22304_ (
    .A(_569_),
    .B(_570_),
    .C(_568_),
    .Y(_575_)
);

AOI21X1 _22305_ (
    .A(_559_),
    .B(_566_),
    .C(_544_),
    .Y(_576_)
);

AOI21X1 _22306_ (
    .A(_394_),
    .B(_397_),
    .C(_387_),
    .Y(_577_)
);

OAI21X1 _22307_ (
    .A(_575_),
    .B(_576_),
    .C(_577_),
    .Y(_578_)
);

NAND3X1 _22308_ (
    .A(_543_),
    .B(_574_),
    .C(_578_),
    .Y(_579_)
);

INVX2 _22309_ (
    .A(_543_),
    .Y(_580_)
);

NAND3X1 _22310_ (
    .A(_567_),
    .B(_572_),
    .C(_577_),
    .Y(_581_)
);

OAI21X1 _22311_ (
    .A(_575_),
    .B(_576_),
    .C(_573_),
    .Y(_583_)
);

NAND3X1 _22312_ (
    .A(_580_),
    .B(_581_),
    .C(_583_),
    .Y(_584_)
);

NAND3X1 _22313_ (
    .A(_542_),
    .B(_579_),
    .C(_584_),
    .Y(_585_)
);

NAND2X1 _22314_ (
    .A(_320_),
    .B(_324_),
    .Y(_586_)
);

NOR2X1 _22315_ (
    .A(_333_),
    .B(_586_),
    .Y(_587_)
);

AOI21X1 _22316_ (
    .A(_296_),
    .B(_334_),
    .C(_587_),
    .Y(_588_)
);

AOI21X1 _22317_ (
    .A(_583_),
    .B(_581_),
    .C(_580_),
    .Y(_589_)
);

AOI21X1 _22318_ (
    .A(_574_),
    .B(_578_),
    .C(_543_),
    .Y(_590_)
);

OAI21X1 _22319_ (
    .A(_589_),
    .B(_590_),
    .C(_588_),
    .Y(_591_)
);

NAND3X1 _22320_ (
    .A(_585_),
    .B(_591_),
    .C(_540_),
    .Y(_592_)
);

NAND2X1 _22321_ (
    .A(_539_),
    .B(_535_),
    .Y(_594_)
);

OAI21X1 _22322_ (
    .A(_589_),
    .B(_590_),
    .C(_542_),
    .Y(_595_)
);

NAND3X1 _22323_ (
    .A(_579_),
    .B(_584_),
    .C(_588_),
    .Y(_596_)
);

NAND3X1 _22324_ (
    .A(_594_),
    .B(_595_),
    .C(_596_),
    .Y(_597_)
);

NAND3X1 _22325_ (
    .A(_441_),
    .B(_597_),
    .C(_592_),
    .Y(_598_)
);

AOI21X1 _22326_ (
    .A(_595_),
    .B(_596_),
    .C(_594_),
    .Y(_599_)
);

AOI21X1 _22327_ (
    .A(_585_),
    .B(_591_),
    .C(_540_),
    .Y(_600_)
);

OAI21X1 _22328_ (
    .A(_599_),
    .B(_600_),
    .C(_433_),
    .Y(_601_)
);

NAND3X1 _22329_ (
    .A(_501_),
    .B(_598_),
    .C(_601_),
    .Y(_602_)
);

NAND2X1 _22330_ (
    .A(_340_),
    .B(_348_),
    .Y(_603_)
);

NAND3X1 _22331_ (
    .A(_433_),
    .B(_597_),
    .C(_592_),
    .Y(_605_)
);

OAI21X1 _22332_ (
    .A(_599_),
    .B(_600_),
    .C(_441_),
    .Y(_606_)
);

NAND3X1 _22333_ (
    .A(_603_),
    .B(_605_),
    .C(_606_),
    .Y(_607_)
);

OAI21X1 _22334_ (
    .A(_428_),
    .B(_430_),
    .C(_426_),
    .Y(_608_)
);

NAND2X1 _22335_ (
    .A(areg_23_bF$buf2),
    .B(breg_23_bF$buf1),
    .Y(_609_)
);

NAND2X1 _22336_ (
    .A(breg_22_bF$buf0),
    .B(areg_24_bF$buf0),
    .Y(_610_)
);

NAND2X1 _22337_ (
    .A(breg_21_bF$buf0),
    .B(areg_25_bF$buf4),
    .Y(_611_)
);

OR2X2 _22338_ (
    .A(_610_),
    .B(_611_),
    .Y(_612_)
);

OAI21X1 _22339_ (
    .A(_4069_),
    .B(_5921__bF$buf2),
    .C(_611_),
    .Y(_613_)
);

NAND2X1 _22340_ (
    .A(_613_),
    .B(_612_),
    .Y(_614_)
);

XNOR2X1 _22341_ (
    .A(_614_),
    .B(_609_),
    .Y(_616_)
);

NOR2X1 _22342_ (
    .A(_379_),
    .B(_383_),
    .Y(_617_)
);

AOI21X1 _22343_ (
    .A(_376_),
    .B(_380_),
    .C(_617_),
    .Y(_618_)
);

INVX2 _22344_ (
    .A(_618_),
    .Y(_619_)
);

NOR2X1 _22345_ (
    .A(_3526_),
    .B(_6686__bF$buf2),
    .Y(_620_)
);

INVX1 _22346_ (
    .A(_620_),
    .Y(_621_)
);

NAND2X1 _22347_ (
    .A(breg_19_bF$buf2),
    .B(areg_28_bF$buf4),
    .Y(_622_)
);

OAI21X1 _22348_ (
    .A(_3529__bF$buf2),
    .B(_7520__bF$buf1),
    .C(_378_),
    .Y(_623_)
);

OAI21X1 _22349_ (
    .A(_383_),
    .B(_622_),
    .C(_623_),
    .Y(_624_)
);

NOR2X1 _22350_ (
    .A(_621_),
    .B(_624_),
    .Y(_625_)
);

NAND2X1 _22351_ (
    .A(breg_18_bF$buf3),
    .B(areg_28_bF$buf3),
    .Y(_627_)
);

XOR2X1 _22352_ (
    .A(_378_),
    .B(_627_),
    .Y(_628_)
);

NOR2X1 _22353_ (
    .A(_620_),
    .B(_628_),
    .Y(_629_)
);

OAI21X1 _22354_ (
    .A(_629_),
    .B(_625_),
    .C(_619_),
    .Y(_630_)
);

NAND2X1 _22355_ (
    .A(_620_),
    .B(_628_),
    .Y(_631_)
);

OAI21X1 _22356_ (
    .A(_3526_),
    .B(_6686__bF$buf1),
    .C(_624_),
    .Y(_632_)
);

NAND3X1 _22357_ (
    .A(_618_),
    .B(_632_),
    .C(_631_),
    .Y(_633_)
);

AOI21X1 _22358_ (
    .A(_633_),
    .B(_630_),
    .C(_616_),
    .Y(_634_)
);

INVX2 _22359_ (
    .A(_609_),
    .Y(_635_)
);

XNOR2X1 _22360_ (
    .A(_614_),
    .B(_635_),
    .Y(_636_)
);

NAND3X1 _22361_ (
    .A(_632_),
    .B(_619_),
    .C(_631_),
    .Y(_638_)
);

OAI21X1 _22362_ (
    .A(_629_),
    .B(_625_),
    .C(_618_),
    .Y(_639_)
);

AOI21X1 _22363_ (
    .A(_638_),
    .B(_639_),
    .C(_636_),
    .Y(_640_)
);

NOR2X1 _22364_ (
    .A(_640_),
    .B(_634_),
    .Y(_641_)
);

OR2X2 _22365_ (
    .A(_410_),
    .B(_406_),
    .Y(_642_)
);

NAND2X1 _22366_ (
    .A(breg_17_bF$buf0),
    .B(areg_29_bF$buf1),
    .Y(_643_)
);

NAND2X1 _22367_ (
    .A(breg_15_bF$buf5),
    .B(areg_31_bF$buf1),
    .Y(_644_)
);

OR2X2 _22368_ (
    .A(_405_),
    .B(_644_),
    .Y(_645_)
);

OAI21X1 _22369_ (
    .A(_2362__bF$buf0),
    .B(_8773_),
    .C(_405_),
    .Y(_646_)
);

NAND2X1 _22370_ (
    .A(_646_),
    .B(_645_),
    .Y(_647_)
);

XOR2X1 _22371_ (
    .A(_647_),
    .B(_643_),
    .Y(_649_)
);

XOR2X1 _22372_ (
    .A(_649_),
    .B(_642_),
    .Y(_650_)
);

OAI21X1 _22373_ (
    .A(_421_),
    .B(_419_),
    .C(_650_),
    .Y(_651_)
);

AOI21X1 _22374_ (
    .A(_402_),
    .B(_415_),
    .C(_419_),
    .Y(_652_)
);

XNOR2X1 _22375_ (
    .A(_649_),
    .B(_642_),
    .Y(_653_)
);

NAND2X1 _22376_ (
    .A(_652_),
    .B(_653_),
    .Y(_654_)
);

NAND3X1 _22377_ (
    .A(_641_),
    .B(_654_),
    .C(_651_),
    .Y(_655_)
);

OR2X2 _22378_ (
    .A(_634_),
    .B(_640_),
    .Y(_656_)
);

NOR2X1 _22379_ (
    .A(_652_),
    .B(_653_),
    .Y(_657_)
);

OAI21X1 _22380_ (
    .A(_420_),
    .B(_417_),
    .C(_412_),
    .Y(_658_)
);

NOR2X1 _22381_ (
    .A(_658_),
    .B(_650_),
    .Y(_660_)
);

OAI21X1 _22382_ (
    .A(_660_),
    .B(_657_),
    .C(_656_),
    .Y(_661_)
);

NAND3X1 _22383_ (
    .A(_655_),
    .B(_661_),
    .C(_608_),
    .Y(_662_)
);

AOI21X1 _22384_ (
    .A(_399_),
    .B(_422_),
    .C(_431_),
    .Y(_663_)
);

NOR3X1 _22385_ (
    .A(_657_),
    .B(_656_),
    .C(_660_),
    .Y(_664_)
);

AOI21X1 _22386_ (
    .A(_654_),
    .B(_651_),
    .C(_641_),
    .Y(_665_)
);

OAI21X1 _22387_ (
    .A(_664_),
    .B(_665_),
    .C(_663_),
    .Y(_666_)
);

NAND2X1 _22388_ (
    .A(_662_),
    .B(_666_),
    .Y(_667_)
);

XNOR2X1 _22389_ (
    .A(_439_),
    .B(_667_),
    .Y(_668_)
);

AOI21X1 _22390_ (
    .A(_602_),
    .B(_607_),
    .C(_668_),
    .Y(_669_)
);

NAND3X1 _22391_ (
    .A(_603_),
    .B(_598_),
    .C(_601_),
    .Y(_670_)
);

NAND3X1 _22392_ (
    .A(_501_),
    .B(_605_),
    .C(_606_),
    .Y(_671_)
);

XOR2X1 _22393_ (
    .A(_439_),
    .B(_667_),
    .Y(_672_)
);

AOI21X1 _22394_ (
    .A(_670_),
    .B(_671_),
    .C(_672_),
    .Y(_673_)
);

OAI21X1 _22395_ (
    .A(_669_),
    .B(_673_),
    .C(_500_),
    .Y(_674_)
);

INVX1 _22396_ (
    .A(_448_),
    .Y(_675_)
);

AOI21X1 _22397_ (
    .A(_456_),
    .B(_455_),
    .C(_675_),
    .Y(_676_)
);

NOR2X1 _22398_ (
    .A(_669_),
    .B(_673_),
    .Y(_677_)
);

NAND2X1 _22399_ (
    .A(_677_),
    .B(_676_),
    .Y(_678_)
);

AOI21X1 _22400_ (
    .A(_674_),
    .B(_678_),
    .C(_499_),
    .Y(_679_)
);

OAI21X1 _22401_ (
    .A(_446_),
    .B(_675_),
    .C(_677_),
    .Y(_681_)
);

OAI21X1 _22402_ (
    .A(_669_),
    .B(_673_),
    .C(_676_),
    .Y(_682_)
);

AOI21X1 _22403_ (
    .A(_681_),
    .B(_682_),
    .C(_498_),
    .Y(_683_)
);

OAI21X1 _22404_ (
    .A(_683_),
    .B(_679_),
    .C(_497_),
    .Y(_684_)
);

NOR3X1 _22405_ (
    .A(_452_),
    .B(_449_),
    .C(_446_),
    .Y(_685_)
);

AOI21X1 _22406_ (
    .A(_247_),
    .B(_463_),
    .C(_685_),
    .Y(_686_)
);

NAND3X1 _22407_ (
    .A(_498_),
    .B(_681_),
    .C(_682_),
    .Y(_687_)
);

NAND3X1 _22408_ (
    .A(_670_),
    .B(_671_),
    .C(_672_),
    .Y(_688_)
);

NAND3X1 _22409_ (
    .A(_602_),
    .B(_607_),
    .C(_668_),
    .Y(_689_)
);

NAND2X1 _22410_ (
    .A(_689_),
    .B(_688_),
    .Y(_690_)
);

NOR2X1 _22411_ (
    .A(_690_),
    .B(_676_),
    .Y(_693_)
);

NOR2X1 _22412_ (
    .A(_500_),
    .B(_677_),
    .Y(_694_)
);

OAI21X1 _22413_ (
    .A(_693_),
    .B(_694_),
    .C(_499_),
    .Y(_695_)
);

NAND3X1 _22414_ (
    .A(_687_),
    .B(_686_),
    .C(_695_),
    .Y(_696_)
);

AOI21X1 _22415_ (
    .A(_684_),
    .B(_696_),
    .C(_495_),
    .Y(_697_)
);

NAND3X1 _22416_ (
    .A(_497_),
    .B(_687_),
    .C(_695_),
    .Y(_698_)
);

OAI21X1 _22417_ (
    .A(_683_),
    .B(_679_),
    .C(_686_),
    .Y(_699_)
);

AOI21X1 _22418_ (
    .A(_699_),
    .B(_698_),
    .C(_493_),
    .Y(_700_)
);

OAI21X1 _22419_ (
    .A(_697_),
    .B(_700_),
    .C(_492_),
    .Y(_701_)
);

NOR3X1 _22420_ (
    .A(_460_),
    .B(_464_),
    .C(_468_),
    .Y(_702_)
);

AOI21X1 _22421_ (
    .A(_243_),
    .B(_475_),
    .C(_702_),
    .Y(_704_)
);

NAND3X1 _22422_ (
    .A(_493_),
    .B(_699_),
    .C(_698_),
    .Y(_705_)
);

NAND3X1 _22423_ (
    .A(_495_),
    .B(_684_),
    .C(_696_),
    .Y(_706_)
);

NAND3X1 _22424_ (
    .A(_705_),
    .B(_706_),
    .C(_704_),
    .Y(_707_)
);

AOI22X1 _22425_ (
    .A(_701_),
    .B(_707_),
    .C(_490_),
    .D(_488_),
    .Y(_708_)
);

INVX1 _22426_ (
    .A(_489_),
    .Y(_709_)
);

OAI21X1 _22427_ (
    .A(_11879_),
    .B(_709_),
    .C(_488_),
    .Y(_710_)
);

NAND2X1 _22428_ (
    .A(_701_),
    .B(_707_),
    .Y(_711_)
);

NOR2X1 _22429_ (
    .A(_711_),
    .B(_710_),
    .Y(_712_)
);

NOR2X1 _22430_ (
    .A(_708_),
    .B(_712_),
    .Y(_0_[46])
);

NOR2X1 _22431_ (
    .A(_700_),
    .B(_697_),
    .Y(_714_)
);

OAI21X1 _22432_ (
    .A(_702_),
    .B(_472_),
    .C(_714_),
    .Y(_715_)
);

INVX1 _22433_ (
    .A(_486_),
    .Y(_716_)
);

INVX1 _22434_ (
    .A(_487_),
    .Y(_717_)
);

OAI21X1 _22435_ (
    .A(_237_),
    .B(_717_),
    .C(_716_),
    .Y(_718_)
);

AOI22X1 _22436_ (
    .A(_11869_),
    .B(_11871_),
    .C(_11312_),
    .D(_11874_),
    .Y(_719_)
);

NAND2X1 _22437_ (
    .A(_11877_),
    .B(_10688_),
    .Y(_720_)
);

AOI21X1 _22438_ (
    .A(_719_),
    .B(_720_),
    .C(_709_),
    .Y(_721_)
);

OAI21X1 _22439_ (
    .A(_721_),
    .B(_718_),
    .C(_711_),
    .Y(_722_)
);

AOI21X1 _22440_ (
    .A(_687_),
    .B(_695_),
    .C(_497_),
    .Y(_723_)
);

OAI21X1 _22441_ (
    .A(_723_),
    .B(_495_),
    .C(_698_),
    .Y(_725_)
);

OAI21X1 _22442_ (
    .A(_530_),
    .B(_503_),
    .C(_537_),
    .Y(_726_)
);

INVX1 _22443_ (
    .A(_726_),
    .Y(_727_)
);

OAI21X1 _22444_ (
    .A(_694_),
    .B(_499_),
    .C(_681_),
    .Y(_728_)
);

NAND2X1 _22445_ (
    .A(_598_),
    .B(_670_),
    .Y(_729_)
);

INVX1 _22446_ (
    .A(_729_),
    .Y(_730_)
);

NOR2X1 _22447_ (
    .A(_667_),
    .B(_439_),
    .Y(_731_)
);

AND2X2 _22448_ (
    .A(_592_),
    .B(_585_),
    .Y(_732_)
);

NOR2X1 _22449_ (
    .A(_2669__bF$buf3),
    .B(_7225__bF$buf3),
    .Y(_733_)
);

INVX1 _22450_ (
    .A(_733_),
    .Y(_734_)
);

OAI21X1 _22451_ (
    .A(_520_),
    .B(_507_),
    .C(_528_),
    .Y(_736_)
);

INVX1 _22452_ (
    .A(_736_),
    .Y(_737_)
);

NOR2X1 _22453_ (
    .A(_2884__bF$buf1),
    .B(_6815__bF$buf2),
    .Y(_738_)
);

INVX1 _22454_ (
    .A(_738_),
    .Y(_739_)
);

OAI21X1 _22455_ (
    .A(_513_),
    .B(_509_),
    .C(_517_),
    .Y(_740_)
);

OAI21X1 _22456_ (
    .A(_3958__bF$buf2),
    .B(_5668__bF$buf3),
    .C(_510_),
    .Y(_741_)
);

NAND2X1 _22457_ (
    .A(areg_20_bF$buf1),
    .B(breg_28_bF$buf0),
    .Y(_742_)
);

OAI21X1 _22458_ (
    .A(_512_),
    .B(_742_),
    .C(_741_),
    .Y(_743_)
);

OAI21X1 _22459_ (
    .A(_3146__bF$buf2),
    .B(_6427_),
    .C(_743_),
    .Y(_744_)
);

NOR2X1 _22460_ (
    .A(_3146__bF$buf1),
    .B(_6427_),
    .Y(_745_)
);

NAND2X1 _22461_ (
    .A(areg_20_bF$buf0),
    .B(breg_27_bF$buf0),
    .Y(_747_)
);

XOR2X1 _22462_ (
    .A(_510_),
    .B(_747_),
    .Y(_748_)
);

NAND2X1 _22463_ (
    .A(_745_),
    .B(_748_),
    .Y(_749_)
);

NAND3X1 _22464_ (
    .A(_740_),
    .B(_744_),
    .C(_749_),
    .Y(_750_)
);

INVX1 _22465_ (
    .A(_740_),
    .Y(_751_)
);

NOR2X1 _22466_ (
    .A(_745_),
    .B(_748_),
    .Y(_752_)
);

INVX1 _22467_ (
    .A(_745_),
    .Y(_753_)
);

NOR2X1 _22468_ (
    .A(_753_),
    .B(_743_),
    .Y(_754_)
);

OAI21X1 _22469_ (
    .A(_752_),
    .B(_754_),
    .C(_751_),
    .Y(_755_)
);

NAND3X1 _22470_ (
    .A(_739_),
    .B(_750_),
    .C(_755_),
    .Y(_756_)
);

OAI21X1 _22471_ (
    .A(_752_),
    .B(_754_),
    .C(_740_),
    .Y(_758_)
);

NAND3X1 _22472_ (
    .A(_744_),
    .B(_749_),
    .C(_751_),
    .Y(_759_)
);

NAND3X1 _22473_ (
    .A(_738_),
    .B(_759_),
    .C(_758_),
    .Y(_760_)
);

AOI21X1 _22474_ (
    .A(_756_),
    .B(_760_),
    .C(_737_),
    .Y(_761_)
);

NAND3X1 _22475_ (
    .A(_738_),
    .B(_750_),
    .C(_755_),
    .Y(_762_)
);

NAND3X1 _22476_ (
    .A(_739_),
    .B(_759_),
    .C(_758_),
    .Y(_763_)
);

AOI21X1 _22477_ (
    .A(_762_),
    .B(_763_),
    .C(_736_),
    .Y(_764_)
);

OAI21X1 _22478_ (
    .A(_761_),
    .B(_764_),
    .C(_734_),
    .Y(_765_)
);

NAND3X1 _22479_ (
    .A(_736_),
    .B(_762_),
    .C(_763_),
    .Y(_766_)
);

NAND3X1 _22480_ (
    .A(_756_),
    .B(_760_),
    .C(_737_),
    .Y(_767_)
);

NAND3X1 _22481_ (
    .A(_733_),
    .B(_766_),
    .C(_767_),
    .Y(_769_)
);

AND2X2 _22482_ (
    .A(_765_),
    .B(_769_),
    .Y(_770_)
);

AOI21X1 _22483_ (
    .A(_572_),
    .B(_567_),
    .C(_573_),
    .Y(_771_)
);

OAI21X1 _22484_ (
    .A(_580_),
    .B(_771_),
    .C(_574_),
    .Y(_772_)
);

NAND2X1 _22485_ (
    .A(_559_),
    .B(_567_),
    .Y(_773_)
);

OAI21X1 _22486_ (
    .A(_554_),
    .B(_561_),
    .C(_550_),
    .Y(_774_)
);

NAND2X1 _22487_ (
    .A(areg_21_bF$buf3),
    .B(breg_26_bF$buf4),
    .Y(_775_)
);

AOI22X1 _22488_ (
    .A(areg_22_bF$buf3),
    .B(breg_25_bF$buf4),
    .C(areg_23_bF$buf1),
    .D(breg_24_bF$buf0),
    .Y(_776_)
);

NAND2X1 _22489_ (
    .A(areg_23_bF$buf0),
    .B(breg_25_bF$buf3),
    .Y(_777_)
);

NOR2X1 _22490_ (
    .A(_547_),
    .B(_777_),
    .Y(_778_)
);

OAI21X1 _22491_ (
    .A(_778_),
    .B(_776_),
    .C(_775_),
    .Y(_780_)
);

INVX1 _22492_ (
    .A(_775_),
    .Y(_781_)
);

INVX1 _22493_ (
    .A(_776_),
    .Y(_782_)
);

NAND2X1 _22494_ (
    .A(areg_23_bF$buf4),
    .B(breg_24_bF$buf5),
    .Y(_783_)
);

OR2X2 _22495_ (
    .A(_553_),
    .B(_783_),
    .Y(_784_)
);

NAND3X1 _22496_ (
    .A(_781_),
    .B(_782_),
    .C(_784_),
    .Y(_785_)
);

AND2X2 _22497_ (
    .A(_610_),
    .B(_611_),
    .Y(_786_)
);

OAI21X1 _22498_ (
    .A(_786_),
    .B(_609_),
    .C(_612_),
    .Y(_787_)
);

NAND3X1 _22499_ (
    .A(_780_),
    .B(_787_),
    .C(_785_),
    .Y(_788_)
);

AOI21X1 _22500_ (
    .A(_782_),
    .B(_784_),
    .C(_781_),
    .Y(_789_)
);

NOR3X1 _22501_ (
    .A(_775_),
    .B(_776_),
    .C(_778_),
    .Y(_791_)
);

NOR2X1 _22502_ (
    .A(_610_),
    .B(_611_),
    .Y(_792_)
);

AOI21X1 _22503_ (
    .A(_635_),
    .B(_613_),
    .C(_792_),
    .Y(_793_)
);

OAI21X1 _22504_ (
    .A(_789_),
    .B(_791_),
    .C(_793_),
    .Y(_794_)
);

NAND3X1 _22505_ (
    .A(_774_),
    .B(_788_),
    .C(_794_),
    .Y(_795_)
);

INVX2 _22506_ (
    .A(_774_),
    .Y(_796_)
);

NAND2X1 _22507_ (
    .A(_788_),
    .B(_794_),
    .Y(_797_)
);

NAND2X1 _22508_ (
    .A(_796_),
    .B(_797_),
    .Y(_798_)
);

AOI21X1 _22509_ (
    .A(_632_),
    .B(_631_),
    .C(_619_),
    .Y(_799_)
);

OAI21X1 _22510_ (
    .A(_799_),
    .B(_616_),
    .C(_638_),
    .Y(_800_)
);

NAND3X1 _22511_ (
    .A(_795_),
    .B(_800_),
    .C(_798_),
    .Y(_802_)
);

NAND3X1 _22512_ (
    .A(_793_),
    .B(_780_),
    .C(_785_),
    .Y(_803_)
);

OAI21X1 _22513_ (
    .A(_789_),
    .B(_791_),
    .C(_787_),
    .Y(_804_)
);

AOI21X1 _22514_ (
    .A(_803_),
    .B(_804_),
    .C(_796_),
    .Y(_805_)
);

AOI21X1 _22515_ (
    .A(_788_),
    .B(_794_),
    .C(_774_),
    .Y(_806_)
);

NOR3X1 _22516_ (
    .A(_625_),
    .B(_618_),
    .C(_629_),
    .Y(_807_)
);

AOI21X1 _22517_ (
    .A(_636_),
    .B(_639_),
    .C(_807_),
    .Y(_808_)
);

OAI21X1 _22518_ (
    .A(_805_),
    .B(_806_),
    .C(_808_),
    .Y(_809_)
);

NAND3X1 _22519_ (
    .A(_773_),
    .B(_809_),
    .C(_802_),
    .Y(_810_)
);

AND2X2 _22520_ (
    .A(_567_),
    .B(_559_),
    .Y(_811_)
);

NAND3X1 _22521_ (
    .A(_795_),
    .B(_798_),
    .C(_808_),
    .Y(_813_)
);

OAI21X1 _22522_ (
    .A(_805_),
    .B(_806_),
    .C(_800_),
    .Y(_814_)
);

NAND3X1 _22523_ (
    .A(_811_),
    .B(_814_),
    .C(_813_),
    .Y(_815_)
);

NAND3X1 _22524_ (
    .A(_772_),
    .B(_810_),
    .C(_815_),
    .Y(_816_)
);

NOR3X1 _22525_ (
    .A(_575_),
    .B(_576_),
    .C(_577_),
    .Y(_817_)
);

AOI21X1 _22526_ (
    .A(_543_),
    .B(_578_),
    .C(_817_),
    .Y(_818_)
);

AOI21X1 _22527_ (
    .A(_814_),
    .B(_813_),
    .C(_811_),
    .Y(_819_)
);

AOI21X1 _22528_ (
    .A(_809_),
    .B(_802_),
    .C(_773_),
    .Y(_820_)
);

OAI21X1 _22529_ (
    .A(_819_),
    .B(_820_),
    .C(_818_),
    .Y(_821_)
);

NAND3X1 _22530_ (
    .A(_816_),
    .B(_821_),
    .C(_770_),
    .Y(_822_)
);

NAND2X1 _22531_ (
    .A(_769_),
    .B(_765_),
    .Y(_824_)
);

OAI21X1 _22532_ (
    .A(_819_),
    .B(_820_),
    .C(_772_),
    .Y(_825_)
);

NAND3X1 _22533_ (
    .A(_810_),
    .B(_815_),
    .C(_818_),
    .Y(_826_)
);

NAND3X1 _22534_ (
    .A(_824_),
    .B(_826_),
    .C(_825_),
    .Y(_827_)
);

NAND3X1 _22535_ (
    .A(_662_),
    .B(_827_),
    .C(_822_),
    .Y(_828_)
);

INVX1 _22536_ (
    .A(_662_),
    .Y(_829_)
);

AOI21X1 _22537_ (
    .A(_826_),
    .B(_825_),
    .C(_824_),
    .Y(_830_)
);

AOI21X1 _22538_ (
    .A(_816_),
    .B(_821_),
    .C(_770_),
    .Y(_831_)
);

OAI21X1 _22539_ (
    .A(_830_),
    .B(_831_),
    .C(_829_),
    .Y(_832_)
);

AOI21X1 _22540_ (
    .A(_828_),
    .B(_832_),
    .C(_732_),
    .Y(_833_)
);

NAND2X1 _22541_ (
    .A(_585_),
    .B(_592_),
    .Y(_835_)
);

NAND3X1 _22542_ (
    .A(_829_),
    .B(_827_),
    .C(_822_),
    .Y(_836_)
);

OAI21X1 _22543_ (
    .A(_830_),
    .B(_831_),
    .C(_662_),
    .Y(_837_)
);

AOI21X1 _22544_ (
    .A(_836_),
    .B(_837_),
    .C(_835_),
    .Y(_838_)
);

NOR2X1 _22545_ (
    .A(_657_),
    .B(_664_),
    .Y(_839_)
);

NOR2X1 _22546_ (
    .A(_5369_),
    .B(_5921__bF$buf1),
    .Y(_840_)
);

NAND2X1 _22547_ (
    .A(breg_22_bF$buf4),
    .B(areg_26_bF$buf3),
    .Y(_841_)
);

NOR2X1 _22548_ (
    .A(_611_),
    .B(_841_),
    .Y(_842_)
);

AOI22X1 _22549_ (
    .A(breg_21_bF$buf4),
    .B(areg_26_bF$buf2),
    .C(breg_22_bF$buf3),
    .D(areg_25_bF$buf3),
    .Y(_843_)
);

NOR2X1 _22550_ (
    .A(_843_),
    .B(_842_),
    .Y(_844_)
);

OR2X2 _22551_ (
    .A(_844_),
    .B(_840_),
    .Y(_846_)
);

NAND2X1 _22552_ (
    .A(_840_),
    .B(_844_),
    .Y(_847_)
);

NAND2X1 _22553_ (
    .A(_847_),
    .B(_846_),
    .Y(_848_)
);

NOR2X1 _22554_ (
    .A(_378_),
    .B(_627_),
    .Y(_849_)
);

NOR2X1 _22555_ (
    .A(_849_),
    .B(_625_),
    .Y(_850_)
);

NAND2X1 _22556_ (
    .A(breg_20_bF$buf2),
    .B(areg_27_bF$buf1),
    .Y(_851_)
);

NAND2X1 _22557_ (
    .A(breg_19_bF$buf1),
    .B(areg_29_bF$buf0),
    .Y(_852_)
);

NAND2X1 _22558_ (
    .A(breg_18_bF$buf2),
    .B(areg_29_bF$buf5),
    .Y(_853_)
);

OAI21X1 _22559_ (
    .A(_3253__bF$buf2),
    .B(_7520__bF$buf0),
    .C(_853_),
    .Y(_854_)
);

OAI21X1 _22560_ (
    .A(_627_),
    .B(_852_),
    .C(_854_),
    .Y(_855_)
);

OR2X2 _22561_ (
    .A(_855_),
    .B(_851_),
    .Y(_857_)
);

OAI21X1 _22562_ (
    .A(_3526_),
    .B(_7100__bF$buf1),
    .C(_855_),
    .Y(_858_)
);

NAND2X1 _22563_ (
    .A(_858_),
    .B(_857_),
    .Y(_859_)
);

OR2X2 _22564_ (
    .A(_859_),
    .B(_850_),
    .Y(_860_)
);

NAND2X1 _22565_ (
    .A(_850_),
    .B(_859_),
    .Y(_861_)
);

NAND2X1 _22566_ (
    .A(_861_),
    .B(_860_),
    .Y(_862_)
);

XNOR2X1 _22567_ (
    .A(_862_),
    .B(_848_),
    .Y(_863_)
);

OAI21X1 _22568_ (
    .A(_406_),
    .B(_410_),
    .C(_649_),
    .Y(_864_)
);

OAI21X1 _22569_ (
    .A(_647_),
    .B(_643_),
    .C(_645_),
    .Y(_865_)
);

NAND2X1 _22570_ (
    .A(breg_17_bF$buf4),
    .B(areg_31_bF$buf0),
    .Y(_866_)
);

NOR2X1 _22571_ (
    .A(_405_),
    .B(_866_),
    .Y(_868_)
);

AOI22X1 _22572_ (
    .A(breg_16_bF$buf3),
    .B(areg_31_bF$buf4),
    .C(breg_17_bF$buf3),
    .D(areg_30_bF$buf5),
    .Y(_869_)
);

NOR2X1 _22573_ (
    .A(_869_),
    .B(_868_),
    .Y(_870_)
);

NAND2X1 _22574_ (
    .A(_870_),
    .B(_865_),
    .Y(_871_)
);

INVX1 _22575_ (
    .A(_871_),
    .Y(_872_)
);

NOR2X1 _22576_ (
    .A(_870_),
    .B(_865_),
    .Y(_873_)
);

NOR2X1 _22577_ (
    .A(_873_),
    .B(_872_),
    .Y(_874_)
);

XOR2X1 _22578_ (
    .A(_874_),
    .B(_864_),
    .Y(_875_)
);

XNOR2X1 _22579_ (
    .A(_863_),
    .B(_875_),
    .Y(_876_)
);

NAND2X1 _22580_ (
    .A(_839_),
    .B(_876_),
    .Y(_877_)
);

OR2X2 _22581_ (
    .A(_876_),
    .B(_839_),
    .Y(_879_)
);

NAND2X1 _22582_ (
    .A(_877_),
    .B(_879_),
    .Y(_880_)
);

OAI21X1 _22583_ (
    .A(_833_),
    .B(_838_),
    .C(_880_),
    .Y(_881_)
);

NAND3X1 _22584_ (
    .A(_836_),
    .B(_835_),
    .C(_837_),
    .Y(_882_)
);

NAND3X1 _22585_ (
    .A(_732_),
    .B(_828_),
    .C(_832_),
    .Y(_883_)
);

AND2X2 _22586_ (
    .A(_879_),
    .B(_877_),
    .Y(_884_)
);

NAND3X1 _22587_ (
    .A(_884_),
    .B(_882_),
    .C(_883_),
    .Y(_885_)
);

NAND2X1 _22588_ (
    .A(_885_),
    .B(_881_),
    .Y(_886_)
);

OAI21X1 _22589_ (
    .A(_731_),
    .B(_669_),
    .C(_886_),
    .Y(_887_)
);

NAND2X1 _22590_ (
    .A(_602_),
    .B(_607_),
    .Y(_888_)
);

AOI21X1 _22591_ (
    .A(_672_),
    .B(_888_),
    .C(_731_),
    .Y(_890_)
);

NAND3X1 _22592_ (
    .A(_881_),
    .B(_885_),
    .C(_890_),
    .Y(_891_)
);

AOI21X1 _22593_ (
    .A(_891_),
    .B(_887_),
    .C(_730_),
    .Y(_892_)
);

INVX1 _22594_ (
    .A(_731_),
    .Y(_893_)
);

NAND2X1 _22595_ (
    .A(_893_),
    .B(_688_),
    .Y(_894_)
);

NAND3X1 _22596_ (
    .A(_881_),
    .B(_885_),
    .C(_894_),
    .Y(_895_)
);

NAND2X1 _22597_ (
    .A(_890_),
    .B(_886_),
    .Y(_896_)
);

AOI21X1 _22598_ (
    .A(_895_),
    .B(_896_),
    .C(_729_),
    .Y(_897_)
);

OAI21X1 _22599_ (
    .A(_892_),
    .B(_897_),
    .C(_728_),
    .Y(_898_)
);

AOI21X1 _22600_ (
    .A(_498_),
    .B(_682_),
    .C(_693_),
    .Y(_899_)
);

NAND3X1 _22601_ (
    .A(_729_),
    .B(_895_),
    .C(_896_),
    .Y(_901_)
);

NAND3X1 _22602_ (
    .A(_730_),
    .B(_891_),
    .C(_887_),
    .Y(_902_)
);

NAND3X1 _22603_ (
    .A(_901_),
    .B(_902_),
    .C(_899_),
    .Y(_903_)
);

AOI21X1 _22604_ (
    .A(_903_),
    .B(_898_),
    .C(_727_),
    .Y(_904_)
);

NAND3X1 _22605_ (
    .A(_901_),
    .B(_902_),
    .C(_728_),
    .Y(_905_)
);

OAI21X1 _22606_ (
    .A(_892_),
    .B(_897_),
    .C(_899_),
    .Y(_906_)
);

AOI21X1 _22607_ (
    .A(_905_),
    .B(_906_),
    .C(_726_),
    .Y(_907_)
);

OAI21X1 _22608_ (
    .A(_907_),
    .B(_904_),
    .C(_725_),
    .Y(_908_)
);

NOR3X1 _22609_ (
    .A(_683_),
    .B(_679_),
    .C(_686_),
    .Y(_909_)
);

AOI21X1 _22610_ (
    .A(_493_),
    .B(_699_),
    .C(_909_),
    .Y(_910_)
);

NAND3X1 _22611_ (
    .A(_726_),
    .B(_905_),
    .C(_906_),
    .Y(_912_)
);

NAND3X1 _22612_ (
    .A(_727_),
    .B(_903_),
    .C(_898_),
    .Y(_913_)
);

NAND3X1 _22613_ (
    .A(_912_),
    .B(_913_),
    .C(_910_),
    .Y(_914_)
);

NAND2X1 _22614_ (
    .A(_908_),
    .B(_914_),
    .Y(_915_)
);

NAND3X1 _22615_ (
    .A(_715_),
    .B(_915_),
    .C(_722_),
    .Y(_916_)
);

AND2X2 _22616_ (
    .A(_714_),
    .B(_492_),
    .Y(_917_)
);

INVX1 _22617_ (
    .A(_915_),
    .Y(_918_)
);

OAI21X1 _22618_ (
    .A(_708_),
    .B(_917_),
    .C(_918_),
    .Y(_919_)
);

NAND2X1 _22619_ (
    .A(_916_),
    .B(_919_),
    .Y(_0_[47])
);

AOI22X1 _22620_ (
    .A(_914_),
    .B(_908_),
    .C(_701_),
    .D(_707_),
    .Y(_920_)
);

NAND2X1 _22621_ (
    .A(_920_),
    .B(_489_),
    .Y(_922_)
);

NOR2X1 _22622_ (
    .A(_11875_),
    .B(_922_),
    .Y(_923_)
);

NAND2X1 _22623_ (
    .A(_923_),
    .B(_10686_),
    .Y(_924_)
);

NOR2X1 _22624_ (
    .A(_9974_),
    .B(_9971_),
    .Y(_925_)
);

OAI21X1 _22625_ (
    .A(_9976_),
    .B(_9618_),
    .C(_925_),
    .Y(_926_)
);

INVX1 _22626_ (
    .A(_9985_),
    .Y(_927_)
);

AOI21X1 _22627_ (
    .A(_9633_),
    .B(_926_),
    .C(_927_),
    .Y(_928_)
);

OAI21X1 _22628_ (
    .A(_10649_),
    .B(_10653_),
    .C(_10656_),
    .Y(_929_)
);

INVX1 _22629_ (
    .A(_10680_),
    .Y(_930_)
);

OAI21X1 _22630_ (
    .A(_9992_),
    .B(_10336_),
    .C(_930_),
    .Y(_931_)
);

AOI22X1 _22631_ (
    .A(_931_),
    .B(_929_),
    .C(_928_),
    .D(_10673_),
    .Y(_933_)
);

OAI21X1 _22632_ (
    .A(_9263_),
    .B(_10685_),
    .C(_933_),
    .Y(_934_)
);

OAI21X1 _22633_ (
    .A(_907_),
    .B(_904_),
    .C(_910_),
    .Y(_935_)
);

NOR2X1 _22634_ (
    .A(_904_),
    .B(_907_),
    .Y(_936_)
);

OAI21X1 _22635_ (
    .A(_909_),
    .B(_697_),
    .C(_936_),
    .Y(_937_)
);

NAND2X1 _22636_ (
    .A(_937_),
    .B(_715_),
    .Y(_938_)
);

AOI22X1 _22637_ (
    .A(_935_),
    .B(_938_),
    .C(_718_),
    .D(_920_),
    .Y(_939_)
);

OAI21X1 _22638_ (
    .A(_719_),
    .B(_922_),
    .C(_939_),
    .Y(_940_)
);

AOI21X1 _22639_ (
    .A(_923_),
    .B(_934_),
    .C(_940_),
    .Y(_941_)
);

OAI21X1 _22640_ (
    .A(_7651_),
    .B(_924_),
    .C(_941_),
    .Y(_942_)
);

NAND2X1 _22641_ (
    .A(_905_),
    .B(_912_),
    .Y(_944_)
);

INVX1 _22642_ (
    .A(_944_),
    .Y(_945_)
);

OAI21X1 _22643_ (
    .A(_764_),
    .B(_734_),
    .C(_766_),
    .Y(_946_)
);

OAI21X1 _22644_ (
    .A(_890_),
    .B(_886_),
    .C(_901_),
    .Y(_947_)
);

INVX1 _22645_ (
    .A(_947_),
    .Y(_948_)
);

NAND2X1 _22646_ (
    .A(_836_),
    .B(_882_),
    .Y(_949_)
);

NAND2X1 _22647_ (
    .A(_816_),
    .B(_822_),
    .Y(_950_)
);

INVX1 _22648_ (
    .A(_879_),
    .Y(_951_)
);

NOR2X1 _22649_ (
    .A(_2884__bF$buf0),
    .B(_7225__bF$buf2),
    .Y(_952_)
);

INVX1 _22650_ (
    .A(_952_),
    .Y(_953_)
);

NAND2X1 _22651_ (
    .A(_750_),
    .B(_762_),
    .Y(_955_)
);

INVX1 _22652_ (
    .A(_955_),
    .Y(_956_)
);

NOR2X1 _22653_ (
    .A(_3146__bF$buf0),
    .B(_6815__bF$buf1),
    .Y(_957_)
);

OAI21X1 _22654_ (
    .A(_510_),
    .B(_747_),
    .C(_749_),
    .Y(_958_)
);

NAND2X1 _22655_ (
    .A(areg_21_bF$buf2),
    .B(breg_28_bF$buf5),
    .Y(_959_)
);

OAI21X1 _22656_ (
    .A(_3961__bF$buf3),
    .B(_5668__bF$buf2),
    .C(_742_),
    .Y(_960_)
);

OAI21X1 _22657_ (
    .A(_747_),
    .B(_959_),
    .C(_960_),
    .Y(_961_)
);

OAI21X1 _22658_ (
    .A(_3402__bF$buf1),
    .B(_6427_),
    .C(_961_),
    .Y(_962_)
);

NOR2X1 _22659_ (
    .A(_3402__bF$buf0),
    .B(_6427_),
    .Y(_963_)
);

NAND2X1 _22660_ (
    .A(areg_21_bF$buf1),
    .B(breg_27_bF$buf5),
    .Y(_964_)
);

OR2X2 _22661_ (
    .A(_742_),
    .B(_964_),
    .Y(_966_)
);

NAND3X1 _22662_ (
    .A(_963_),
    .B(_960_),
    .C(_966_),
    .Y(_967_)
);

NAND2X1 _22663_ (
    .A(_967_),
    .B(_962_),
    .Y(_968_)
);

XNOR2X1 _22664_ (
    .A(_958_),
    .B(_968_),
    .Y(_969_)
);

XNOR2X1 _22665_ (
    .A(_969_),
    .B(_957_),
    .Y(_970_)
);

NOR2X1 _22666_ (
    .A(_956_),
    .B(_970_),
    .Y(_971_)
);

XOR2X1 _22667_ (
    .A(_969_),
    .B(_957_),
    .Y(_972_)
);

NOR2X1 _22668_ (
    .A(_955_),
    .B(_972_),
    .Y(_973_)
);

OAI21X1 _22669_ (
    .A(_973_),
    .B(_971_),
    .C(_953_),
    .Y(_974_)
);

NAND2X1 _22670_ (
    .A(_955_),
    .B(_972_),
    .Y(_975_)
);

NAND2X1 _22671_ (
    .A(_956_),
    .B(_970_),
    .Y(_977_)
);

NAND3X1 _22672_ (
    .A(_952_),
    .B(_977_),
    .C(_975_),
    .Y(_978_)
);

AND2X2 _22673_ (
    .A(_974_),
    .B(_978_),
    .Y(_979_)
);

NAND2X1 _22674_ (
    .A(_802_),
    .B(_810_),
    .Y(_980_)
);

OAI21X1 _22675_ (
    .A(_797_),
    .B(_796_),
    .C(_788_),
    .Y(_981_)
);

OAI21X1 _22676_ (
    .A(_775_),
    .B(_776_),
    .C(_784_),
    .Y(_982_)
);

OAI21X1 _22677_ (
    .A(_5921__bF$buf0),
    .B(_5315__bF$buf3),
    .C(_777_),
    .Y(_983_)
);

NAND2X1 _22678_ (
    .A(areg_24_bF$buf4),
    .B(breg_25_bF$buf2),
    .Y(_984_)
);

OAI21X1 _22679_ (
    .A(_783_),
    .B(_984_),
    .C(_983_),
    .Y(_985_)
);

OAI21X1 _22680_ (
    .A(_4551__bF$buf4),
    .B(_5676_),
    .C(_985_),
    .Y(_986_)
);

NOR2X1 _22681_ (
    .A(_4551__bF$buf3),
    .B(_5676_),
    .Y(_988_)
);

NAND2X1 _22682_ (
    .A(areg_24_bF$buf3),
    .B(breg_24_bF$buf4),
    .Y(_989_)
);

OR2X2 _22683_ (
    .A(_777_),
    .B(_989_),
    .Y(_990_)
);

NAND3X1 _22684_ (
    .A(_988_),
    .B(_983_),
    .C(_990_),
    .Y(_991_)
);

NAND2X1 _22685_ (
    .A(_991_),
    .B(_986_),
    .Y(_992_)
);

OAI21X1 _22686_ (
    .A(_611_),
    .B(_841_),
    .C(_847_),
    .Y(_993_)
);

XNOR2X1 _22687_ (
    .A(_993_),
    .B(_992_),
    .Y(_994_)
);

XOR2X1 _22688_ (
    .A(_994_),
    .B(_982_),
    .Y(_995_)
);

OAI21X1 _22689_ (
    .A(_862_),
    .B(_848_),
    .C(_860_),
    .Y(_996_)
);

NAND2X1 _22690_ (
    .A(_996_),
    .B(_995_),
    .Y(_997_)
);

XNOR2X1 _22691_ (
    .A(_994_),
    .B(_982_),
    .Y(_999_)
);

INVX1 _22692_ (
    .A(_848_),
    .Y(_1000_)
);

INVX1 _22693_ (
    .A(_860_),
    .Y(_1001_)
);

AOI21X1 _22694_ (
    .A(_1000_),
    .B(_861_),
    .C(_1001_),
    .Y(_1002_)
);

NAND2X1 _22695_ (
    .A(_1002_),
    .B(_999_),
    .Y(_1003_)
);

NAND3X1 _22696_ (
    .A(_981_),
    .B(_1003_),
    .C(_997_),
    .Y(_1004_)
);

INVX2 _22697_ (
    .A(_981_),
    .Y(_1005_)
);

NOR2X1 _22698_ (
    .A(_1002_),
    .B(_999_),
    .Y(_1006_)
);

NOR2X1 _22699_ (
    .A(_996_),
    .B(_995_),
    .Y(_1007_)
);

OAI21X1 _22700_ (
    .A(_1007_),
    .B(_1006_),
    .C(_1005_),
    .Y(_1008_)
);

NAND3X1 _22701_ (
    .A(_980_),
    .B(_1004_),
    .C(_1008_),
    .Y(_1010_)
);

INVX1 _22702_ (
    .A(_980_),
    .Y(_1011_)
);

NAND2X1 _22703_ (
    .A(_1002_),
    .B(_995_),
    .Y(_1012_)
);

NAND2X1 _22704_ (
    .A(_996_),
    .B(_999_),
    .Y(_1013_)
);

AOI21X1 _22705_ (
    .A(_1013_),
    .B(_1012_),
    .C(_1005_),
    .Y(_1014_)
);

AOI21X1 _22706_ (
    .A(_1003_),
    .B(_997_),
    .C(_981_),
    .Y(_1015_)
);

OAI21X1 _22707_ (
    .A(_1014_),
    .B(_1015_),
    .C(_1011_),
    .Y(_1016_)
);

NAND3X1 _22708_ (
    .A(_1016_),
    .B(_1010_),
    .C(_979_),
    .Y(_1017_)
);

NAND2X1 _22709_ (
    .A(_978_),
    .B(_974_),
    .Y(_1018_)
);

OAI21X1 _22710_ (
    .A(_1014_),
    .B(_1015_),
    .C(_980_),
    .Y(_1019_)
);

NAND3X1 _22711_ (
    .A(_1011_),
    .B(_1004_),
    .C(_1008_),
    .Y(_1021_)
);

NAND3X1 _22712_ (
    .A(_1018_),
    .B(_1019_),
    .C(_1021_),
    .Y(_1022_)
);

NAND3X1 _22713_ (
    .A(_951_),
    .B(_1022_),
    .C(_1017_),
    .Y(_1023_)
);

AOI21X1 _22714_ (
    .A(_1019_),
    .B(_1021_),
    .C(_1018_),
    .Y(_1024_)
);

AOI21X1 _22715_ (
    .A(_1016_),
    .B(_1010_),
    .C(_979_),
    .Y(_1025_)
);

OAI21X1 _22716_ (
    .A(_1024_),
    .B(_1025_),
    .C(_879_),
    .Y(_1026_)
);

NAND3X1 _22717_ (
    .A(_950_),
    .B(_1023_),
    .C(_1026_),
    .Y(_1027_)
);

INVX1 _22718_ (
    .A(_950_),
    .Y(_1028_)
);

NAND3X1 _22719_ (
    .A(_879_),
    .B(_1022_),
    .C(_1017_),
    .Y(_1029_)
);

OAI21X1 _22720_ (
    .A(_1024_),
    .B(_1025_),
    .C(_951_),
    .Y(_1030_)
);

NAND3X1 _22721_ (
    .A(_1028_),
    .B(_1029_),
    .C(_1030_),
    .Y(_1032_)
);

INVX1 _22722_ (
    .A(_874_),
    .Y(_1033_)
);

NOR2X1 _22723_ (
    .A(_864_),
    .B(_1033_),
    .Y(_1034_)
);

NOR2X1 _22724_ (
    .A(_875_),
    .B(_863_),
    .Y(_1035_)
);

NOR2X1 _22725_ (
    .A(_1034_),
    .B(_1035_),
    .Y(_1036_)
);

NOR2X1 _22726_ (
    .A(_5369_),
    .B(_6300__bF$buf0),
    .Y(_1037_)
);

NAND2X1 _22727_ (
    .A(breg_21_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_1038_)
);

XOR2X1 _22728_ (
    .A(_841_),
    .B(_1038_),
    .Y(_1039_)
);

XOR2X1 _22729_ (
    .A(_1039_),
    .B(_1037_),
    .Y(_1040_)
);

OR2X2 _22730_ (
    .A(_622_),
    .B(_853_),
    .Y(_1041_)
);

AND2X2 _22731_ (
    .A(_857_),
    .B(_1041_),
    .Y(_1043_)
);

NAND2X1 _22732_ (
    .A(breg_20_bF$buf1),
    .B(areg_28_bF$buf2),
    .Y(_1044_)
);

NAND2X1 _22733_ (
    .A(breg_19_bF$buf0),
    .B(areg_30_bF$buf4),
    .Y(_1045_)
);

OAI21X1 _22734_ (
    .A(_3529__bF$buf1),
    .B(_8759_),
    .C(_852_),
    .Y(_1046_)
);

OAI21X1 _22735_ (
    .A(_853_),
    .B(_1045_),
    .C(_1046_),
    .Y(_1047_)
);

XNOR2X1 _22736_ (
    .A(_1047_),
    .B(_1044_),
    .Y(_1048_)
);

OR2X2 _22737_ (
    .A(_1043_),
    .B(_1048_),
    .Y(_1049_)
);

NAND2X1 _22738_ (
    .A(_1048_),
    .B(_1043_),
    .Y(_1050_)
);

NAND2X1 _22739_ (
    .A(_1050_),
    .B(_1049_),
    .Y(_1051_)
);

XNOR2X1 _22740_ (
    .A(_1051_),
    .B(_1040_),
    .Y(_1052_)
);

OAI21X1 _22741_ (
    .A(_866_),
    .B(_868_),
    .C(_871_),
    .Y(_1054_)
);

NOR2X1 _22742_ (
    .A(_866_),
    .B(_868_),
    .Y(_1055_)
);

NAND2X1 _22743_ (
    .A(_1055_),
    .B(_872_),
    .Y(_1056_)
);

AND2X2 _22744_ (
    .A(_1056_),
    .B(_1054_),
    .Y(_1057_)
);

XNOR2X1 _22745_ (
    .A(_1052_),
    .B(_1057_),
    .Y(_1058_)
);

NOR2X1 _22746_ (
    .A(_1036_),
    .B(_1058_),
    .Y(_1059_)
);

INVX2 _22747_ (
    .A(_1059_),
    .Y(_1060_)
);

NAND2X1 _22748_ (
    .A(_1036_),
    .B(_1058_),
    .Y(_1061_)
);

NAND2X1 _22749_ (
    .A(_1061_),
    .B(_1060_),
    .Y(_1062_)
);

INVX1 _22750_ (
    .A(_1062_),
    .Y(_1063_)
);

AOI21X1 _22751_ (
    .A(_1027_),
    .B(_1032_),
    .C(_1063_),
    .Y(_1065_)
);

AOI21X1 _22752_ (
    .A(_1029_),
    .B(_1030_),
    .C(_1028_),
    .Y(_1066_)
);

AOI21X1 _22753_ (
    .A(_1023_),
    .B(_1026_),
    .C(_950_),
    .Y(_1067_)
);

NOR3X1 _22754_ (
    .A(_1066_),
    .B(_1062_),
    .C(_1067_),
    .Y(_1068_)
);

OAI21X1 _22755_ (
    .A(_1068_),
    .B(_1065_),
    .C(_885_),
    .Y(_1069_)
);

INVX1 _22756_ (
    .A(_885_),
    .Y(_1070_)
);

OAI21X1 _22757_ (
    .A(_1066_),
    .B(_1067_),
    .C(_1062_),
    .Y(_1071_)
);

NAND3X1 _22758_ (
    .A(_1063_),
    .B(_1027_),
    .C(_1032_),
    .Y(_1072_)
);

NAND3X1 _22759_ (
    .A(_1070_),
    .B(_1072_),
    .C(_1071_),
    .Y(_1073_)
);

AOI21X1 _22760_ (
    .A(_1073_),
    .B(_1069_),
    .C(_949_),
    .Y(_1074_)
);

INVX2 _22761_ (
    .A(_949_),
    .Y(_1076_)
);

AOI21X1 _22762_ (
    .A(_1072_),
    .B(_1071_),
    .C(_1070_),
    .Y(_1077_)
);

NOR3X1 _22763_ (
    .A(_885_),
    .B(_1065_),
    .C(_1068_),
    .Y(_1078_)
);

NOR3X1 _22764_ (
    .A(_1076_),
    .B(_1077_),
    .C(_1078_),
    .Y(_1079_)
);

OAI21X1 _22765_ (
    .A(_1079_),
    .B(_1074_),
    .C(_948_),
    .Y(_1080_)
);

OAI21X1 _22766_ (
    .A(_1078_),
    .B(_1077_),
    .C(_1076_),
    .Y(_1081_)
);

NAND3X1 _22767_ (
    .A(_949_),
    .B(_1073_),
    .C(_1069_),
    .Y(_1082_)
);

NAND3X1 _22768_ (
    .A(_947_),
    .B(_1082_),
    .C(_1081_),
    .Y(_1083_)
);

AOI21X1 _22769_ (
    .A(_1083_),
    .B(_1080_),
    .C(_946_),
    .Y(_1084_)
);

INVX2 _22770_ (
    .A(_946_),
    .Y(_1085_)
);

NAND2X1 _22771_ (
    .A(_1083_),
    .B(_1080_),
    .Y(_1087_)
);

NOR2X1 _22772_ (
    .A(_1085_),
    .B(_1087_),
    .Y(_1088_)
);

OAI21X1 _22773_ (
    .A(_1088_),
    .B(_1084_),
    .C(_945_),
    .Y(_1089_)
);

INVX1 _22774_ (
    .A(_1084_),
    .Y(_1090_)
);

OR2X2 _22775_ (
    .A(_1087_),
    .B(_1085_),
    .Y(_1091_)
);

NAND3X1 _22776_ (
    .A(_944_),
    .B(_1090_),
    .C(_1091_),
    .Y(_1092_)
);

NAND2X1 _22777_ (
    .A(_1089_),
    .B(_1092_),
    .Y(_1093_)
);

XNOR2X1 _22778_ (
    .A(_942_),
    .B(_1093_),
    .Y(_0_[48])
);

NOR3X1 _22779_ (
    .A(_945_),
    .B(_1084_),
    .C(_1088_),
    .Y(_1094_)
);

AOI21X1 _22780_ (
    .A(_1089_),
    .B(_942_),
    .C(_1094_),
    .Y(_1095_)
);

AOI21X1 _22781_ (
    .A(_1082_),
    .B(_1081_),
    .C(_947_),
    .Y(_1097_)
);

OAI21X1 _22782_ (
    .A(_1097_),
    .B(_1085_),
    .C(_1083_),
    .Y(_1098_)
);

OAI21X1 _22783_ (
    .A(_973_),
    .B(_953_),
    .C(_975_),
    .Y(_1099_)
);

INVX2 _22784_ (
    .A(_1099_),
    .Y(_1100_)
);

OAI21X1 _22785_ (
    .A(_1077_),
    .B(_1076_),
    .C(_1073_),
    .Y(_1101_)
);

NAND2X1 _22786_ (
    .A(_1023_),
    .B(_1027_),
    .Y(_1102_)
);

INVX2 _22787_ (
    .A(_1102_),
    .Y(_1103_)
);

NAND2X1 _22788_ (
    .A(_1010_),
    .B(_1017_),
    .Y(_1104_)
);

NOR2X1 _22789_ (
    .A(_3146__bF$buf3),
    .B(_7225__bF$buf1),
    .Y(_1105_)
);

INVX1 _22790_ (
    .A(_1105_),
    .Y(_1106_)
);

NAND3X1 _22791_ (
    .A(_962_),
    .B(_967_),
    .C(_958_),
    .Y(_1108_)
);

NAND2X1 _22792_ (
    .A(_957_),
    .B(_969_),
    .Y(_1109_)
);

NAND2X1 _22793_ (
    .A(_1108_),
    .B(_1109_),
    .Y(_1110_)
);

NOR2X1 _22794_ (
    .A(_3402__bF$buf3),
    .B(_6815__bF$buf0),
    .Y(_1111_)
);

OAI21X1 _22795_ (
    .A(_747_),
    .B(_959_),
    .C(_967_),
    .Y(_1112_)
);

NAND2X1 _22796_ (
    .A(areg_22_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_1113_)
);

OAI21X1 _22797_ (
    .A(_4551__bF$buf2),
    .B(_5668__bF$buf1),
    .C(_959_),
    .Y(_1114_)
);

OAI21X1 _22798_ (
    .A(_964_),
    .B(_1113_),
    .C(_1114_),
    .Y(_1115_)
);

OAI21X1 _22799_ (
    .A(_3958__bF$buf1),
    .B(_6427_),
    .C(_1115_),
    .Y(_1116_)
);

NOR2X1 _22800_ (
    .A(_3958__bF$buf0),
    .B(_6427_),
    .Y(_1117_)
);

NAND2X1 _22801_ (
    .A(areg_22_bF$buf1),
    .B(breg_27_bF$buf4),
    .Y(_1119_)
);

OR2X2 _22802_ (
    .A(_959_),
    .B(_1119_),
    .Y(_1120_)
);

NAND3X1 _22803_ (
    .A(_1117_),
    .B(_1114_),
    .C(_1120_),
    .Y(_1121_)
);

NAND2X1 _22804_ (
    .A(_1121_),
    .B(_1116_),
    .Y(_1122_)
);

XNOR2X1 _22805_ (
    .A(_1122_),
    .B(_1112_),
    .Y(_1123_)
);

XOR2X1 _22806_ (
    .A(_1123_),
    .B(_1111_),
    .Y(_1124_)
);

AND2X2 _22807_ (
    .A(_1110_),
    .B(_1124_),
    .Y(_1125_)
);

NOR2X1 _22808_ (
    .A(_1124_),
    .B(_1110_),
    .Y(_1126_)
);

OAI21X1 _22809_ (
    .A(_1125_),
    .B(_1126_),
    .C(_1106_),
    .Y(_1127_)
);

NAND2X1 _22810_ (
    .A(_1124_),
    .B(_1110_),
    .Y(_1128_)
);

OR2X2 _22811_ (
    .A(_1110_),
    .B(_1124_),
    .Y(_1130_)
);

NAND3X1 _22812_ (
    .A(_1105_),
    .B(_1128_),
    .C(_1130_),
    .Y(_1131_)
);

AND2X2 _22813_ (
    .A(_1131_),
    .B(_1127_),
    .Y(_1132_)
);

OAI21X1 _22814_ (
    .A(_1007_),
    .B(_1005_),
    .C(_997_),
    .Y(_1133_)
);

NAND3X1 _22815_ (
    .A(_986_),
    .B(_991_),
    .C(_993_),
    .Y(_1134_)
);

OAI21X1 _22816_ (
    .A(_778_),
    .B(_791_),
    .C(_994_),
    .Y(_1135_)
);

NAND2X1 _22817_ (
    .A(_1134_),
    .B(_1135_),
    .Y(_1136_)
);

OAI21X1 _22818_ (
    .A(_777_),
    .B(_989_),
    .C(_991_),
    .Y(_1137_)
);

OAI21X1 _22819_ (
    .A(_5315__bF$buf2),
    .B(_6300__bF$buf3),
    .C(_984_),
    .Y(_1138_)
);

NAND2X1 _22820_ (
    .A(areg_25_bF$buf2),
    .B(breg_25_bF$buf1),
    .Y(_1139_)
);

OAI21X1 _22821_ (
    .A(_989_),
    .B(_1139_),
    .C(_1138_),
    .Y(_1141_)
);

OAI21X1 _22822_ (
    .A(_4541__bF$buf0),
    .B(_5676_),
    .C(_1141_),
    .Y(_1142_)
);

NOR2X1 _22823_ (
    .A(_4541__bF$buf4),
    .B(_5676_),
    .Y(_1143_)
);

NAND2X1 _22824_ (
    .A(breg_24_bF$buf3),
    .B(areg_25_bF$buf1),
    .Y(_1144_)
);

OR2X2 _22825_ (
    .A(_984_),
    .B(_1144_),
    .Y(_1145_)
);

NAND3X1 _22826_ (
    .A(_1143_),
    .B(_1138_),
    .C(_1145_),
    .Y(_1146_)
);

NAND2X1 _22827_ (
    .A(_1146_),
    .B(_1142_),
    .Y(_1147_)
);

NAND2X1 _22828_ (
    .A(_1037_),
    .B(_1039_),
    .Y(_1148_)
);

OAI21X1 _22829_ (
    .A(_841_),
    .B(_1038_),
    .C(_1148_),
    .Y(_1149_)
);

XNOR2X1 _22830_ (
    .A(_1149_),
    .B(_1147_),
    .Y(_1150_)
);

XOR2X1 _22831_ (
    .A(_1150_),
    .B(_1137_),
    .Y(_1152_)
);

INVX1 _22832_ (
    .A(_1040_),
    .Y(_1153_)
);

OAI21X1 _22833_ (
    .A(_1051_),
    .B(_1153_),
    .C(_1049_),
    .Y(_1154_)
);

NAND2X1 _22834_ (
    .A(_1152_),
    .B(_1154_),
    .Y(_1155_)
);

XNOR2X1 _22835_ (
    .A(_1150_),
    .B(_1137_),
    .Y(_1156_)
);

INVX1 _22836_ (
    .A(_1049_),
    .Y(_1157_)
);

AOI21X1 _22837_ (
    .A(_1040_),
    .B(_1050_),
    .C(_1157_),
    .Y(_1158_)
);

NAND2X1 _22838_ (
    .A(_1158_),
    .B(_1156_),
    .Y(_1159_)
);

NAND3X1 _22839_ (
    .A(_1136_),
    .B(_1159_),
    .C(_1155_),
    .Y(_1160_)
);

INVX2 _22840_ (
    .A(_1136_),
    .Y(_1161_)
);

NOR2X1 _22841_ (
    .A(_1158_),
    .B(_1156_),
    .Y(_1163_)
);

NOR2X1 _22842_ (
    .A(_1152_),
    .B(_1154_),
    .Y(_1164_)
);

OAI21X1 _22843_ (
    .A(_1164_),
    .B(_1163_),
    .C(_1161_),
    .Y(_1165_)
);

NAND3X1 _22844_ (
    .A(_1160_),
    .B(_1133_),
    .C(_1165_),
    .Y(_1166_)
);

AOI21X1 _22845_ (
    .A(_981_),
    .B(_1003_),
    .C(_1006_),
    .Y(_1167_)
);

NAND2X1 _22846_ (
    .A(_1158_),
    .B(_1152_),
    .Y(_1168_)
);

NAND2X1 _22847_ (
    .A(_1156_),
    .B(_1154_),
    .Y(_1169_)
);

AOI21X1 _22848_ (
    .A(_1168_),
    .B(_1169_),
    .C(_1161_),
    .Y(_1170_)
);

AOI21X1 _22849_ (
    .A(_1159_),
    .B(_1155_),
    .C(_1136_),
    .Y(_1171_)
);

OAI21X1 _22850_ (
    .A(_1170_),
    .B(_1171_),
    .C(_1167_),
    .Y(_1172_)
);

NAND3X1 _22851_ (
    .A(_1166_),
    .B(_1172_),
    .C(_1132_),
    .Y(_1174_)
);

NAND2X1 _22852_ (
    .A(_1127_),
    .B(_1131_),
    .Y(_1175_)
);

OAI21X1 _22853_ (
    .A(_1170_),
    .B(_1171_),
    .C(_1133_),
    .Y(_1176_)
);

NAND3X1 _22854_ (
    .A(_1167_),
    .B(_1160_),
    .C(_1165_),
    .Y(_1177_)
);

NAND3X1 _22855_ (
    .A(_1175_),
    .B(_1176_),
    .C(_1177_),
    .Y(_1178_)
);

NAND3X1 _22856_ (
    .A(_1059_),
    .B(_1178_),
    .C(_1174_),
    .Y(_1179_)
);

AOI21X1 _22857_ (
    .A(_1176_),
    .B(_1177_),
    .C(_1175_),
    .Y(_1180_)
);

AOI21X1 _22858_ (
    .A(_1166_),
    .B(_1172_),
    .C(_1132_),
    .Y(_1181_)
);

OAI21X1 _22859_ (
    .A(_1181_),
    .B(_1180_),
    .C(_1060_),
    .Y(_1182_)
);

NAND3X1 _22860_ (
    .A(_1104_),
    .B(_1179_),
    .C(_1182_),
    .Y(_1183_)
);

AND2X2 _22861_ (
    .A(_1017_),
    .B(_1010_),
    .Y(_1185_)
);

NAND3X1 _22862_ (
    .A(_1060_),
    .B(_1178_),
    .C(_1174_),
    .Y(_1186_)
);

OAI21X1 _22863_ (
    .A(_1181_),
    .B(_1180_),
    .C(_1059_),
    .Y(_1187_)
);

NAND3X1 _22864_ (
    .A(_1185_),
    .B(_1186_),
    .C(_1187_),
    .Y(_1188_)
);

INVX1 _22865_ (
    .A(_1056_),
    .Y(_1189_)
);

AOI21X1 _22866_ (
    .A(_1054_),
    .B(_1052_),
    .C(_1189_),
    .Y(_1190_)
);

NOR2X1 _22867_ (
    .A(_5369_),
    .B(_6686__bF$buf0),
    .Y(_1191_)
);

NAND2X1 _22868_ (
    .A(breg_22_bF$buf2),
    .B(areg_28_bF$buf1),
    .Y(_1192_)
);

NOR2X1 _22869_ (
    .A(_1038_),
    .B(_1192_),
    .Y(_1193_)
);

AOI22X1 _22870_ (
    .A(breg_21_bF$buf2),
    .B(areg_28_bF$buf0),
    .C(breg_22_bF$buf1),
    .D(areg_27_bF$buf5),
    .Y(_1194_)
);

NOR2X1 _22871_ (
    .A(_1194_),
    .B(_1193_),
    .Y(_1196_)
);

OR2X2 _22872_ (
    .A(_1196_),
    .B(_1191_),
    .Y(_1197_)
);

NAND2X1 _22873_ (
    .A(_1191_),
    .B(_1196_),
    .Y(_1198_)
);

AND2X2 _22874_ (
    .A(_1197_),
    .B(_1198_),
    .Y(_1199_)
);

INVX1 _22875_ (
    .A(_1044_),
    .Y(_1200_)
);

NOR2X1 _22876_ (
    .A(_853_),
    .B(_1045_),
    .Y(_1201_)
);

AOI21X1 _22877_ (
    .A(_1200_),
    .B(_1046_),
    .C(_1201_),
    .Y(_1202_)
);

NOR2X1 _22878_ (
    .A(_3526_),
    .B(_9153_),
    .Y(_1203_)
);

NAND2X1 _22879_ (
    .A(breg_18_bF$buf1),
    .B(areg_31_bF$buf3),
    .Y(_1204_)
);

OR2X2 _22880_ (
    .A(_1045_),
    .B(_1204_),
    .Y(_1205_)
);

OAI21X1 _22881_ (
    .A(_3529__bF$buf0),
    .B(_8773_),
    .C(_1045_),
    .Y(_1207_)
);

NAND3X1 _22882_ (
    .A(_1203_),
    .B(_1207_),
    .C(_1205_),
    .Y(_1208_)
);

NAND2X1 _22883_ (
    .A(_1207_),
    .B(_1205_),
    .Y(_1209_)
);

OAI21X1 _22884_ (
    .A(_3526_),
    .B(_9153_),
    .C(_1209_),
    .Y(_1210_)
);

NAND2X1 _22885_ (
    .A(_1208_),
    .B(_1210_),
    .Y(_1211_)
);

XOR2X1 _22886_ (
    .A(_1211_),
    .B(_1202_),
    .Y(_1212_)
);

XOR2X1 _22887_ (
    .A(_1212_),
    .B(_1199_),
    .Y(_1213_)
);

XNOR2X1 _22888_ (
    .A(_1213_),
    .B(_868_),
    .Y(_1214_)
);

NAND2X1 _22889_ (
    .A(_1214_),
    .B(_1190_),
    .Y(_1215_)
);

NOR2X1 _22890_ (
    .A(_1214_),
    .B(_1190_),
    .Y(_1216_)
);

INVX2 _22891_ (
    .A(_1216_),
    .Y(_1218_)
);

NAND2X1 _22892_ (
    .A(_1215_),
    .B(_1218_),
    .Y(_1219_)
);

NAND3X1 _22893_ (
    .A(_1219_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1220_)
);

AOI21X1 _22894_ (
    .A(_1186_),
    .B(_1187_),
    .C(_1185_),
    .Y(_1221_)
);

AOI21X1 _22895_ (
    .A(_1179_),
    .B(_1182_),
    .C(_1104_),
    .Y(_1222_)
);

INVX1 _22896_ (
    .A(_1219_),
    .Y(_1223_)
);

OAI21X1 _22897_ (
    .A(_1221_),
    .B(_1222_),
    .C(_1223_),
    .Y(_1224_)
);

AOI21X1 _22898_ (
    .A(_1220_),
    .B(_1224_),
    .C(_1072_),
    .Y(_1225_)
);

NAND3X1 _22899_ (
    .A(_1223_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1226_)
);

OAI21X1 _22900_ (
    .A(_1221_),
    .B(_1222_),
    .C(_1219_),
    .Y(_1227_)
);

AOI21X1 _22901_ (
    .A(_1226_),
    .B(_1227_),
    .C(_1068_),
    .Y(_1229_)
);

NOR3X1 _22902_ (
    .A(_1225_),
    .B(_1103_),
    .C(_1229_),
    .Y(_1230_)
);

NAND3X1 _22903_ (
    .A(_1226_),
    .B(_1227_),
    .C(_1068_),
    .Y(_1231_)
);

NAND3X1 _22904_ (
    .A(_1072_),
    .B(_1220_),
    .C(_1224_),
    .Y(_1232_)
);

AOI21X1 _22905_ (
    .A(_1232_),
    .B(_1231_),
    .C(_1102_),
    .Y(_1233_)
);

OAI21X1 _22906_ (
    .A(_1230_),
    .B(_1233_),
    .C(_1101_),
    .Y(_1234_)
);

AOI21X1 _22907_ (
    .A(_1069_),
    .B(_949_),
    .C(_1078_),
    .Y(_1235_)
);

NAND3X1 _22908_ (
    .A(_1102_),
    .B(_1232_),
    .C(_1231_),
    .Y(_1236_)
);

OAI21X1 _22909_ (
    .A(_1229_),
    .B(_1225_),
    .C(_1103_),
    .Y(_1237_)
);

NAND3X1 _22910_ (
    .A(_1236_),
    .B(_1237_),
    .C(_1235_),
    .Y(_1238_)
);

AOI21X1 _22911_ (
    .A(_1238_),
    .B(_1234_),
    .C(_1100_),
    .Y(_1240_)
);

NAND3X1 _22912_ (
    .A(_1101_),
    .B(_1236_),
    .C(_1237_),
    .Y(_1241_)
);

OAI21X1 _22913_ (
    .A(_1230_),
    .B(_1233_),
    .C(_1235_),
    .Y(_1242_)
);

AOI21X1 _22914_ (
    .A(_1241_),
    .B(_1242_),
    .C(_1099_),
    .Y(_1243_)
);

OAI21X1 _22915_ (
    .A(_1240_),
    .B(_1243_),
    .C(_1098_),
    .Y(_1244_)
);

NOR3X1 _22916_ (
    .A(_948_),
    .B(_1074_),
    .C(_1079_),
    .Y(_1245_)
);

AOI21X1 _22917_ (
    .A(_946_),
    .B(_1080_),
    .C(_1245_),
    .Y(_1246_)
);

NAND3X1 _22918_ (
    .A(_1099_),
    .B(_1241_),
    .C(_1242_),
    .Y(_1247_)
);

NOR3X1 _22919_ (
    .A(_1235_),
    .B(_1233_),
    .C(_1230_),
    .Y(_1248_)
);

AOI21X1 _22920_ (
    .A(_1236_),
    .B(_1237_),
    .C(_1101_),
    .Y(_1249_)
);

OAI21X1 _22921_ (
    .A(_1248_),
    .B(_1249_),
    .C(_1100_),
    .Y(_1251_)
);

NAND3X1 _22922_ (
    .A(_1247_),
    .B(_1251_),
    .C(_1246_),
    .Y(_1252_)
);

NAND2X1 _22923_ (
    .A(_1244_),
    .B(_1252_),
    .Y(_1253_)
);

XNOR2X1 _22924_ (
    .A(_1095_),
    .B(_1253_),
    .Y(_0_[49])
);

NAND3X1 _22925_ (
    .A(_1098_),
    .B(_1247_),
    .C(_1251_),
    .Y(_1254_)
);

OAI21X1 _22926_ (
    .A(_1240_),
    .B(_1243_),
    .C(_1246_),
    .Y(_1255_)
);

NAND2X1 _22927_ (
    .A(_1255_),
    .B(_1254_),
    .Y(_1256_)
);

OAI21X1 _22928_ (
    .A(_1092_),
    .B(_1256_),
    .C(_1254_),
    .Y(_1257_)
);

NAND3X1 _22929_ (
    .A(_1089_),
    .B(_1253_),
    .C(_1092_),
    .Y(_1258_)
);

INVX1 _22930_ (
    .A(_1258_),
    .Y(_1259_)
);

AOI21X1 _22931_ (
    .A(_1259_),
    .B(_942_),
    .C(_1257_),
    .Y(_1261_)
);

OAI21X1 _22932_ (
    .A(_1249_),
    .B(_1100_),
    .C(_1241_),
    .Y(_1262_)
);

OAI21X1 _22933_ (
    .A(_1126_),
    .B(_1106_),
    .C(_1128_),
    .Y(_1263_)
);

INVX1 _22934_ (
    .A(_1263_),
    .Y(_1264_)
);

OAI21X1 _22935_ (
    .A(_1229_),
    .B(_1103_),
    .C(_1231_),
    .Y(_1265_)
);

NAND2X1 _22936_ (
    .A(_1179_),
    .B(_1183_),
    .Y(_1266_)
);

INVX2 _22937_ (
    .A(_1266_),
    .Y(_1267_)
);

NAND2X1 _22938_ (
    .A(_1166_),
    .B(_1174_),
    .Y(_1268_)
);

NAND3X1 _22939_ (
    .A(_1116_),
    .B(_1121_),
    .C(_1112_),
    .Y(_1269_)
);

NAND2X1 _22940_ (
    .A(_1111_),
    .B(_1123_),
    .Y(_1270_)
);

NAND2X1 _22941_ (
    .A(_1269_),
    .B(_1270_),
    .Y(_1272_)
);

NOR2X1 _22942_ (
    .A(_3958__bF$buf3),
    .B(_6815__bF$buf4),
    .Y(_1273_)
);

AND2X2 _22943_ (
    .A(_1121_),
    .B(_1120_),
    .Y(_1274_)
);

NAND2X1 _22944_ (
    .A(areg_23_bF$buf3),
    .B(breg_28_bF$buf3),
    .Y(_1275_)
);

OAI21X1 _22945_ (
    .A(_4541__bF$buf3),
    .B(_5668__bF$buf0),
    .C(_1113_),
    .Y(_1276_)
);

OAI21X1 _22946_ (
    .A(_1119_),
    .B(_1275_),
    .C(_1276_),
    .Y(_1277_)
);

OAI21X1 _22947_ (
    .A(_3961__bF$buf2),
    .B(_6427_),
    .C(_1277_),
    .Y(_1278_)
);

NAND2X1 _22948_ (
    .A(areg_21_bF$buf0),
    .B(breg_29_bF$buf1),
    .Y(_1279_)
);

OR2X2 _22949_ (
    .A(_1277_),
    .B(_1279_),
    .Y(_1280_)
);

NAND2X1 _22950_ (
    .A(_1278_),
    .B(_1280_),
    .Y(_1281_)
);

XOR2X1 _22951_ (
    .A(_1281_),
    .B(_1274_),
    .Y(_1283_)
);

XOR2X1 _22952_ (
    .A(_1283_),
    .B(_1273_),
    .Y(_1284_)
);

NAND2X1 _22953_ (
    .A(_1272_),
    .B(_1284_),
    .Y(_1285_)
);

AND2X2 _22954_ (
    .A(_1270_),
    .B(_1269_),
    .Y(_1286_)
);

XNOR2X1 _22955_ (
    .A(_1283_),
    .B(_1273_),
    .Y(_1287_)
);

NAND2X1 _22956_ (
    .A(_1286_),
    .B(_1287_),
    .Y(_1288_)
);

NAND2X1 _22957_ (
    .A(_1288_),
    .B(_1285_),
    .Y(_1289_)
);

OAI21X1 _22958_ (
    .A(_3402__bF$buf2),
    .B(_7225__bF$buf0),
    .C(_1289_),
    .Y(_1290_)
);

NOR2X1 _22959_ (
    .A(_3402__bF$buf1),
    .B(_7225__bF$buf4),
    .Y(_1291_)
);

NAND3X1 _22960_ (
    .A(_1291_),
    .B(_1288_),
    .C(_1285_),
    .Y(_1292_)
);

AND2X2 _22961_ (
    .A(_1290_),
    .B(_1292_),
    .Y(_1294_)
);

OAI21X1 _22962_ (
    .A(_1164_),
    .B(_1161_),
    .C(_1155_),
    .Y(_1295_)
);

NAND3X1 _22963_ (
    .A(_1142_),
    .B(_1146_),
    .C(_1149_),
    .Y(_1296_)
);

NAND2X1 _22964_ (
    .A(_1137_),
    .B(_1150_),
    .Y(_1297_)
);

NAND2X1 _22965_ (
    .A(_1296_),
    .B(_1297_),
    .Y(_1298_)
);

OAI21X1 _22966_ (
    .A(_989_),
    .B(_1139_),
    .C(_1146_),
    .Y(_1299_)
);

OAI21X1 _22967_ (
    .A(_5315__bF$buf1),
    .B(_6686__bF$buf3),
    .C(_1139_),
    .Y(_1300_)
);

NAND2X1 _22968_ (
    .A(breg_25_bF$buf0),
    .B(areg_26_bF$buf1),
    .Y(_1301_)
);

OAI21X1 _22969_ (
    .A(_1144_),
    .B(_1301_),
    .C(_1300_),
    .Y(_1302_)
);

OAI21X1 _22970_ (
    .A(_5921__bF$buf3),
    .B(_5676_),
    .C(_1302_),
    .Y(_1303_)
);

NOR2X1 _22971_ (
    .A(_5921__bF$buf2),
    .B(_5676_),
    .Y(_1304_)
);

NAND2X1 _22972_ (
    .A(breg_24_bF$buf2),
    .B(areg_26_bF$buf0),
    .Y(_1305_)
);

OR2X2 _22973_ (
    .A(_1139_),
    .B(_1305_),
    .Y(_1306_)
);

NAND3X1 _22974_ (
    .A(_1304_),
    .B(_1300_),
    .C(_1306_),
    .Y(_1307_)
);

NAND2X1 _22975_ (
    .A(_1307_),
    .B(_1303_),
    .Y(_1308_)
);

OAI21X1 _22976_ (
    .A(_1038_),
    .B(_1192_),
    .C(_1198_),
    .Y(_1309_)
);

XNOR2X1 _22977_ (
    .A(_1309_),
    .B(_1308_),
    .Y(_1310_)
);

XOR2X1 _22978_ (
    .A(_1310_),
    .B(_1299_),
    .Y(_1311_)
);

NOR2X1 _22979_ (
    .A(_1202_),
    .B(_1211_),
    .Y(_1312_)
);

AOI21X1 _22980_ (
    .A(_1199_),
    .B(_1212_),
    .C(_1312_),
    .Y(_1313_)
);

INVX1 _22981_ (
    .A(_1313_),
    .Y(_1315_)
);

NAND2X1 _22982_ (
    .A(_1311_),
    .B(_1315_),
    .Y(_1316_)
);

XNOR2X1 _22983_ (
    .A(_1310_),
    .B(_1299_),
    .Y(_1317_)
);

NAND2X1 _22984_ (
    .A(_1313_),
    .B(_1317_),
    .Y(_1318_)
);

NAND3X1 _22985_ (
    .A(_1298_),
    .B(_1318_),
    .C(_1316_),
    .Y(_1319_)
);

INVX2 _22986_ (
    .A(_1298_),
    .Y(_1320_)
);

NOR2X1 _22987_ (
    .A(_1313_),
    .B(_1317_),
    .Y(_1321_)
);

NOR2X1 _22988_ (
    .A(_1311_),
    .B(_1315_),
    .Y(_1322_)
);

OAI21X1 _22989_ (
    .A(_1322_),
    .B(_1321_),
    .C(_1320_),
    .Y(_1323_)
);

NAND3X1 _22990_ (
    .A(_1319_),
    .B(_1323_),
    .C(_1295_),
    .Y(_1324_)
);

AOI21X1 _22991_ (
    .A(_1136_),
    .B(_1159_),
    .C(_1163_),
    .Y(_1326_)
);

NOR3X1 _22992_ (
    .A(_1321_),
    .B(_1320_),
    .C(_1322_),
    .Y(_1327_)
);

AOI21X1 _22993_ (
    .A(_1318_),
    .B(_1316_),
    .C(_1298_),
    .Y(_1328_)
);

OAI21X1 _22994_ (
    .A(_1327_),
    .B(_1328_),
    .C(_1326_),
    .Y(_1329_)
);

NAND3X1 _22995_ (
    .A(_1324_),
    .B(_1329_),
    .C(_1294_),
    .Y(_1330_)
);

NAND2X1 _22996_ (
    .A(_1292_),
    .B(_1290_),
    .Y(_1331_)
);

OAI21X1 _22997_ (
    .A(_1327_),
    .B(_1328_),
    .C(_1295_),
    .Y(_1332_)
);

NAND3X1 _22998_ (
    .A(_1326_),
    .B(_1319_),
    .C(_1323_),
    .Y(_1333_)
);

NAND3X1 _22999_ (
    .A(_1333_),
    .B(_1331_),
    .C(_1332_),
    .Y(_1334_)
);

NAND3X1 _23000_ (
    .A(_1216_),
    .B(_1334_),
    .C(_1330_),
    .Y(_1335_)
);

AOI21X1 _23001_ (
    .A(_1333_),
    .B(_1332_),
    .C(_1331_),
    .Y(_1337_)
);

AOI21X1 _23002_ (
    .A(_1324_),
    .B(_1329_),
    .C(_1294_),
    .Y(_1338_)
);

OAI21X1 _23003_ (
    .A(_1338_),
    .B(_1337_),
    .C(_1218_),
    .Y(_1339_)
);

NAND3X1 _23004_ (
    .A(_1268_),
    .B(_1335_),
    .C(_1339_),
    .Y(_1340_)
);

INVX1 _23005_ (
    .A(_1268_),
    .Y(_1341_)
);

NAND3X1 _23006_ (
    .A(_1218_),
    .B(_1334_),
    .C(_1330_),
    .Y(_1342_)
);

OAI21X1 _23007_ (
    .A(_1338_),
    .B(_1337_),
    .C(_1216_),
    .Y(_1343_)
);

NAND3X1 _23008_ (
    .A(_1342_),
    .B(_1343_),
    .C(_1341_),
    .Y(_1344_)
);

NAND2X1 _23009_ (
    .A(_868_),
    .B(_1213_),
    .Y(_1345_)
);

NAND2X1 _23010_ (
    .A(breg_23_bF$buf0),
    .B(areg_27_bF$buf4),
    .Y(_1346_)
);

NAND2X1 _23011_ (
    .A(breg_21_bF$buf1),
    .B(areg_29_bF$buf4),
    .Y(_1348_)
);

XOR2X1 _23012_ (
    .A(_1192_),
    .B(_1348_),
    .Y(_1349_)
);

XNOR2X1 _23013_ (
    .A(_1349_),
    .B(_1346_),
    .Y(_1350_)
);

OAI21X1 _23014_ (
    .A(_1045_),
    .B(_1204_),
    .C(_1208_),
    .Y(_1351_)
);

NAND2X1 _23015_ (
    .A(breg_20_bF$buf0),
    .B(areg_31_bF$buf2),
    .Y(_1352_)
);

NOR2X1 _23016_ (
    .A(_1045_),
    .B(_1352_),
    .Y(_1353_)
);

AOI22X1 _23017_ (
    .A(breg_19_bF$buf5),
    .B(areg_31_bF$buf1),
    .C(breg_20_bF$buf4),
    .D(areg_30_bF$buf3),
    .Y(_1354_)
);

NOR2X1 _23018_ (
    .A(_1354_),
    .B(_1353_),
    .Y(_1355_)
);

XOR2X1 _23019_ (
    .A(_1351_),
    .B(_1355_),
    .Y(_1356_)
);

XOR2X1 _23020_ (
    .A(_1356_),
    .B(_1350_),
    .Y(_1357_)
);

INVX1 _23021_ (
    .A(_1357_),
    .Y(_1359_)
);

NAND2X1 _23022_ (
    .A(_1359_),
    .B(_1345_),
    .Y(_1360_)
);

NOR2X1 _23023_ (
    .A(_1359_),
    .B(_1345_),
    .Y(_1361_)
);

INVX2 _23024_ (
    .A(_1361_),
    .Y(_1362_)
);

AND2X2 _23025_ (
    .A(_1362_),
    .B(_1360_),
    .Y(_1363_)
);

NAND3X1 _23026_ (
    .A(_1363_),
    .B(_1340_),
    .C(_1344_),
    .Y(_1364_)
);

AOI21X1 _23027_ (
    .A(_1342_),
    .B(_1343_),
    .C(_1341_),
    .Y(_1365_)
);

AOI21X1 _23028_ (
    .A(_1335_),
    .B(_1339_),
    .C(_1268_),
    .Y(_1366_)
);

INVX2 _23029_ (
    .A(_1363_),
    .Y(_1367_)
);

OAI21X1 _23030_ (
    .A(_1365_),
    .B(_1366_),
    .C(_1367_),
    .Y(_1368_)
);

NAND3X1 _23031_ (
    .A(_1226_),
    .B(_1364_),
    .C(_1368_),
    .Y(_1370_)
);

NOR3X1 _23032_ (
    .A(_1221_),
    .B(_1219_),
    .C(_1222_),
    .Y(_1371_)
);

NAND3X1 _23033_ (
    .A(_1367_),
    .B(_1340_),
    .C(_1344_),
    .Y(_1372_)
);

OAI21X1 _23034_ (
    .A(_1365_),
    .B(_1366_),
    .C(_1363_),
    .Y(_1373_)
);

NAND3X1 _23035_ (
    .A(_1371_),
    .B(_1372_),
    .C(_1373_),
    .Y(_1374_)
);

AOI21X1 _23036_ (
    .A(_1370_),
    .B(_1374_),
    .C(_1267_),
    .Y(_1375_)
);

NAND3X1 _23037_ (
    .A(_1371_),
    .B(_1364_),
    .C(_1368_),
    .Y(_1376_)
);

NAND3X1 _23038_ (
    .A(_1226_),
    .B(_1372_),
    .C(_1373_),
    .Y(_1377_)
);

AOI21X1 _23039_ (
    .A(_1377_),
    .B(_1376_),
    .C(_1266_),
    .Y(_1378_)
);

OAI21X1 _23040_ (
    .A(_1375_),
    .B(_1378_),
    .C(_1265_),
    .Y(_1379_)
);

AOI21X1 _23041_ (
    .A(_1102_),
    .B(_1232_),
    .C(_1225_),
    .Y(_1381_)
);

NAND3X1 _23042_ (
    .A(_1266_),
    .B(_1377_),
    .C(_1376_),
    .Y(_1382_)
);

AOI21X1 _23043_ (
    .A(_1372_),
    .B(_1373_),
    .C(_1226_),
    .Y(_1383_)
);

AOI21X1 _23044_ (
    .A(_1364_),
    .B(_1368_),
    .C(_1371_),
    .Y(_1384_)
);

OAI21X1 _23045_ (
    .A(_1383_),
    .B(_1384_),
    .C(_1267_),
    .Y(_1385_)
);

NAND3X1 _23046_ (
    .A(_1381_),
    .B(_1382_),
    .C(_1385_),
    .Y(_1386_)
);

AOI21X1 _23047_ (
    .A(_1386_),
    .B(_1379_),
    .C(_1264_),
    .Y(_1387_)
);

NAND3X1 _23048_ (
    .A(_1265_),
    .B(_1382_),
    .C(_1385_),
    .Y(_1388_)
);

OAI21X1 _23049_ (
    .A(_1375_),
    .B(_1378_),
    .C(_1381_),
    .Y(_1389_)
);

AOI21X1 _23050_ (
    .A(_1388_),
    .B(_1389_),
    .C(_1263_),
    .Y(_1390_)
);

OAI21X1 _23051_ (
    .A(_1387_),
    .B(_1390_),
    .C(_1262_),
    .Y(_1392_)
);

AOI21X1 _23052_ (
    .A(_1099_),
    .B(_1242_),
    .C(_1248_),
    .Y(_1393_)
);

NAND3X1 _23053_ (
    .A(_1263_),
    .B(_1388_),
    .C(_1389_),
    .Y(_1394_)
);

NAND3X1 _23054_ (
    .A(_1264_),
    .B(_1386_),
    .C(_1379_),
    .Y(_1395_)
);

NAND3X1 _23055_ (
    .A(_1394_),
    .B(_1395_),
    .C(_1393_),
    .Y(_1396_)
);

NAND2X1 _23056_ (
    .A(_1396_),
    .B(_1392_),
    .Y(_1397_)
);

XNOR2X1 _23057_ (
    .A(_1261_),
    .B(_1397_),
    .Y(_0_[50])
);

NAND3X1 _23058_ (
    .A(_1262_),
    .B(_1394_),
    .C(_1395_),
    .Y(_1398_)
);

OAI21X1 _23059_ (
    .A(_1387_),
    .B(_1390_),
    .C(_1393_),
    .Y(_1399_)
);

NAND2X1 _23060_ (
    .A(_1398_),
    .B(_1399_),
    .Y(_1400_)
);

OAI21X1 _23061_ (
    .A(_1261_),
    .B(_1400_),
    .C(_1398_),
    .Y(_1402_)
);

INVX1 _23062_ (
    .A(_1388_),
    .Y(_1403_)
);

AOI21X1 _23063_ (
    .A(_1263_),
    .B(_1389_),
    .C(_1403_),
    .Y(_1404_)
);

OAI21X1 _23064_ (
    .A(_1286_),
    .B(_1287_),
    .C(_1292_),
    .Y(_1405_)
);

AOI21X1 _23065_ (
    .A(_1266_),
    .B(_1377_),
    .C(_1383_),
    .Y(_1406_)
);

NAND2X1 _23066_ (
    .A(_1335_),
    .B(_1340_),
    .Y(_1407_)
);

NAND2X1 _23067_ (
    .A(_1324_),
    .B(_1330_),
    .Y(_1408_)
);

NOR2X1 _23068_ (
    .A(_3958__bF$buf2),
    .B(_7225__bF$buf3),
    .Y(_1409_)
);

INVX1 _23069_ (
    .A(_1409_),
    .Y(_1410_)
);

NOR2X1 _23070_ (
    .A(_1274_),
    .B(_1281_),
    .Y(_1411_)
);

AOI21X1 _23071_ (
    .A(_1273_),
    .B(_1283_),
    .C(_1411_),
    .Y(_1413_)
);

NOR2X1 _23072_ (
    .A(_3961__bF$buf1),
    .B(_6815__bF$buf3),
    .Y(_1414_)
);

OAI21X1 _23073_ (
    .A(_1119_),
    .B(_1275_),
    .C(_1280_),
    .Y(_1415_)
);

NAND2X1 _23074_ (
    .A(areg_23_bF$buf2),
    .B(breg_27_bF$buf3),
    .Y(_1416_)
);

NAND2X1 _23075_ (
    .A(areg_24_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_1417_)
);

OAI21X1 _23076_ (
    .A(_5921__bF$buf1),
    .B(_5668__bF$buf5),
    .C(_1275_),
    .Y(_1418_)
);

OAI21X1 _23077_ (
    .A(_1416_),
    .B(_1417_),
    .C(_1418_),
    .Y(_1419_)
);

OAI21X1 _23078_ (
    .A(_4551__bF$buf1),
    .B(_6427_),
    .C(_1419_),
    .Y(_1420_)
);

NAND2X1 _23079_ (
    .A(areg_22_bF$buf0),
    .B(breg_29_bF$buf0),
    .Y(_1421_)
);

OR2X2 _23080_ (
    .A(_1419_),
    .B(_1421_),
    .Y(_1422_)
);

NAND2X1 _23081_ (
    .A(_1420_),
    .B(_1422_),
    .Y(_1424_)
);

XNOR2X1 _23082_ (
    .A(_1415_),
    .B(_1424_),
    .Y(_1425_)
);

XNOR2X1 _23083_ (
    .A(_1425_),
    .B(_1414_),
    .Y(_1426_)
);

NOR2X1 _23084_ (
    .A(_1413_),
    .B(_1426_),
    .Y(_1427_)
);

INVX1 _23085_ (
    .A(_1413_),
    .Y(_1428_)
);

XOR2X1 _23086_ (
    .A(_1425_),
    .B(_1414_),
    .Y(_1429_)
);

NOR2X1 _23087_ (
    .A(_1428_),
    .B(_1429_),
    .Y(_1430_)
);

OAI21X1 _23088_ (
    .A(_1430_),
    .B(_1427_),
    .C(_1410_),
    .Y(_1431_)
);

NAND2X1 _23089_ (
    .A(_1428_),
    .B(_1429_),
    .Y(_1432_)
);

NAND2X1 _23090_ (
    .A(_1413_),
    .B(_1426_),
    .Y(_1433_)
);

NAND3X1 _23091_ (
    .A(_1409_),
    .B(_1433_),
    .C(_1432_),
    .Y(_1435_)
);

AND2X2 _23092_ (
    .A(_1431_),
    .B(_1435_),
    .Y(_1436_)
);

OAI21X1 _23093_ (
    .A(_1322_),
    .B(_1320_),
    .C(_1316_),
    .Y(_1437_)
);

NAND3X1 _23094_ (
    .A(_1303_),
    .B(_1307_),
    .C(_1309_),
    .Y(_1438_)
);

NAND2X1 _23095_ (
    .A(_1299_),
    .B(_1310_),
    .Y(_1439_)
);

NAND2X1 _23096_ (
    .A(_1438_),
    .B(_1439_),
    .Y(_1440_)
);

OAI21X1 _23097_ (
    .A(_1144_),
    .B(_1301_),
    .C(_1307_),
    .Y(_1441_)
);

OAI21X1 _23098_ (
    .A(_5315__bF$buf0),
    .B(_7100__bF$buf0),
    .C(_1301_),
    .Y(_1442_)
);

NAND2X1 _23099_ (
    .A(breg_25_bF$buf5),
    .B(areg_27_bF$buf3),
    .Y(_1443_)
);

OAI21X1 _23100_ (
    .A(_1305_),
    .B(_1443_),
    .C(_1442_),
    .Y(_1444_)
);

OAI21X1 _23101_ (
    .A(_6300__bF$buf2),
    .B(_5676_),
    .C(_1444_),
    .Y(_1446_)
);

NOR2X1 _23102_ (
    .A(_6300__bF$buf1),
    .B(_5676_),
    .Y(_1447_)
);

NAND2X1 _23103_ (
    .A(breg_24_bF$buf1),
    .B(areg_27_bF$buf2),
    .Y(_1448_)
);

OR2X2 _23104_ (
    .A(_1301_),
    .B(_1448_),
    .Y(_1449_)
);

NAND3X1 _23105_ (
    .A(_1447_),
    .B(_1442_),
    .C(_1449_),
    .Y(_1450_)
);

NAND2X1 _23106_ (
    .A(_1450_),
    .B(_1446_),
    .Y(_1451_)
);

NAND3X1 _23107_ (
    .A(breg_23_bF$buf3),
    .B(areg_27_bF$buf1),
    .C(_1349_),
    .Y(_1452_)
);

OAI21X1 _23108_ (
    .A(_1192_),
    .B(_1348_),
    .C(_1452_),
    .Y(_1453_)
);

XNOR2X1 _23109_ (
    .A(_1453_),
    .B(_1451_),
    .Y(_1454_)
);

XOR2X1 _23110_ (
    .A(_1454_),
    .B(_1441_),
    .Y(_1455_)
);

NAND2X1 _23111_ (
    .A(_1355_),
    .B(_1351_),
    .Y(_1457_)
);

NAND2X1 _23112_ (
    .A(_1350_),
    .B(_1356_),
    .Y(_1458_)
);

NAND2X1 _23113_ (
    .A(_1457_),
    .B(_1458_),
    .Y(_1459_)
);

NAND2X1 _23114_ (
    .A(_1459_),
    .B(_1455_),
    .Y(_1460_)
);

XNOR2X1 _23115_ (
    .A(_1454_),
    .B(_1441_),
    .Y(_1461_)
);

INVX1 _23116_ (
    .A(_1459_),
    .Y(_1462_)
);

NAND2X1 _23117_ (
    .A(_1462_),
    .B(_1461_),
    .Y(_1463_)
);

NAND3X1 _23118_ (
    .A(_1440_),
    .B(_1463_),
    .C(_1460_),
    .Y(_1464_)
);

INVX2 _23119_ (
    .A(_1440_),
    .Y(_1465_)
);

NOR2X1 _23120_ (
    .A(_1462_),
    .B(_1461_),
    .Y(_1466_)
);

NOR2X1 _23121_ (
    .A(_1459_),
    .B(_1455_),
    .Y(_1468_)
);

OAI21X1 _23122_ (
    .A(_1468_),
    .B(_1466_),
    .C(_1465_),
    .Y(_1469_)
);

NAND3X1 _23123_ (
    .A(_1464_),
    .B(_1437_),
    .C(_1469_),
    .Y(_1470_)
);

AOI21X1 _23124_ (
    .A(_1298_),
    .B(_1318_),
    .C(_1321_),
    .Y(_1471_)
);

NAND2X1 _23125_ (
    .A(_1462_),
    .B(_1455_),
    .Y(_1472_)
);

NAND2X1 _23126_ (
    .A(_1459_),
    .B(_1461_),
    .Y(_1473_)
);

AOI21X1 _23127_ (
    .A(_1473_),
    .B(_1472_),
    .C(_1465_),
    .Y(_1474_)
);

AOI21X1 _23128_ (
    .A(_1463_),
    .B(_1460_),
    .C(_1440_),
    .Y(_1475_)
);

OAI21X1 _23129_ (
    .A(_1474_),
    .B(_1475_),
    .C(_1471_),
    .Y(_1476_)
);

NAND3X1 _23130_ (
    .A(_1470_),
    .B(_1476_),
    .C(_1436_),
    .Y(_1477_)
);

NAND2X1 _23131_ (
    .A(_1435_),
    .B(_1431_),
    .Y(_1479_)
);

NOR3X1 _23132_ (
    .A(_1474_),
    .B(_1471_),
    .C(_1475_),
    .Y(_1480_)
);

AOI21X1 _23133_ (
    .A(_1464_),
    .B(_1469_),
    .C(_1437_),
    .Y(_1481_)
);

OAI21X1 _23134_ (
    .A(_1480_),
    .B(_1481_),
    .C(_1479_),
    .Y(_1482_)
);

NAND3X1 _23135_ (
    .A(_1361_),
    .B(_1482_),
    .C(_1477_),
    .Y(_1483_)
);

OAI21X1 _23136_ (
    .A(_1474_),
    .B(_1475_),
    .C(_1437_),
    .Y(_1484_)
);

NAND3X1 _23137_ (
    .A(_1471_),
    .B(_1464_),
    .C(_1469_),
    .Y(_1485_)
);

AOI21X1 _23138_ (
    .A(_1484_),
    .B(_1485_),
    .C(_1479_),
    .Y(_1486_)
);

AOI21X1 _23139_ (
    .A(_1470_),
    .B(_1476_),
    .C(_1436_),
    .Y(_1487_)
);

OAI21X1 _23140_ (
    .A(_1487_),
    .B(_1486_),
    .C(_1362_),
    .Y(_1488_)
);

NAND3X1 _23141_ (
    .A(_1408_),
    .B(_1483_),
    .C(_1488_),
    .Y(_1490_)
);

AND2X2 _23142_ (
    .A(_1330_),
    .B(_1324_),
    .Y(_1491_)
);

NAND3X1 _23143_ (
    .A(_1362_),
    .B(_1482_),
    .C(_1477_),
    .Y(_1492_)
);

OAI21X1 _23144_ (
    .A(_1487_),
    .B(_1486_),
    .C(_1361_),
    .Y(_1493_)
);

NAND3X1 _23145_ (
    .A(_1492_),
    .B(_1493_),
    .C(_1491_),
    .Y(_1494_)
);

NAND2X1 _23146_ (
    .A(breg_23_bF$buf2),
    .B(areg_28_bF$buf5),
    .Y(_1495_)
);

NAND2X1 _23147_ (
    .A(breg_22_bF$buf0),
    .B(areg_30_bF$buf2),
    .Y(_1496_)
);

NOR2X1 _23148_ (
    .A(_1348_),
    .B(_1496_),
    .Y(_1497_)
);

AOI22X1 _23149_ (
    .A(breg_21_bF$buf0),
    .B(areg_30_bF$buf1),
    .C(breg_22_bF$buf4),
    .D(areg_29_bF$buf3),
    .Y(_1498_)
);

NOR2X1 _23150_ (
    .A(_1498_),
    .B(_1497_),
    .Y(_1499_)
);

XNOR2X1 _23151_ (
    .A(_1499_),
    .B(_1495_),
    .Y(_1501_)
);

NOR2X1 _23152_ (
    .A(_1352_),
    .B(_1353_),
    .Y(_1502_)
);

XOR2X1 _23153_ (
    .A(_1501_),
    .B(_1502_),
    .Y(_1503_)
);

AOI21X1 _23154_ (
    .A(_1490_),
    .B(_1494_),
    .C(_1503_),
    .Y(_1504_)
);

AOI21X1 _23155_ (
    .A(_1492_),
    .B(_1493_),
    .C(_1491_),
    .Y(_1505_)
);

AOI21X1 _23156_ (
    .A(_1483_),
    .B(_1488_),
    .C(_1408_),
    .Y(_1506_)
);

INVX1 _23157_ (
    .A(_1503_),
    .Y(_1507_)
);

NOR3X1 _23158_ (
    .A(_1506_),
    .B(_1507_),
    .C(_1505_),
    .Y(_1508_)
);

OAI21X1 _23159_ (
    .A(_1508_),
    .B(_1504_),
    .C(_1364_),
    .Y(_1509_)
);

NOR3X1 _23160_ (
    .A(_1365_),
    .B(_1367_),
    .C(_1366_),
    .Y(_1510_)
);

OAI21X1 _23161_ (
    .A(_1505_),
    .B(_1506_),
    .C(_1507_),
    .Y(_1512_)
);

NAND3X1 _23162_ (
    .A(_1490_),
    .B(_1503_),
    .C(_1494_),
    .Y(_1513_)
);

NAND3X1 _23163_ (
    .A(_1512_),
    .B(_1513_),
    .C(_1510_),
    .Y(_1514_)
);

AOI21X1 _23164_ (
    .A(_1509_),
    .B(_1514_),
    .C(_1407_),
    .Y(_1515_)
);

INVX2 _23165_ (
    .A(_1407_),
    .Y(_1516_)
);

AOI21X1 _23166_ (
    .A(_1512_),
    .B(_1513_),
    .C(_1510_),
    .Y(_1517_)
);

NOR3X1 _23167_ (
    .A(_1364_),
    .B(_1504_),
    .C(_1508_),
    .Y(_1518_)
);

NOR3X1 _23168_ (
    .A(_1517_),
    .B(_1516_),
    .C(_1518_),
    .Y(_1519_)
);

OAI21X1 _23169_ (
    .A(_1519_),
    .B(_1515_),
    .C(_1406_),
    .Y(_1520_)
);

OAI21X1 _23170_ (
    .A(_1384_),
    .B(_1267_),
    .C(_1376_),
    .Y(_1521_)
);

OAI21X1 _23171_ (
    .A(_1518_),
    .B(_1517_),
    .C(_1516_),
    .Y(_1523_)
);

NAND3X1 _23172_ (
    .A(_1407_),
    .B(_1509_),
    .C(_1514_),
    .Y(_1524_)
);

NAND3X1 _23173_ (
    .A(_1521_),
    .B(_1524_),
    .C(_1523_),
    .Y(_1525_)
);

AOI21X1 _23174_ (
    .A(_1525_),
    .B(_1520_),
    .C(_1405_),
    .Y(_1526_)
);

INVX2 _23175_ (
    .A(_1405_),
    .Y(_1527_)
);

AOI21X1 _23176_ (
    .A(_1524_),
    .B(_1523_),
    .C(_1521_),
    .Y(_1528_)
);

NOR3X1 _23177_ (
    .A(_1515_),
    .B(_1406_),
    .C(_1519_),
    .Y(_1529_)
);

NOR3X1 _23178_ (
    .A(_1527_),
    .B(_1528_),
    .C(_1529_),
    .Y(_1530_)
);

OAI21X1 _23179_ (
    .A(_1530_),
    .B(_1526_),
    .C(_1404_),
    .Y(_1531_)
);

NAND2X1 _23180_ (
    .A(_1388_),
    .B(_1394_),
    .Y(_1532_)
);

OAI21X1 _23181_ (
    .A(_1529_),
    .B(_1528_),
    .C(_1527_),
    .Y(_1534_)
);

NAND3X1 _23182_ (
    .A(_1405_),
    .B(_1525_),
    .C(_1520_),
    .Y(_1535_)
);

NAND3X1 _23183_ (
    .A(_1534_),
    .B(_1535_),
    .C(_1532_),
    .Y(_1536_)
);

NAND2X1 _23184_ (
    .A(_1531_),
    .B(_1536_),
    .Y(_1537_)
);

XNOR2X1 _23185_ (
    .A(_1402_),
    .B(_1537_),
    .Y(_0_[51])
);

INVX1 _23186_ (
    .A(_1254_),
    .Y(_1538_)
);

AOI21X1 _23187_ (
    .A(_1255_),
    .B(_1094_),
    .C(_1538_),
    .Y(_1539_)
);

NAND3X1 _23188_ (
    .A(_1531_),
    .B(_1536_),
    .C(_1397_),
    .Y(_1540_)
);

INVX1 _23189_ (
    .A(_1398_),
    .Y(_1541_)
);

NOR3X1 _23190_ (
    .A(_1404_),
    .B(_1526_),
    .C(_1530_),
    .Y(_1542_)
);

AOI21X1 _23191_ (
    .A(_1541_),
    .B(_1531_),
    .C(_1542_),
    .Y(_1544_)
);

OAI21X1 _23192_ (
    .A(_1539_),
    .B(_1540_),
    .C(_1544_),
    .Y(_1545_)
);

NOR2X1 _23193_ (
    .A(_1540_),
    .B(_1258_),
    .Y(_1546_)
);

AOI21X1 _23194_ (
    .A(_1546_),
    .B(_942_),
    .C(_1545_),
    .Y(_1547_)
);

OAI21X1 _23195_ (
    .A(_1528_),
    .B(_1527_),
    .C(_1525_),
    .Y(_1548_)
);

OAI21X1 _23196_ (
    .A(_1430_),
    .B(_1410_),
    .C(_1432_),
    .Y(_1549_)
);

INVX2 _23197_ (
    .A(_1549_),
    .Y(_1550_)
);

OAI21X1 _23198_ (
    .A(_1517_),
    .B(_1516_),
    .C(_1514_),
    .Y(_1551_)
);

NAND2X1 _23199_ (
    .A(_1483_),
    .B(_1490_),
    .Y(_1552_)
);

INVX2 _23200_ (
    .A(_1552_),
    .Y(_1553_)
);

OAI21X1 _23201_ (
    .A(_1479_),
    .B(_1481_),
    .C(_1470_),
    .Y(_1555_)
);

NOR2X1 _23202_ (
    .A(_3961__bF$buf0),
    .B(_7225__bF$buf2),
    .Y(_1556_)
);

NAND3X1 _23203_ (
    .A(_1420_),
    .B(_1422_),
    .C(_1415_),
    .Y(_1557_)
);

NAND2X1 _23204_ (
    .A(_1414_),
    .B(_1425_),
    .Y(_1558_)
);

NAND2X1 _23205_ (
    .A(_1557_),
    .B(_1558_),
    .Y(_1559_)
);

NOR2X1 _23206_ (
    .A(_4551__bF$buf0),
    .B(_6815__bF$buf2),
    .Y(_1560_)
);

OAI21X1 _23207_ (
    .A(_1416_),
    .B(_1417_),
    .C(_1422_),
    .Y(_1561_)
);

NAND2X1 _23208_ (
    .A(areg_23_bF$buf1),
    .B(breg_29_bF$buf4),
    .Y(_1562_)
);

NAND2X1 _23209_ (
    .A(areg_24_bF$buf1),
    .B(breg_27_bF$buf2),
    .Y(_1563_)
);

NAND2X1 _23210_ (
    .A(areg_25_bF$buf0),
    .B(breg_28_bF$buf1),
    .Y(_1564_)
);

OAI21X1 _23211_ (
    .A(_6300__bF$buf0),
    .B(_5668__bF$buf4),
    .C(_1417_),
    .Y(_1566_)
);

OAI21X1 _23212_ (
    .A(_1563_),
    .B(_1564_),
    .C(_1566_),
    .Y(_1567_)
);

XNOR2X1 _23213_ (
    .A(_1567_),
    .B(_1562_),
    .Y(_1568_)
);

XNOR2X1 _23214_ (
    .A(_1561_),
    .B(_1568_),
    .Y(_1569_)
);

XNOR2X1 _23215_ (
    .A(_1569_),
    .B(_1560_),
    .Y(_1570_)
);

XNOR2X1 _23216_ (
    .A(_1559_),
    .B(_1570_),
    .Y(_1571_)
);

XOR2X1 _23217_ (
    .A(_1571_),
    .B(_1556_),
    .Y(_1572_)
);

AOI21X1 _23218_ (
    .A(_1440_),
    .B(_1463_),
    .C(_1466_),
    .Y(_1573_)
);

NAND3X1 _23219_ (
    .A(_1446_),
    .B(_1450_),
    .C(_1453_),
    .Y(_1574_)
);

NAND2X1 _23220_ (
    .A(_1441_),
    .B(_1454_),
    .Y(_1575_)
);

NAND2X1 _23221_ (
    .A(_1574_),
    .B(_1575_),
    .Y(_1576_)
);

OAI21X1 _23222_ (
    .A(_1305_),
    .B(_1443_),
    .C(_1450_),
    .Y(_1577_)
);

NAND2X1 _23223_ (
    .A(breg_25_bF$buf4),
    .B(areg_28_bF$buf4),
    .Y(_1578_)
);

OAI21X1 _23224_ (
    .A(_5315__bF$buf4),
    .B(_7520__bF$buf3),
    .C(_1443_),
    .Y(_1579_)
);

OAI21X1 _23225_ (
    .A(_1448_),
    .B(_1578_),
    .C(_1579_),
    .Y(_1580_)
);

OAI21X1 _23226_ (
    .A(_6686__bF$buf2),
    .B(_5676_),
    .C(_1580_),
    .Y(_1581_)
);

NOR2X1 _23227_ (
    .A(_6686__bF$buf1),
    .B(_5676_),
    .Y(_1582_)
);

OR2X2 _23228_ (
    .A(_1448_),
    .B(_1578_),
    .Y(_1583_)
);

NAND3X1 _23229_ (
    .A(_1582_),
    .B(_1579_),
    .C(_1583_),
    .Y(_1584_)
);

NAND2X1 _23230_ (
    .A(_1584_),
    .B(_1581_),
    .Y(_1585_)
);

OAI22X1 _23231_ (
    .A(_1348_),
    .B(_1496_),
    .C(_1498_),
    .D(_1495_),
    .Y(_1588_)
);

XNOR2X1 _23232_ (
    .A(_1585_),
    .B(_1588_),
    .Y(_1589_)
);

XOR2X1 _23233_ (
    .A(_1589_),
    .B(_1577_),
    .Y(_1590_)
);

AOI21X1 _23234_ (
    .A(_1502_),
    .B(_1501_),
    .C(_1353_),
    .Y(_1591_)
);

INVX1 _23235_ (
    .A(_1591_),
    .Y(_1592_)
);

NAND2X1 _23236_ (
    .A(_1592_),
    .B(_1590_),
    .Y(_1593_)
);

XNOR2X1 _23237_ (
    .A(_1589_),
    .B(_1577_),
    .Y(_1594_)
);

NAND2X1 _23238_ (
    .A(_1591_),
    .B(_1594_),
    .Y(_1595_)
);

NAND3X1 _23239_ (
    .A(_1576_),
    .B(_1595_),
    .C(_1593_),
    .Y(_1596_)
);

INVX1 _23240_ (
    .A(_1576_),
    .Y(_1597_)
);

NOR2X1 _23241_ (
    .A(_1591_),
    .B(_1594_),
    .Y(_1599_)
);

NOR2X1 _23242_ (
    .A(_1592_),
    .B(_1590_),
    .Y(_1600_)
);

OAI21X1 _23243_ (
    .A(_1600_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1601_)
);

NAND2X1 _23244_ (
    .A(_1596_),
    .B(_1601_),
    .Y(_1602_)
);

NAND2X1 _23245_ (
    .A(_1573_),
    .B(_1602_),
    .Y(_1603_)
);

OAI21X1 _23246_ (
    .A(_1468_),
    .B(_1465_),
    .C(_1460_),
    .Y(_1604_)
);

NAND3X1 _23247_ (
    .A(_1596_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1605_)
);

NAND3X1 _23248_ (
    .A(_1603_),
    .B(_1605_),
    .C(_1572_),
    .Y(_1606_)
);

XNOR2X1 _23249_ (
    .A(_1571_),
    .B(_1556_),
    .Y(_1607_)
);

AOI21X1 _23250_ (
    .A(_1596_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1608_)
);

NOR2X1 _23251_ (
    .A(_1573_),
    .B(_1602_),
    .Y(_1610_)
);

OAI21X1 _23252_ (
    .A(_1610_),
    .B(_1608_),
    .C(_1607_),
    .Y(_1611_)
);

NAND3X1 _23253_ (
    .A(_1555_),
    .B(_1611_),
    .C(_1606_),
    .Y(_1612_)
);

AOI21X1 _23254_ (
    .A(_1476_),
    .B(_1436_),
    .C(_1480_),
    .Y(_1613_)
);

OAI21X1 _23255_ (
    .A(_1610_),
    .B(_1608_),
    .C(_1572_),
    .Y(_1614_)
);

NAND3X1 _23256_ (
    .A(_1603_),
    .B(_1605_),
    .C(_1607_),
    .Y(_1615_)
);

NAND3X1 _23257_ (
    .A(_1613_),
    .B(_1614_),
    .C(_1615_),
    .Y(_1616_)
);

NOR2X1 _23258_ (
    .A(_5369_),
    .B(_9153_),
    .Y(_1617_)
);

NAND2X1 _23259_ (
    .A(breg_21_bF$buf4),
    .B(areg_31_bF$buf0),
    .Y(_1618_)
);

XOR2X1 _23260_ (
    .A(_1496_),
    .B(_1618_),
    .Y(_1619_)
);

XOR2X1 _23261_ (
    .A(_1619_),
    .B(_1617_),
    .Y(_1621_)
);

NAND3X1 _23262_ (
    .A(_1621_),
    .B(_1612_),
    .C(_1616_),
    .Y(_1622_)
);

AOI21X1 _23263_ (
    .A(_1614_),
    .B(_1615_),
    .C(_1613_),
    .Y(_1623_)
);

AOI21X1 _23264_ (
    .A(_1611_),
    .B(_1606_),
    .C(_1555_),
    .Y(_1624_)
);

INVX1 _23265_ (
    .A(_1621_),
    .Y(_1625_)
);

OAI21X1 _23266_ (
    .A(_1624_),
    .B(_1623_),
    .C(_1625_),
    .Y(_1626_)
);

NAND2X1 _23267_ (
    .A(_1622_),
    .B(_1626_),
    .Y(_1627_)
);

NOR2X1 _23268_ (
    .A(_1627_),
    .B(_1513_),
    .Y(_1628_)
);

AND2X2 _23269_ (
    .A(_1513_),
    .B(_1627_),
    .Y(_1629_)
);

NOR3X1 _23270_ (
    .A(_1628_),
    .B(_1553_),
    .C(_1629_),
    .Y(_1630_)
);

OR2X2 _23271_ (
    .A(_1513_),
    .B(_1627_),
    .Y(_1632_)
);

NAND2X1 _23272_ (
    .A(_1627_),
    .B(_1513_),
    .Y(_1633_)
);

AOI21X1 _23273_ (
    .A(_1633_),
    .B(_1632_),
    .C(_1552_),
    .Y(_1634_)
);

OAI21X1 _23274_ (
    .A(_1630_),
    .B(_1634_),
    .C(_1551_),
    .Y(_1635_)
);

AOI21X1 _23275_ (
    .A(_1407_),
    .B(_1509_),
    .C(_1518_),
    .Y(_1636_)
);

NAND3X1 _23276_ (
    .A(_1552_),
    .B(_1633_),
    .C(_1632_),
    .Y(_1637_)
);

OAI21X1 _23277_ (
    .A(_1629_),
    .B(_1628_),
    .C(_1553_),
    .Y(_1638_)
);

NAND3X1 _23278_ (
    .A(_1637_),
    .B(_1638_),
    .C(_1636_),
    .Y(_1639_)
);

AOI21X1 _23279_ (
    .A(_1635_),
    .B(_1639_),
    .C(_1550_),
    .Y(_1640_)
);

NAND3X1 _23280_ (
    .A(_1637_),
    .B(_1638_),
    .C(_1551_),
    .Y(_1641_)
);

OAI21X1 _23281_ (
    .A(_1630_),
    .B(_1634_),
    .C(_1636_),
    .Y(_1643_)
);

AOI21X1 _23282_ (
    .A(_1643_),
    .B(_1641_),
    .C(_1549_),
    .Y(_1644_)
);

OAI21X1 _23283_ (
    .A(_1644_),
    .B(_1640_),
    .C(_1548_),
    .Y(_1645_)
);

AOI21X1 _23284_ (
    .A(_1405_),
    .B(_1520_),
    .C(_1529_),
    .Y(_1646_)
);

NAND3X1 _23285_ (
    .A(_1549_),
    .B(_1643_),
    .C(_1641_),
    .Y(_1647_)
);

NOR3X1 _23286_ (
    .A(_1630_),
    .B(_1634_),
    .C(_1636_),
    .Y(_1648_)
);

AOI21X1 _23287_ (
    .A(_1637_),
    .B(_1638_),
    .C(_1551_),
    .Y(_1649_)
);

OAI21X1 _23288_ (
    .A(_1648_),
    .B(_1649_),
    .C(_1550_),
    .Y(_1650_)
);

NAND3X1 _23289_ (
    .A(_1647_),
    .B(_1650_),
    .C(_1646_),
    .Y(_1651_)
);

NAND2X1 _23290_ (
    .A(_1645_),
    .B(_1651_),
    .Y(_1652_)
);

XNOR2X1 _23291_ (
    .A(_1547_),
    .B(_1652_),
    .Y(_0_[52])
);

NAND3X1 _23292_ (
    .A(_1647_),
    .B(_1548_),
    .C(_1650_),
    .Y(_1654_)
);

INVX1 _23293_ (
    .A(_1652_),
    .Y(_1655_)
);

OAI21X1 _23294_ (
    .A(_1547_),
    .B(_1655_),
    .C(_1654_),
    .Y(_1656_)
);

AOI21X1 _23295_ (
    .A(_1549_),
    .B(_1643_),
    .C(_1648_),
    .Y(_1657_)
);

AOI21X1 _23296_ (
    .A(_1557_),
    .B(_1558_),
    .C(_1570_),
    .Y(_1658_)
);

AND2X2 _23297_ (
    .A(_1571_),
    .B(_1556_),
    .Y(_1659_)
);

NOR2X1 _23298_ (
    .A(_1658_),
    .B(_1659_),
    .Y(_1660_)
);

INVX2 _23299_ (
    .A(_1660_),
    .Y(_1661_)
);

AOI21X1 _23300_ (
    .A(_1552_),
    .B(_1633_),
    .C(_1628_),
    .Y(_1662_)
);

OAI21X1 _23301_ (
    .A(_1607_),
    .B(_1608_),
    .C(_1605_),
    .Y(_1664_)
);

NOR2X1 _23302_ (
    .A(_4551__bF$buf4),
    .B(_7225__bF$buf1),
    .Y(_1665_)
);

INVX1 _23303_ (
    .A(_1665_),
    .Y(_1666_)
);

OAI21X1 _23304_ (
    .A(_4541__bF$buf2),
    .B(_6427_),
    .C(_1567_),
    .Y(_1667_)
);

OR2X2 _23305_ (
    .A(_1567_),
    .B(_1562_),
    .Y(_1668_)
);

NAND3X1 _23306_ (
    .A(_1667_),
    .B(_1668_),
    .C(_1561_),
    .Y(_1669_)
);

NAND2X1 _23307_ (
    .A(_1560_),
    .B(_1569_),
    .Y(_1670_)
);

NAND2X1 _23308_ (
    .A(_1669_),
    .B(_1670_),
    .Y(_1671_)
);

NOR2X1 _23309_ (
    .A(_4541__bF$buf1),
    .B(_6815__bF$buf1),
    .Y(_1672_)
);

INVX1 _23310_ (
    .A(_1562_),
    .Y(_1673_)
);

NAND2X1 _23311_ (
    .A(areg_25_bF$buf4),
    .B(breg_27_bF$buf1),
    .Y(_1675_)
);

NOR2X1 _23312_ (
    .A(_1417_),
    .B(_1675_),
    .Y(_1676_)
);

AOI21X1 _23313_ (
    .A(_1673_),
    .B(_1566_),
    .C(_1676_),
    .Y(_1677_)
);

NAND2X1 _23314_ (
    .A(areg_24_bF$buf0),
    .B(breg_29_bF$buf3),
    .Y(_1678_)
);

NAND2X1 _23315_ (
    .A(areg_26_bF$buf4),
    .B(breg_28_bF$buf0),
    .Y(_1679_)
);

OAI21X1 _23316_ (
    .A(_6686__bF$buf0),
    .B(_5668__bF$buf3),
    .C(_1564_),
    .Y(_1680_)
);

OAI21X1 _23317_ (
    .A(_1675_),
    .B(_1679_),
    .C(_1680_),
    .Y(_1681_)
);

XOR2X1 _23318_ (
    .A(_1681_),
    .B(_1678_),
    .Y(_1682_)
);

XNOR2X1 _23319_ (
    .A(_1682_),
    .B(_1677_),
    .Y(_1683_)
);

XOR2X1 _23320_ (
    .A(_1683_),
    .B(_1672_),
    .Y(_1684_)
);

NOR2X1 _23321_ (
    .A(_1684_),
    .B(_1671_),
    .Y(_1686_)
);

AND2X2 _23322_ (
    .A(_1671_),
    .B(_1684_),
    .Y(_1687_)
);

OAI21X1 _23323_ (
    .A(_1687_),
    .B(_1686_),
    .C(_1666_),
    .Y(_1688_)
);

OR2X2 _23324_ (
    .A(_1671_),
    .B(_1684_),
    .Y(_1689_)
);

NAND2X1 _23325_ (
    .A(_1684_),
    .B(_1671_),
    .Y(_1690_)
);

NAND3X1 _23326_ (
    .A(_1665_),
    .B(_1690_),
    .C(_1689_),
    .Y(_1691_)
);

NAND2X1 _23327_ (
    .A(_1688_),
    .B(_1691_),
    .Y(_1692_)
);

INVX2 _23328_ (
    .A(_1692_),
    .Y(_1693_)
);

OAI21X1 _23329_ (
    .A(_1597_),
    .B(_1600_),
    .C(_1593_),
    .Y(_1694_)
);

NAND3X1 _23330_ (
    .A(_1584_),
    .B(_1588_),
    .C(_1581_),
    .Y(_1695_)
);

NAND2X1 _23331_ (
    .A(_1577_),
    .B(_1589_),
    .Y(_1697_)
);

NAND2X1 _23332_ (
    .A(_1695_),
    .B(_1697_),
    .Y(_1698_)
);

INVX1 _23333_ (
    .A(_1698_),
    .Y(_1699_)
);

INVX1 _23334_ (
    .A(_1582_),
    .Y(_1700_)
);

OAI21X1 _23335_ (
    .A(_1580_),
    .B(_1700_),
    .C(_1583_),
    .Y(_1701_)
);

NAND2X1 _23336_ (
    .A(breg_26_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_1702_)
);

NAND2X1 _23337_ (
    .A(breg_24_bF$buf0),
    .B(areg_29_bF$buf2),
    .Y(_1703_)
);

NOR2X1 _23338_ (
    .A(_1578_),
    .B(_1703_),
    .Y(_1704_)
);

AND2X2 _23339_ (
    .A(_1578_),
    .B(_1703_),
    .Y(_1705_)
);

OR2X2 _23340_ (
    .A(_1705_),
    .B(_1704_),
    .Y(_1706_)
);

XNOR2X1 _23341_ (
    .A(_1706_),
    .B(_1702_),
    .Y(_1708_)
);

NAND2X1 _23342_ (
    .A(_1617_),
    .B(_1619_),
    .Y(_1709_)
);

OAI21X1 _23343_ (
    .A(_1496_),
    .B(_1618_),
    .C(_1709_),
    .Y(_1710_)
);

XNOR2X1 _23344_ (
    .A(_1708_),
    .B(_1710_),
    .Y(_1711_)
);

NOR2X1 _23345_ (
    .A(_1701_),
    .B(_1711_),
    .Y(_1712_)
);

INVX1 _23346_ (
    .A(_1701_),
    .Y(_1713_)
);

XOR2X1 _23347_ (
    .A(_1708_),
    .B(_1710_),
    .Y(_1714_)
);

NOR2X1 _23348_ (
    .A(_1713_),
    .B(_1714_),
    .Y(_1715_)
);

OAI21X1 _23349_ (
    .A(_1712_),
    .B(_1715_),
    .C(_1699_),
    .Y(_1716_)
);

NOR2X1 _23350_ (
    .A(_1712_),
    .B(_1715_),
    .Y(_1717_)
);

NAND2X1 _23351_ (
    .A(_1698_),
    .B(_1717_),
    .Y(_1719_)
);

NAND2X1 _23352_ (
    .A(_1716_),
    .B(_1719_),
    .Y(_1720_)
);

XNOR2X1 _23353_ (
    .A(_1720_),
    .B(_1694_),
    .Y(_1721_)
);

NAND2X1 _23354_ (
    .A(_1693_),
    .B(_1721_),
    .Y(_1722_)
);

AND2X2 _23355_ (
    .A(_1719_),
    .B(_1716_),
    .Y(_1723_)
);

NOR2X1 _23356_ (
    .A(_1694_),
    .B(_1723_),
    .Y(_1724_)
);

AOI21X1 _23357_ (
    .A(_1593_),
    .B(_1596_),
    .C(_1720_),
    .Y(_1725_)
);

OAI21X1 _23358_ (
    .A(_1724_),
    .B(_1725_),
    .C(_1692_),
    .Y(_1726_)
);

NAND3X1 _23359_ (
    .A(_1722_),
    .B(_1726_),
    .C(_1664_),
    .Y(_1727_)
);

AOI21X1 _23360_ (
    .A(_1603_),
    .B(_1572_),
    .C(_1610_),
    .Y(_1728_)
);

OAI21X1 _23361_ (
    .A(_1724_),
    .B(_1725_),
    .C(_1693_),
    .Y(_1730_)
);

NAND2X1 _23362_ (
    .A(_1692_),
    .B(_1721_),
    .Y(_1731_)
);

NAND3X1 _23363_ (
    .A(_1730_),
    .B(_1731_),
    .C(_1728_),
    .Y(_1732_)
);

NAND2X1 _23364_ (
    .A(breg_23_bF$buf1),
    .B(areg_31_bF$buf4),
    .Y(_1733_)
);

OAI22X1 _23365_ (
    .A(_4069_),
    .B(_8773_),
    .C(_5369_),
    .D(_8759_),
    .Y(_1734_)
);

OAI21X1 _23366_ (
    .A(_1496_),
    .B(_1733_),
    .C(_1734_),
    .Y(_1735_)
);

INVX1 _23367_ (
    .A(_1735_),
    .Y(_1736_)
);

AOI21X1 _23368_ (
    .A(_1727_),
    .B(_1732_),
    .C(_1736_),
    .Y(_1737_)
);

AOI21X1 _23369_ (
    .A(_1731_),
    .B(_1730_),
    .C(_1728_),
    .Y(_1738_)
);

AOI21X1 _23370_ (
    .A(_1726_),
    .B(_1722_),
    .C(_1664_),
    .Y(_1739_)
);

NOR3X1 _23371_ (
    .A(_1739_),
    .B(_1735_),
    .C(_1738_),
    .Y(_1741_)
);

OAI21X1 _23372_ (
    .A(_1741_),
    .B(_1737_),
    .C(_1622_),
    .Y(_1742_)
);

INVX1 _23373_ (
    .A(_1622_),
    .Y(_1743_)
);

OAI21X1 _23374_ (
    .A(_1738_),
    .B(_1739_),
    .C(_1735_),
    .Y(_1744_)
);

NAND3X1 _23375_ (
    .A(_1736_),
    .B(_1727_),
    .C(_1732_),
    .Y(_1745_)
);

NAND3X1 _23376_ (
    .A(_1745_),
    .B(_1744_),
    .C(_1743_),
    .Y(_1746_)
);

AOI21X1 _23377_ (
    .A(_1742_),
    .B(_1746_),
    .C(_1623_),
    .Y(_1747_)
);

NOR2X1 _23378_ (
    .A(_1623_),
    .B(_1624_),
    .Y(_1748_)
);

AOI22X1 _23379_ (
    .A(_1748_),
    .B(_1621_),
    .C(_1744_),
    .D(_1745_),
    .Y(_1749_)
);

NOR3X1 _23380_ (
    .A(_1622_),
    .B(_1737_),
    .C(_1741_),
    .Y(_1750_)
);

NOR3X1 _23381_ (
    .A(_1612_),
    .B(_1749_),
    .C(_1750_),
    .Y(_1752_)
);

OAI21X1 _23382_ (
    .A(_1752_),
    .B(_1747_),
    .C(_1662_),
    .Y(_1753_)
);

OAI21X1 _23383_ (
    .A(_1629_),
    .B(_1553_),
    .C(_1632_),
    .Y(_1754_)
);

OAI21X1 _23384_ (
    .A(_1750_),
    .B(_1749_),
    .C(_1612_),
    .Y(_1755_)
);

NAND3X1 _23385_ (
    .A(_1623_),
    .B(_1742_),
    .C(_1746_),
    .Y(_1756_)
);

NAND3X1 _23386_ (
    .A(_1755_),
    .B(_1756_),
    .C(_1754_),
    .Y(_1757_)
);

AOI21X1 _23387_ (
    .A(_1753_),
    .B(_1757_),
    .C(_1661_),
    .Y(_1758_)
);

AOI21X1 _23388_ (
    .A(_1755_),
    .B(_1756_),
    .C(_1754_),
    .Y(_1759_)
);

NOR3X1 _23389_ (
    .A(_1747_),
    .B(_1752_),
    .C(_1662_),
    .Y(_1760_)
);

NOR3X1 _23390_ (
    .A(_1759_),
    .B(_1660_),
    .C(_1760_),
    .Y(_1761_)
);

OAI21X1 _23391_ (
    .A(_1761_),
    .B(_1758_),
    .C(_1657_),
    .Y(_1763_)
);

OAI21X1 _23392_ (
    .A(_1649_),
    .B(_1550_),
    .C(_1641_),
    .Y(_1764_)
);

OAI21X1 _23393_ (
    .A(_1760_),
    .B(_1759_),
    .C(_1660_),
    .Y(_1765_)
);

NAND3X1 _23394_ (
    .A(_1661_),
    .B(_1753_),
    .C(_1757_),
    .Y(_1766_)
);

NAND3X1 _23395_ (
    .A(_1765_),
    .B(_1766_),
    .C(_1764_),
    .Y(_1767_)
);

NAND2X1 _23396_ (
    .A(_1767_),
    .B(_1763_),
    .Y(_1768_)
);

XNOR2X1 _23397_ (
    .A(_1656_),
    .B(_1768_),
    .Y(_0_[53])
);

NAND2X1 _23398_ (
    .A(_1767_),
    .B(_1654_),
    .Y(_1769_)
);

NAND2X1 _23399_ (
    .A(_1763_),
    .B(_1769_),
    .Y(_1770_)
);

NOR2X1 _23400_ (
    .A(_1768_),
    .B(_1655_),
    .Y(_1771_)
);

INVX1 _23401_ (
    .A(_1771_),
    .Y(_1773_)
);

OAI21X1 _23402_ (
    .A(_1547_),
    .B(_1773_),
    .C(_1770_),
    .Y(_1774_)
);

AOI21X1 _23403_ (
    .A(_1661_),
    .B(_1753_),
    .C(_1760_),
    .Y(_1775_)
);

INVX1 _23404_ (
    .A(_1775_),
    .Y(_1776_)
);

OAI21X1 _23405_ (
    .A(_1686_),
    .B(_1666_),
    .C(_1690_),
    .Y(_1777_)
);

OAI21X1 _23406_ (
    .A(_1749_),
    .B(_1612_),
    .C(_1746_),
    .Y(_1778_)
);

INVX1 _23407_ (
    .A(_1733_),
    .Y(_1779_)
);

INVX1 _23408_ (
    .A(_1725_),
    .Y(_1780_)
);

OAI21X1 _23409_ (
    .A(_1724_),
    .B(_1692_),
    .C(_1780_),
    .Y(_1781_)
);

NOR2X1 _23410_ (
    .A(_4541__bF$buf0),
    .B(_7225__bF$buf0),
    .Y(_1782_)
);

INVX1 _23411_ (
    .A(_1677_),
    .Y(_1784_)
);

NAND2X1 _23412_ (
    .A(_1784_),
    .B(_1682_),
    .Y(_1785_)
);

NAND2X1 _23413_ (
    .A(_1672_),
    .B(_1683_),
    .Y(_1786_)
);

NAND2X1 _23414_ (
    .A(_1785_),
    .B(_1786_),
    .Y(_1787_)
);

NOR2X1 _23415_ (
    .A(_5921__bF$buf0),
    .B(_6815__bF$buf0),
    .Y(_1788_)
);

NAND2X1 _23416_ (
    .A(areg_26_bF$buf3),
    .B(breg_27_bF$buf0),
    .Y(_1789_)
);

NOR2X1 _23417_ (
    .A(_1564_),
    .B(_1789_),
    .Y(_1790_)
);

NOR2X1 _23418_ (
    .A(_1678_),
    .B(_1681_),
    .Y(_1791_)
);

NOR2X1 _23419_ (
    .A(_1790_),
    .B(_1791_),
    .Y(_1792_)
);

NAND2X1 _23420_ (
    .A(areg_25_bF$buf3),
    .B(breg_29_bF$buf2),
    .Y(_1793_)
);

NAND2X1 _23421_ (
    .A(areg_27_bF$buf5),
    .B(breg_28_bF$buf5),
    .Y(_1795_)
);

OAI21X1 _23422_ (
    .A(_7100__bF$buf3),
    .B(_5668__bF$buf2),
    .C(_1679_),
    .Y(_1796_)
);

OAI21X1 _23423_ (
    .A(_1789_),
    .B(_1795_),
    .C(_1796_),
    .Y(_1797_)
);

XNOR2X1 _23424_ (
    .A(_1797_),
    .B(_1793_),
    .Y(_1798_)
);

XOR2X1 _23425_ (
    .A(_1792_),
    .B(_1798_),
    .Y(_1799_)
);

XNOR2X1 _23426_ (
    .A(_1799_),
    .B(_1788_),
    .Y(_1800_)
);

XNOR2X1 _23427_ (
    .A(_1800_),
    .B(_1787_),
    .Y(_1801_)
);

XOR2X1 _23428_ (
    .A(_1801_),
    .B(_1782_),
    .Y(_1802_)
);

INVX1 _23429_ (
    .A(_1708_),
    .Y(_1803_)
);

NAND2X1 _23430_ (
    .A(_1710_),
    .B(_1803_),
    .Y(_1804_)
);

OAI21X1 _23431_ (
    .A(_1714_),
    .B(_1713_),
    .C(_1804_),
    .Y(_1806_)
);

INVX1 _23432_ (
    .A(_1704_),
    .Y(_1807_)
);

OAI21X1 _23433_ (
    .A(_1705_),
    .B(_1702_),
    .C(_1807_),
    .Y(_1808_)
);

NOR2X1 _23434_ (
    .A(_1496_),
    .B(_1733_),
    .Y(_1809_)
);

NAND2X1 _23435_ (
    .A(breg_26_bF$buf2),
    .B(areg_28_bF$buf3),
    .Y(_1810_)
);

NAND2X1 _23436_ (
    .A(breg_25_bF$buf3),
    .B(areg_30_bF$buf0),
    .Y(_1811_)
);

NAND2X1 _23437_ (
    .A(breg_24_bF$buf5),
    .B(areg_30_bF$buf5),
    .Y(_1812_)
);

OAI21X1 _23438_ (
    .A(_5318_),
    .B(_9153_),
    .C(_1812_),
    .Y(_1813_)
);

OAI21X1 _23439_ (
    .A(_1703_),
    .B(_1811_),
    .C(_1813_),
    .Y(_1814_)
);

XOR2X1 _23440_ (
    .A(_1814_),
    .B(_1810_),
    .Y(_1815_)
);

XOR2X1 _23441_ (
    .A(_1815_),
    .B(_1809_),
    .Y(_1817_)
);

XOR2X1 _23442_ (
    .A(_1817_),
    .B(_1808_),
    .Y(_1818_)
);

XNOR2X1 _23443_ (
    .A(_1818_),
    .B(_1806_),
    .Y(_1819_)
);

NAND2X1 _23444_ (
    .A(_1719_),
    .B(_1819_),
    .Y(_1820_)
);

XOR2X1 _23445_ (
    .A(_1818_),
    .B(_1806_),
    .Y(_1821_)
);

NAND3X1 _23446_ (
    .A(_1698_),
    .B(_1717_),
    .C(_1821_),
    .Y(_1822_)
);

AND2X2 _23447_ (
    .A(_1822_),
    .B(_1820_),
    .Y(_1823_)
);

NAND2X1 _23448_ (
    .A(_1802_),
    .B(_1823_),
    .Y(_1824_)
);

XNOR2X1 _23449_ (
    .A(_1801_),
    .B(_1782_),
    .Y(_1825_)
);

NAND2X1 _23450_ (
    .A(_1820_),
    .B(_1822_),
    .Y(_1826_)
);

NAND2X1 _23451_ (
    .A(_1825_),
    .B(_1826_),
    .Y(_1828_)
);

NAND3X1 _23452_ (
    .A(_1824_),
    .B(_1828_),
    .C(_1781_),
    .Y(_1829_)
);

AOI21X1 _23453_ (
    .A(_1693_),
    .B(_1721_),
    .C(_1725_),
    .Y(_1830_)
);

NOR2X1 _23454_ (
    .A(_1825_),
    .B(_1826_),
    .Y(_1831_)
);

NOR2X1 _23455_ (
    .A(_1802_),
    .B(_1823_),
    .Y(_1832_)
);

OAI21X1 _23456_ (
    .A(_1832_),
    .B(_1831_),
    .C(_1830_),
    .Y(_1833_)
);

NAND3X1 _23457_ (
    .A(_1779_),
    .B(_1829_),
    .C(_1833_),
    .Y(_1834_)
);

NAND2X1 _23458_ (
    .A(_1802_),
    .B(_1826_),
    .Y(_1835_)
);

NAND2X1 _23459_ (
    .A(_1825_),
    .B(_1823_),
    .Y(_1836_)
);

AOI21X1 _23460_ (
    .A(_1835_),
    .B(_1836_),
    .C(_1830_),
    .Y(_1837_)
);

AOI21X1 _23461_ (
    .A(_1828_),
    .B(_1824_),
    .C(_1781_),
    .Y(_1839_)
);

OAI21X1 _23462_ (
    .A(_1837_),
    .B(_1839_),
    .C(_1733_),
    .Y(_1840_)
);

AOI21X1 _23463_ (
    .A(_1834_),
    .B(_1840_),
    .C(_1741_),
    .Y(_1841_)
);

NOR3X1 _23464_ (
    .A(_1733_),
    .B(_1839_),
    .C(_1837_),
    .Y(_1842_)
);

AOI21X1 _23465_ (
    .A(_1829_),
    .B(_1833_),
    .C(_1779_),
    .Y(_1843_)
);

NOR3X1 _23466_ (
    .A(_1843_),
    .B(_1745_),
    .C(_1842_),
    .Y(_1844_)
);

OAI21X1 _23467_ (
    .A(_1844_),
    .B(_1841_),
    .C(_1727_),
    .Y(_1845_)
);

OAI21X1 _23468_ (
    .A(_1842_),
    .B(_1843_),
    .C(_1745_),
    .Y(_1846_)
);

NAND3X1 _23469_ (
    .A(_1834_),
    .B(_1840_),
    .C(_1741_),
    .Y(_1847_)
);

NAND3X1 _23470_ (
    .A(_1738_),
    .B(_1847_),
    .C(_1846_),
    .Y(_1848_)
);

NAND3X1 _23471_ (
    .A(_1848_),
    .B(_1778_),
    .C(_1845_),
    .Y(_1850_)
);

AOI21X1 _23472_ (
    .A(_1623_),
    .B(_1742_),
    .C(_1750_),
    .Y(_1851_)
);

AOI21X1 _23473_ (
    .A(_1847_),
    .B(_1846_),
    .C(_1738_),
    .Y(_1852_)
);

NOR3X1 _23474_ (
    .A(_1841_),
    .B(_1727_),
    .C(_1844_),
    .Y(_1853_)
);

OAI21X1 _23475_ (
    .A(_1853_),
    .B(_1852_),
    .C(_1851_),
    .Y(_1854_)
);

NAND3X1 _23476_ (
    .A(_1777_),
    .B(_1850_),
    .C(_1854_),
    .Y(_1855_)
);

INVX1 _23477_ (
    .A(_1777_),
    .Y(_1856_)
);

NOR3X1 _23478_ (
    .A(_1851_),
    .B(_1852_),
    .C(_1853_),
    .Y(_1857_)
);

AOI21X1 _23479_ (
    .A(_1848_),
    .B(_1845_),
    .C(_1778_),
    .Y(_1858_)
);

OAI21X1 _23480_ (
    .A(_1857_),
    .B(_1858_),
    .C(_1856_),
    .Y(_1859_)
);

NAND2X1 _23481_ (
    .A(_1855_),
    .B(_1859_),
    .Y(_1861_)
);

NAND2X1 _23482_ (
    .A(_1776_),
    .B(_1861_),
    .Y(_1862_)
);

NAND3X1 _23483_ (
    .A(_1855_),
    .B(_1859_),
    .C(_1775_),
    .Y(_1863_)
);

NAND2X1 _23484_ (
    .A(_1863_),
    .B(_1862_),
    .Y(_1864_)
);

XOR2X1 _23485_ (
    .A(_1774_),
    .B(_1864_),
    .Y(_0_[54])
);

NOR2X1 _23486_ (
    .A(_1775_),
    .B(_1861_),
    .Y(_1865_)
);

AOI21X1 _23487_ (
    .A(_1864_),
    .B(_1774_),
    .C(_1865_),
    .Y(_1866_)
);

AOI21X1 _23488_ (
    .A(_1777_),
    .B(_1854_),
    .C(_1857_),
    .Y(_1867_)
);

INVX1 _23489_ (
    .A(_1800_),
    .Y(_1868_)
);

NAND2X1 _23490_ (
    .A(_1787_),
    .B(_1868_),
    .Y(_1869_)
);

NAND2X1 _23491_ (
    .A(_1782_),
    .B(_1801_),
    .Y(_1871_)
);

NAND2X1 _23492_ (
    .A(_1869_),
    .B(_1871_),
    .Y(_1872_)
);

AOI21X1 _23493_ (
    .A(_1738_),
    .B(_1846_),
    .C(_1844_),
    .Y(_1873_)
);

INVX1 _23494_ (
    .A(_1822_),
    .Y(_1874_)
);

AOI21X1 _23495_ (
    .A(_1820_),
    .B(_1802_),
    .C(_1874_),
    .Y(_1875_)
);

NOR2X1 _23496_ (
    .A(_1798_),
    .B(_1792_),
    .Y(_1876_)
);

AND2X2 _23497_ (
    .A(_1799_),
    .B(_1788_),
    .Y(_1877_)
);

NOR2X1 _23498_ (
    .A(_1876_),
    .B(_1877_),
    .Y(_1878_)
);

NOR2X1 _23499_ (
    .A(_6300__bF$buf3),
    .B(_6815__bF$buf4),
    .Y(_1879_)
);

NAND2X1 _23500_ (
    .A(areg_27_bF$buf4),
    .B(breg_27_bF$buf5),
    .Y(_1880_)
);

NOR2X1 _23501_ (
    .A(_1679_),
    .B(_1880_),
    .Y(_1882_)
);

NOR2X1 _23502_ (
    .A(_1793_),
    .B(_1797_),
    .Y(_1883_)
);

NOR2X1 _23503_ (
    .A(_1882_),
    .B(_1883_),
    .Y(_1884_)
);

NAND2X1 _23504_ (
    .A(areg_26_bF$buf2),
    .B(breg_29_bF$buf1),
    .Y(_1885_)
);

NAND2X1 _23505_ (
    .A(areg_28_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_1886_)
);

OAI21X1 _23506_ (
    .A(_5668__bF$buf1),
    .B(_7520__bF$buf2),
    .C(_1795_),
    .Y(_1887_)
);

OAI21X1 _23507_ (
    .A(_1880_),
    .B(_1886_),
    .C(_1887_),
    .Y(_1888_)
);

XOR2X1 _23508_ (
    .A(_1888_),
    .B(_1885_),
    .Y(_1889_)
);

XNOR2X1 _23509_ (
    .A(_1884_),
    .B(_1889_),
    .Y(_1890_)
);

XOR2X1 _23510_ (
    .A(_1890_),
    .B(_1879_),
    .Y(_1891_)
);

XOR2X1 _23511_ (
    .A(_1878_),
    .B(_1891_),
    .Y(_1892_)
);

OAI21X1 _23512_ (
    .A(_5921__bF$buf3),
    .B(_7225__bF$buf4),
    .C(_1892_),
    .Y(_1893_)
);

NOR2X1 _23513_ (
    .A(_5921__bF$buf2),
    .B(_7225__bF$buf3),
    .Y(_1894_)
);

XNOR2X1 _23514_ (
    .A(_1878_),
    .B(_1891_),
    .Y(_1895_)
);

NAND2X1 _23515_ (
    .A(_1894_),
    .B(_1895_),
    .Y(_1896_)
);

NAND2X1 _23516_ (
    .A(_1806_),
    .B(_1818_),
    .Y(_1897_)
);

NAND2X1 _23517_ (
    .A(_1809_),
    .B(_1815_),
    .Y(_1898_)
);

NAND2X1 _23518_ (
    .A(_1808_),
    .B(_1817_),
    .Y(_1899_)
);

NAND2X1 _23519_ (
    .A(_1898_),
    .B(_1899_),
    .Y(_1900_)
);

OAI22X1 _23520_ (
    .A(_1703_),
    .B(_1811_),
    .C(_1814_),
    .D(_1810_),
    .Y(_1901_)
);

NAND2X1 _23521_ (
    .A(breg_26_bF$buf1),
    .B(areg_29_bF$buf1),
    .Y(_1903_)
);

NAND2X1 _23522_ (
    .A(breg_25_bF$buf2),
    .B(areg_31_bF$buf3),
    .Y(_1904_)
);

NOR2X1 _23523_ (
    .A(_1812_),
    .B(_1904_),
    .Y(_1905_)
);

INVX2 _23524_ (
    .A(_1811_),
    .Y(_1906_)
);

AOI21X1 _23525_ (
    .A(breg_24_bF$buf4),
    .B(areg_31_bF$buf2),
    .C(_1906_),
    .Y(_1907_)
);

NOR2X1 _23526_ (
    .A(_1905_),
    .B(_1907_),
    .Y(_1908_)
);

XNOR2X1 _23527_ (
    .A(_1908_),
    .B(_1903_),
    .Y(_1909_)
);

XNOR2X1 _23528_ (
    .A(_1909_),
    .B(_1901_),
    .Y(_1910_)
);

XNOR2X1 _23529_ (
    .A(_1900_),
    .B(_1910_),
    .Y(_1911_)
);

XNOR2X1 _23530_ (
    .A(_1911_),
    .B(_1897_),
    .Y(_1912_)
);

AOI21X1 _23531_ (
    .A(_1896_),
    .B(_1893_),
    .C(_1912_),
    .Y(_1915_)
);

NAND2X1 _23532_ (
    .A(_1896_),
    .B(_1893_),
    .Y(_1916_)
);

INVX2 _23533_ (
    .A(_1912_),
    .Y(_1917_)
);

NOR2X1 _23534_ (
    .A(_1917_),
    .B(_1916_),
    .Y(_1918_)
);

OAI21X1 _23535_ (
    .A(_1918_),
    .B(_1915_),
    .C(_1875_),
    .Y(_1919_)
);

OAI21X1 _23536_ (
    .A(_1826_),
    .B(_1825_),
    .C(_1822_),
    .Y(_1920_)
);

INVX1 _23537_ (
    .A(_1915_),
    .Y(_1921_)
);

OR2X2 _23538_ (
    .A(_1916_),
    .B(_1917_),
    .Y(_1922_)
);

NAND3X1 _23539_ (
    .A(_1921_),
    .B(_1920_),
    .C(_1922_),
    .Y(_1923_)
);

NAND2X1 _23540_ (
    .A(_1919_),
    .B(_1923_),
    .Y(_1924_)
);

NAND2X1 _23541_ (
    .A(_1924_),
    .B(_1834_),
    .Y(_1926_)
);

OR2X2 _23542_ (
    .A(_1834_),
    .B(_1924_),
    .Y(_1927_)
);

AOI21X1 _23543_ (
    .A(_1926_),
    .B(_1927_),
    .C(_1837_),
    .Y(_1928_)
);

NOR2X1 _23544_ (
    .A(_1829_),
    .B(_1924_),
    .Y(_1929_)
);

OAI21X1 _23545_ (
    .A(_1928_),
    .B(_1929_),
    .C(_1873_),
    .Y(_1930_)
);

OAI21X1 _23546_ (
    .A(_1841_),
    .B(_1727_),
    .C(_1847_),
    .Y(_1931_)
);

AND2X2 _23547_ (
    .A(_1834_),
    .B(_1924_),
    .Y(_1932_)
);

NOR2X1 _23548_ (
    .A(_1924_),
    .B(_1834_),
    .Y(_1933_)
);

OAI21X1 _23549_ (
    .A(_1932_),
    .B(_1933_),
    .C(_1829_),
    .Y(_1934_)
);

INVX1 _23550_ (
    .A(_1929_),
    .Y(_1935_)
);

NAND3X1 _23551_ (
    .A(_1934_),
    .B(_1935_),
    .C(_1931_),
    .Y(_1937_)
);

AOI21X1 _23552_ (
    .A(_1930_),
    .B(_1937_),
    .C(_1872_),
    .Y(_1938_)
);

INVX2 _23553_ (
    .A(_1872_),
    .Y(_1939_)
);

AOI21X1 _23554_ (
    .A(_1934_),
    .B(_1935_),
    .C(_1931_),
    .Y(_1940_)
);

NOR3X1 _23555_ (
    .A(_1928_),
    .B(_1929_),
    .C(_1873_),
    .Y(_1941_)
);

NOR3X1 _23556_ (
    .A(_1939_),
    .B(_1940_),
    .C(_1941_),
    .Y(_1942_)
);

OAI21X1 _23557_ (
    .A(_1942_),
    .B(_1938_),
    .C(_1867_),
    .Y(_1943_)
);

OAI21X1 _23558_ (
    .A(_1858_),
    .B(_1856_),
    .C(_1850_),
    .Y(_1944_)
);

OAI21X1 _23559_ (
    .A(_1941_),
    .B(_1940_),
    .C(_1939_),
    .Y(_1945_)
);

NAND3X1 _23560_ (
    .A(_1872_),
    .B(_1930_),
    .C(_1937_),
    .Y(_1946_)
);

NAND3X1 _23561_ (
    .A(_1946_),
    .B(_1944_),
    .C(_1945_),
    .Y(_1948_)
);

NAND2X1 _23562_ (
    .A(_1948_),
    .B(_1943_),
    .Y(_1949_)
);

INVX1 _23563_ (
    .A(_1949_),
    .Y(_1950_)
);

XNOR2X1 _23564_ (
    .A(_1866_),
    .B(_1950_),
    .Y(_0_[55])
);

INVX1 _23565_ (
    .A(_7644_),
    .Y(_1951_)
);

INVX1 _23566_ (
    .A(_6804_),
    .Y(_1952_)
);

NAND3X1 _23567_ (
    .A(_7633_),
    .B(_7637_),
    .C(_7213_),
    .Y(_1953_)
);

INVX1 _23568_ (
    .A(_7647_),
    .Y(_1954_)
);

OAI21X1 _23569_ (
    .A(_1952_),
    .B(_1953_),
    .C(_1954_),
    .Y(_1955_)
);

AOI21X1 _23570_ (
    .A(_6038_),
    .B(_1951_),
    .C(_1955_),
    .Y(_1956_)
);

AOI21X1 _23571_ (
    .A(_2746_),
    .B(_2747_),
    .C(_2745_),
    .Y(_1958_)
);

OAI21X1 _23572_ (
    .A(_2975_),
    .B(_2752_),
    .C(_1958_),
    .Y(_1959_)
);

NAND2X1 _23573_ (
    .A(_2969_),
    .B(_1959_),
    .Y(_1960_)
);

AOI21X1 _23574_ (
    .A(_3234_),
    .B(_3237_),
    .C(_3498_),
    .Y(_1961_)
);

AOI22X1 _23575_ (
    .A(_3497_),
    .B(_3511_),
    .C(_1961_),
    .D(_1960_),
    .Y(_1962_)
);

AOI21X1 _23576_ (
    .A(_3766_),
    .B(_3769_),
    .C(_4050_),
    .Y(_1963_)
);

AND2X2 _23577_ (
    .A(_4639_),
    .B(_4636_),
    .Y(_1964_)
);

NAND3X1 _23578_ (
    .A(_4343_),
    .B(_1964_),
    .C(_1963_),
    .Y(_1965_)
);

OAI21X1 _23579_ (
    .A(_1962_),
    .B(_1965_),
    .C(_4646_),
    .Y(_1966_)
);

NOR2X1 _23580_ (
    .A(_2750_),
    .B(_2974_),
    .Y(_1967_)
);

NAND2X1 _23581_ (
    .A(_1961_),
    .B(_1967_),
    .Y(_1969_)
);

NOR3X1 _23582_ (
    .A(_1969_),
    .B(_1965_),
    .C(_2545_),
    .Y(_1970_)
);

OAI21X1 _23583_ (
    .A(_1966_),
    .B(_1970_),
    .C(_7650_),
    .Y(_1971_)
);

AOI21X1 _23584_ (
    .A(_1956_),
    .B(_1971_),
    .C(_924_),
    .Y(_1972_)
);

INVX1 _23585_ (
    .A(_922_),
    .Y(_1973_)
);

NAND2X1 _23586_ (
    .A(_11877_),
    .B(_1973_),
    .Y(_1974_)
);

INVX1 _23587_ (
    .A(_920_),
    .Y(_1975_)
);

AND2X2 _23588_ (
    .A(_936_),
    .B(_725_),
    .Y(_1976_)
);

OAI21X1 _23589_ (
    .A(_917_),
    .B(_1976_),
    .C(_935_),
    .Y(_1977_)
);

OAI21X1 _23590_ (
    .A(_1975_),
    .B(_488_),
    .C(_1977_),
    .Y(_1978_)
);

AOI21X1 _23591_ (
    .A(_1973_),
    .B(_11873_),
    .C(_1978_),
    .Y(_1980_)
);

OAI21X1 _23592_ (
    .A(_10684_),
    .B(_1974_),
    .C(_1980_),
    .Y(_1981_)
);

AND2X2 _23593_ (
    .A(_1763_),
    .B(_1767_),
    .Y(_1982_)
);

AOI21X1 _23594_ (
    .A(_1862_),
    .B(_1863_),
    .C(_1949_),
    .Y(_1983_)
);

NAND3X1 _23595_ (
    .A(_1982_),
    .B(_1652_),
    .C(_1983_),
    .Y(_1984_)
);

NOR3X1 _23596_ (
    .A(_1258_),
    .B(_1540_),
    .C(_1984_),
    .Y(_1985_)
);

OAI21X1 _23597_ (
    .A(_1972_),
    .B(_1981_),
    .C(_1985_),
    .Y(_1986_)
);

INVX1 _23598_ (
    .A(_1984_),
    .Y(_1987_)
);

INVX1 _23599_ (
    .A(_1983_),
    .Y(_1988_)
);

NAND2X1 _23600_ (
    .A(_1943_),
    .B(_1865_),
    .Y(_1989_)
);

AND2X2 _23601_ (
    .A(_1989_),
    .B(_1948_),
    .Y(_1991_)
);

OAI21X1 _23602_ (
    .A(_1988_),
    .B(_1770_),
    .C(_1991_),
    .Y(_1992_)
);

AOI21X1 _23603_ (
    .A(_1987_),
    .B(_1545_),
    .C(_1992_),
    .Y(_1993_)
);

NAND2X1 _23604_ (
    .A(_1993_),
    .B(_1986_),
    .Y(_1994_)
);

OAI21X1 _23605_ (
    .A(_1940_),
    .B(_1939_),
    .C(_1937_),
    .Y(_1995_)
);

OAI21X1 _23606_ (
    .A(_1876_),
    .B(_1877_),
    .C(_1891_),
    .Y(_1996_)
);

NAND2X1 _23607_ (
    .A(_1996_),
    .B(_1896_),
    .Y(_1997_)
);

OAI21X1 _23608_ (
    .A(_1829_),
    .B(_1924_),
    .C(_1927_),
    .Y(_1998_)
);

NAND3X1 _23609_ (
    .A(_1806_),
    .B(_1818_),
    .C(_1911_),
    .Y(_1999_)
);

OAI21X1 _23610_ (
    .A(_1916_),
    .B(_1917_),
    .C(_1999_),
    .Y(_2000_)
);

NOR2X1 _23611_ (
    .A(_6300__bF$buf2),
    .B(_7225__bF$buf2),
    .Y(_2002_)
);

OAI21X1 _23612_ (
    .A(_1882_),
    .B(_1883_),
    .C(_1889_),
    .Y(_2003_)
);

INVX1 _23613_ (
    .A(_2003_),
    .Y(_2004_)
);

AND2X2 _23614_ (
    .A(_1890_),
    .B(_1879_),
    .Y(_2005_)
);

NOR2X1 _23615_ (
    .A(_2004_),
    .B(_2005_),
    .Y(_2006_)
);

NOR2X1 _23616_ (
    .A(_6686__bF$buf3),
    .B(_6815__bF$buf3),
    .Y(_2007_)
);

NOR2X1 _23617_ (
    .A(_1880_),
    .B(_1886_),
    .Y(_2008_)
);

NOR2X1 _23618_ (
    .A(_1885_),
    .B(_1888_),
    .Y(_2009_)
);

NOR2X1 _23619_ (
    .A(_2008_),
    .B(_2009_),
    .Y(_2010_)
);

NAND2X1 _23620_ (
    .A(areg_27_bF$buf3),
    .B(breg_29_bF$buf0),
    .Y(_2011_)
);

NAND2X1 _23621_ (
    .A(breg_27_bF$buf4),
    .B(areg_29_bF$buf0),
    .Y(_2013_)
);

NOR2X1 _23622_ (
    .A(_1886_),
    .B(_2013_),
    .Y(_2014_)
);

AND2X2 _23623_ (
    .A(_1886_),
    .B(_2013_),
    .Y(_2015_)
);

NOR2X1 _23624_ (
    .A(_2014_),
    .B(_2015_),
    .Y(_2016_)
);

XNOR2X1 _23625_ (
    .A(_2016_),
    .B(_2011_),
    .Y(_2017_)
);

XNOR2X1 _23626_ (
    .A(_2017_),
    .B(_2010_),
    .Y(_2018_)
);

NOR2X1 _23627_ (
    .A(_2007_),
    .B(_2018_),
    .Y(_2019_)
);

AND2X2 _23628_ (
    .A(_2018_),
    .B(_2007_),
    .Y(_2020_)
);

OAI21X1 _23629_ (
    .A(_2019_),
    .B(_2020_),
    .C(_2006_),
    .Y(_2021_)
);

NOR2X1 _23630_ (
    .A(_2019_),
    .B(_2020_),
    .Y(_2022_)
);

OAI21X1 _23631_ (
    .A(_2004_),
    .B(_2005_),
    .C(_2022_),
    .Y(_2024_)
);

AND2X2 _23632_ (
    .A(_2024_),
    .B(_2021_),
    .Y(_2025_)
);

XOR2X1 _23633_ (
    .A(_2025_),
    .B(_2002_),
    .Y(_2026_)
);

AOI21X1 _23634_ (
    .A(_1898_),
    .B(_1899_),
    .C(_1910_),
    .Y(_2027_)
);

NAND2X1 _23635_ (
    .A(_1901_),
    .B(_1909_),
    .Y(_2028_)
);

INVX1 _23636_ (
    .A(_1905_),
    .Y(_2029_)
);

OAI21X1 _23637_ (
    .A(_1907_),
    .B(_1903_),
    .C(_2029_),
    .Y(_2030_)
);

NOR2X1 _23638_ (
    .A(_5676_),
    .B(_8773_),
    .Y(_2031_)
);

AOI22X1 _23639_ (
    .A(breg_25_bF$buf1),
    .B(areg_31_bF$buf1),
    .C(breg_26_bF$buf0),
    .D(areg_30_bF$buf4),
    .Y(_2032_)
);

AOI21X1 _23640_ (
    .A(_1906_),
    .B(_2031_),
    .C(_2032_),
    .Y(_2033_)
);

NAND2X1 _23641_ (
    .A(_2033_),
    .B(_2030_),
    .Y(_2035_)
);

INVX1 _23642_ (
    .A(_2035_),
    .Y(_2036_)
);

NOR2X1 _23643_ (
    .A(_2033_),
    .B(_2030_),
    .Y(_2037_)
);

NOR2X1 _23644_ (
    .A(_2037_),
    .B(_2036_),
    .Y(_2038_)
);

XNOR2X1 _23645_ (
    .A(_2038_),
    .B(_2028_),
    .Y(_2039_)
);

OR2X2 _23646_ (
    .A(_2027_),
    .B(_2039_),
    .Y(_2040_)
);

NAND2X1 _23647_ (
    .A(_2039_),
    .B(_2027_),
    .Y(_2041_)
);

AND2X2 _23648_ (
    .A(_2040_),
    .B(_2041_),
    .Y(_2042_)
);

XNOR2X1 _23649_ (
    .A(_2026_),
    .B(_2042_),
    .Y(_2043_)
);

XNOR2X1 _23650_ (
    .A(_2043_),
    .B(_2000_),
    .Y(_2044_)
);

XNOR2X1 _23651_ (
    .A(_2044_),
    .B(_1923_),
    .Y(_2046_)
);

XOR2X1 _23652_ (
    .A(_2046_),
    .B(_1998_),
    .Y(_2047_)
);

XNOR2X1 _23653_ (
    .A(_2047_),
    .B(_1997_),
    .Y(_2048_)
);

XNOR2X1 _23654_ (
    .A(_2048_),
    .B(_1995_),
    .Y(_2049_)
);

AND2X2 _23655_ (
    .A(_1994_),
    .B(_2049_),
    .Y(_2050_)
);

NOR2X1 _23656_ (
    .A(_2049_),
    .B(_1994_),
    .Y(_2051_)
);

NOR2X1 _23657_ (
    .A(_2051_),
    .B(_2050_),
    .Y(_0_[56])
);

AOI21X1 _23658_ (
    .A(_1937_),
    .B(_1946_),
    .C(_2048_),
    .Y(_2052_)
);

NOR2X1 _23659_ (
    .A(_2052_),
    .B(_2050_),
    .Y(_2053_)
);

AND2X2 _23660_ (
    .A(_2046_),
    .B(_1998_),
    .Y(_2054_)
);

AOI21X1 _23661_ (
    .A(_1997_),
    .B(_2047_),
    .C(_2054_),
    .Y(_2056_)
);

NAND2X1 _23662_ (
    .A(_2002_),
    .B(_2025_),
    .Y(_2057_)
);

NAND2X1 _23663_ (
    .A(_2024_),
    .B(_2057_),
    .Y(_2058_)
);

INVX1 _23664_ (
    .A(_1923_),
    .Y(_2059_)
);

NAND2X1 _23665_ (
    .A(_2059_),
    .B(_2044_),
    .Y(_2060_)
);

AOI21X1 _23666_ (
    .A(_1999_),
    .B(_1922_),
    .C(_2043_),
    .Y(_2061_)
);

NAND2X1 _23667_ (
    .A(_2042_),
    .B(_2026_),
    .Y(_2062_)
);

NAND2X1 _23668_ (
    .A(_2041_),
    .B(_2062_),
    .Y(_2063_)
);

NOR2X1 _23669_ (
    .A(_6686__bF$buf2),
    .B(_7225__bF$buf1),
    .Y(_2064_)
);

INVX1 _23670_ (
    .A(_2010_),
    .Y(_2065_)
);

AOI21X1 _23671_ (
    .A(_2065_),
    .B(_2017_),
    .C(_2020_),
    .Y(_2067_)
);

NOR2X1 _23672_ (
    .A(_7100__bF$buf2),
    .B(_6815__bF$buf2),
    .Y(_2068_)
);

INVX1 _23673_ (
    .A(_2014_),
    .Y(_2069_)
);

OAI21X1 _23674_ (
    .A(_2015_),
    .B(_2011_),
    .C(_2069_),
    .Y(_2070_)
);

NAND2X1 _23675_ (
    .A(areg_28_bF$buf1),
    .B(breg_29_bF$buf4),
    .Y(_2071_)
);

NAND2X1 _23676_ (
    .A(breg_28_bF$buf3),
    .B(areg_30_bF$buf3),
    .Y(_2072_)
);

NOR2X1 _23677_ (
    .A(_2013_),
    .B(_2072_),
    .Y(_2073_)
);

AOI22X1 _23678_ (
    .A(breg_27_bF$buf3),
    .B(areg_30_bF$buf2),
    .C(breg_28_bF$buf2),
    .D(areg_29_bF$buf5),
    .Y(_2074_)
);

OAI21X1 _23679_ (
    .A(_2073_),
    .B(_2074_),
    .C(_2071_),
    .Y(_2075_)
);

NOR2X1 _23680_ (
    .A(_2074_),
    .B(_2073_),
    .Y(_2076_)
);

NAND3X1 _23681_ (
    .A(areg_28_bF$buf0),
    .B(breg_29_bF$buf3),
    .C(_2076_),
    .Y(_2078_)
);

NAND2X1 _23682_ (
    .A(_2075_),
    .B(_2078_),
    .Y(_2079_)
);

XNOR2X1 _23683_ (
    .A(_2079_),
    .B(_2070_),
    .Y(_2080_)
);

XOR2X1 _23684_ (
    .A(_2080_),
    .B(_2068_),
    .Y(_2081_)
);

XNOR2X1 _23685_ (
    .A(_2067_),
    .B(_2081_),
    .Y(_2082_)
);

XNOR2X1 _23686_ (
    .A(_2082_),
    .B(_2064_),
    .Y(_2083_)
);

INVX1 _23687_ (
    .A(_2038_),
    .Y(_2084_)
);

NOR2X1 _23688_ (
    .A(_2028_),
    .B(_2084_),
    .Y(_2085_)
);

INVX1 _23689_ (
    .A(_2031_),
    .Y(_2086_)
);

OAI21X1 _23690_ (
    .A(_1906_),
    .B(_2086_),
    .C(_2035_),
    .Y(_2087_)
);

NAND3X1 _23691_ (
    .A(_1811_),
    .B(_2031_),
    .C(_2036_),
    .Y(_2089_)
);

AND2X2 _23692_ (
    .A(_2089_),
    .B(_2087_),
    .Y(_2090_)
);

XOR2X1 _23693_ (
    .A(_2085_),
    .B(_2090_),
    .Y(_2091_)
);

INVX1 _23694_ (
    .A(_2091_),
    .Y(_2092_)
);

OR2X2 _23695_ (
    .A(_2083_),
    .B(_2092_),
    .Y(_2093_)
);

NAND2X1 _23696_ (
    .A(_2092_),
    .B(_2083_),
    .Y(_2094_)
);

NAND2X1 _23697_ (
    .A(_2094_),
    .B(_2093_),
    .Y(_2095_)
);

XNOR2X1 _23698_ (
    .A(_2095_),
    .B(_2063_),
    .Y(_2096_)
);

XNOR2X1 _23699_ (
    .A(_2096_),
    .B(_2061_),
    .Y(_2097_)
);

NAND2X1 _23700_ (
    .A(_2060_),
    .B(_2097_),
    .Y(_2098_)
);

OR2X2 _23701_ (
    .A(_2097_),
    .B(_2060_),
    .Y(_2100_)
);

NAND2X1 _23702_ (
    .A(_2098_),
    .B(_2100_),
    .Y(_2101_)
);

XOR2X1 _23703_ (
    .A(_2101_),
    .B(_2058_),
    .Y(_2102_)
);

NAND2X1 _23704_ (
    .A(_2056_),
    .B(_2102_),
    .Y(_2103_)
);

OR2X2 _23705_ (
    .A(_2102_),
    .B(_2056_),
    .Y(_2104_)
);

AND2X2 _23706_ (
    .A(_2104_),
    .B(_2103_),
    .Y(_2105_)
);

XNOR2X1 _23707_ (
    .A(_2053_),
    .B(_2105_),
    .Y(_0_[57])
);

AOI21X1 _23708_ (
    .A(_1534_),
    .B(_1535_),
    .C(_1532_),
    .Y(_2106_)
);

NOR3X1 _23709_ (
    .A(_1542_),
    .B(_2106_),
    .C(_1400_),
    .Y(_2107_)
);

OAI21X1 _23710_ (
    .A(_2106_),
    .B(_1398_),
    .C(_1536_),
    .Y(_2108_)
);

AOI21X1 _23711_ (
    .A(_1257_),
    .B(_2107_),
    .C(_2108_),
    .Y(_2110_)
);

OAI21X1 _23712_ (
    .A(_1768_),
    .B(_1654_),
    .C(_1767_),
    .Y(_2111_)
);

NAND2X1 _23713_ (
    .A(_1948_),
    .B(_1989_),
    .Y(_2112_)
);

AOI21X1 _23714_ (
    .A(_1983_),
    .B(_2111_),
    .C(_2112_),
    .Y(_2113_)
);

OAI21X1 _23715_ (
    .A(_2110_),
    .B(_1984_),
    .C(_2113_),
    .Y(_2114_)
);

AOI21X1 _23716_ (
    .A(_1985_),
    .B(_942_),
    .C(_2114_),
    .Y(_2115_)
);

NOR2X1 _23717_ (
    .A(_2056_),
    .B(_2102_),
    .Y(_2116_)
);

AOI21X1 _23718_ (
    .A(_2052_),
    .B(_2103_),
    .C(_2116_),
    .Y(_2117_)
);

NAND2X1 _23719_ (
    .A(_2049_),
    .B(_2105_),
    .Y(_2118_)
);

OAI21X1 _23720_ (
    .A(_2115_),
    .B(_2118_),
    .C(_2117_),
    .Y(_2119_)
);

INVX1 _23721_ (
    .A(_2100_),
    .Y(_2121_)
);

AOI21X1 _23722_ (
    .A(_2058_),
    .B(_2098_),
    .C(_2121_),
    .Y(_2122_)
);

INVX1 _23723_ (
    .A(_2081_),
    .Y(_2123_)
);

NOR2X1 _23724_ (
    .A(_2067_),
    .B(_2123_),
    .Y(_2124_)
);

AOI21X1 _23725_ (
    .A(_2064_),
    .B(_2082_),
    .C(_2124_),
    .Y(_2125_)
);

NAND2X1 _23726_ (
    .A(_2061_),
    .B(_2096_),
    .Y(_2126_)
);

AOI21X1 _23727_ (
    .A(_2041_),
    .B(_2062_),
    .C(_2095_),
    .Y(_2127_)
);

NOR2X1 _23728_ (
    .A(_2092_),
    .B(_2083_),
    .Y(_2128_)
);

AOI21X1 _23729_ (
    .A(_2085_),
    .B(_2090_),
    .C(_2128_),
    .Y(_2129_)
);

NOR2X1 _23730_ (
    .A(_7100__bF$buf1),
    .B(_7225__bF$buf0),
    .Y(_2130_)
);

NAND3X1 _23731_ (
    .A(_2070_),
    .B(_2075_),
    .C(_2078_),
    .Y(_2132_)
);

NAND2X1 _23732_ (
    .A(_2068_),
    .B(_2080_),
    .Y(_2133_)
);

NAND2X1 _23733_ (
    .A(_2132_),
    .B(_2133_),
    .Y(_2134_)
);

NOR2X1 _23734_ (
    .A(_7520__bF$buf1),
    .B(_6815__bF$buf1),
    .Y(_2135_)
);

OAI21X1 _23735_ (
    .A(_2013_),
    .B(_2072_),
    .C(_2078_),
    .Y(_2136_)
);

NAND2X1 _23736_ (
    .A(areg_29_bF$buf4),
    .B(breg_29_bF$buf2),
    .Y(_2137_)
);

NAND2X1 _23737_ (
    .A(breg_27_bF$buf2),
    .B(areg_30_bF$buf1),
    .Y(_2138_)
);

NAND2X1 _23738_ (
    .A(breg_28_bF$buf1),
    .B(areg_31_bF$buf0),
    .Y(_2139_)
);

OAI21X1 _23739_ (
    .A(_5668__bF$buf0),
    .B(_8773_),
    .C(_2072_),
    .Y(_2140_)
);

OAI21X1 _23740_ (
    .A(_2138_),
    .B(_2139_),
    .C(_2140_),
    .Y(_2141_)
);

XNOR2X1 _23741_ (
    .A(_2141_),
    .B(_2137_),
    .Y(_2143_)
);

XNOR2X1 _23742_ (
    .A(_2136_),
    .B(_2143_),
    .Y(_2144_)
);

XNOR2X1 _23743_ (
    .A(_2144_),
    .B(_2135_),
    .Y(_2145_)
);

XNOR2X1 _23744_ (
    .A(_2145_),
    .B(_2134_),
    .Y(_2146_)
);

XOR2X1 _23745_ (
    .A(_2146_),
    .B(_2130_),
    .Y(_2147_)
);

OAI21X1 _23746_ (
    .A(_1811_),
    .B(_2086_),
    .C(_2089_),
    .Y(_2148_)
);

XNOR2X1 _23747_ (
    .A(_2147_),
    .B(_2148_),
    .Y(_2149_)
);

XOR2X1 _23748_ (
    .A(_2129_),
    .B(_2149_),
    .Y(_2150_)
);

XNOR2X1 _23749_ (
    .A(_2150_),
    .B(_2127_),
    .Y(_2151_)
);

XNOR2X1 _23750_ (
    .A(_2151_),
    .B(_2126_),
    .Y(_2152_)
);

XNOR2X1 _23751_ (
    .A(_2152_),
    .B(_2125_),
    .Y(_2154_)
);

NOR2X1 _23752_ (
    .A(_2122_),
    .B(_2154_),
    .Y(_2155_)
);

INVX1 _23753_ (
    .A(_2155_),
    .Y(_2156_)
);

NAND2X1 _23754_ (
    .A(_2122_),
    .B(_2154_),
    .Y(_2157_)
);

NAND2X1 _23755_ (
    .A(_2157_),
    .B(_2156_),
    .Y(_2158_)
);

INVX2 _23756_ (
    .A(_2158_),
    .Y(_2159_)
);

AND2X2 _23757_ (
    .A(_2119_),
    .B(_2159_),
    .Y(_2160_)
);

NOR2X1 _23758_ (
    .A(_2159_),
    .B(_2119_),
    .Y(_2161_)
);

NOR2X1 _23759_ (
    .A(_2161_),
    .B(_2160_),
    .Y(_0_[58])
);

NOR2X1 _23760_ (
    .A(_2126_),
    .B(_2151_),
    .Y(_2162_)
);

NOR2X1 _23761_ (
    .A(_2125_),
    .B(_2152_),
    .Y(_2164_)
);

NOR2X1 _23762_ (
    .A(_2162_),
    .B(_2164_),
    .Y(_2165_)
);

INVX1 _23763_ (
    .A(_2134_),
    .Y(_2166_)
);

NAND2X1 _23764_ (
    .A(_2130_),
    .B(_2146_),
    .Y(_2167_)
);

OAI21X1 _23765_ (
    .A(_2166_),
    .B(_2145_),
    .C(_2167_),
    .Y(_2168_)
);

NAND2X1 _23766_ (
    .A(_2127_),
    .B(_2150_),
    .Y(_2169_)
);

NAND2X1 _23767_ (
    .A(_2148_),
    .B(_2147_),
    .Y(_2170_)
);

NOR2X1 _23768_ (
    .A(_7520__bF$buf0),
    .B(_7225__bF$buf4),
    .Y(_2171_)
);

INVX1 _23769_ (
    .A(_2143_),
    .Y(_2172_)
);

NAND2X1 _23770_ (
    .A(_2136_),
    .B(_2172_),
    .Y(_2173_)
);

NAND2X1 _23771_ (
    .A(_2135_),
    .B(_2144_),
    .Y(_2175_)
);

NAND2X1 _23772_ (
    .A(_2173_),
    .B(_2175_),
    .Y(_2176_)
);

NOR2X1 _23773_ (
    .A(_9153_),
    .B(_6815__bF$buf0),
    .Y(_2177_)
);

OAI22X1 _23774_ (
    .A(_2138_),
    .B(_2139_),
    .C(_2141_),
    .D(_2137_),
    .Y(_2178_)
);

NAND2X1 _23775_ (
    .A(breg_29_bF$buf1),
    .B(areg_30_bF$buf0),
    .Y(_2179_)
);

XOR2X1 _23776_ (
    .A(_2139_),
    .B(_2179_),
    .Y(_2180_)
);

XOR2X1 _23777_ (
    .A(_2178_),
    .B(_2180_),
    .Y(_2181_)
);

XNOR2X1 _23778_ (
    .A(_2181_),
    .B(_2177_),
    .Y(_2182_)
);

XNOR2X1 _23779_ (
    .A(_2176_),
    .B(_2182_),
    .Y(_2183_)
);

XNOR2X1 _23780_ (
    .A(_2183_),
    .B(_2171_),
    .Y(_2184_)
);

NOR2X1 _23781_ (
    .A(_2184_),
    .B(_2170_),
    .Y(_2186_)
);

INVX1 _23782_ (
    .A(_2186_),
    .Y(_2187_)
);

NAND2X1 _23783_ (
    .A(_2184_),
    .B(_2170_),
    .Y(_2188_)
);

NAND2X1 _23784_ (
    .A(_2188_),
    .B(_2187_),
    .Y(_2189_)
);

OAI21X1 _23785_ (
    .A(_2129_),
    .B(_2149_),
    .C(_2189_),
    .Y(_2190_)
);

OR2X2 _23786_ (
    .A(_2129_),
    .B(_2149_),
    .Y(_2191_)
);

OR2X2 _23787_ (
    .A(_2191_),
    .B(_2189_),
    .Y(_2192_)
);

NAND2X1 _23788_ (
    .A(_2190_),
    .B(_2192_),
    .Y(_2193_)
);

NAND2X1 _23789_ (
    .A(_2169_),
    .B(_2193_),
    .Y(_2194_)
);

OR2X2 _23790_ (
    .A(_2193_),
    .B(_2169_),
    .Y(_2195_)
);

NAND2X1 _23791_ (
    .A(_2194_),
    .B(_2195_),
    .Y(_2197_)
);

XOR2X1 _23792_ (
    .A(_2197_),
    .B(_2168_),
    .Y(_2198_)
);

NOR2X1 _23793_ (
    .A(_2198_),
    .B(_2165_),
    .Y(_2199_)
);

INVX1 _23794_ (
    .A(_2199_),
    .Y(_2200_)
);

NAND2X1 _23795_ (
    .A(_2198_),
    .B(_2165_),
    .Y(_2201_)
);

AND2X2 _23796_ (
    .A(_2200_),
    .B(_2201_),
    .Y(_2202_)
);

INVX1 _23797_ (
    .A(_2202_),
    .Y(_2203_)
);

OAI21X1 _23798_ (
    .A(_2160_),
    .B(_2155_),
    .C(_2203_),
    .Y(_2204_)
);

NAND2X1 _23799_ (
    .A(_2159_),
    .B(_2119_),
    .Y(_2205_)
);

NAND3X1 _23800_ (
    .A(_2156_),
    .B(_2202_),
    .C(_2205_),
    .Y(_2206_)
);

NAND2X1 _23801_ (
    .A(_2206_),
    .B(_2204_),
    .Y(_0_[59])
);

NAND2X1 _23802_ (
    .A(_2202_),
    .B(_2159_),
    .Y(_2208_)
);

OR2X2 _23803_ (
    .A(_2208_),
    .B(_2118_),
    .Y(_2209_)
);

OAI21X1 _23804_ (
    .A(_2199_),
    .B(_2155_),
    .C(_2201_),
    .Y(_2210_)
);

OAI21X1 _23805_ (
    .A(_2208_),
    .B(_2117_),
    .C(_2210_),
    .Y(_2211_)
);

INVX1 _23806_ (
    .A(_2211_),
    .Y(_2212_)
);

OAI21X1 _23807_ (
    .A(_2115_),
    .B(_2209_),
    .C(_2212_),
    .Y(_2213_)
);

NAND3X1 _23808_ (
    .A(_2168_),
    .B(_2194_),
    .C(_2195_),
    .Y(_2214_)
);

OAI21X1 _23809_ (
    .A(_2169_),
    .B(_2193_),
    .C(_2214_),
    .Y(_2215_)
);

INVX1 _23810_ (
    .A(_2176_),
    .Y(_2216_)
);

NAND2X1 _23811_ (
    .A(_2171_),
    .B(_2183_),
    .Y(_2218_)
);

OAI21X1 _23812_ (
    .A(_2216_),
    .B(_2182_),
    .C(_2218_),
    .Y(_2219_)
);

NAND2X1 _23813_ (
    .A(_2180_),
    .B(_2178_),
    .Y(_2220_)
);

NAND2X1 _23814_ (
    .A(_2177_),
    .B(_2181_),
    .Y(_2221_)
);

NAND2X1 _23815_ (
    .A(_2220_),
    .B(_2221_),
    .Y(_2222_)
);

NOR2X1 _23816_ (
    .A(_8759_),
    .B(_6815__bF$buf4),
    .Y(_2223_)
);

NAND3X1 _23817_ (
    .A(breg_29_bF$buf0),
    .B(areg_31_bF$buf4),
    .C(_2072_),
    .Y(_2224_)
);

XNOR2X1 _23818_ (
    .A(_2224_),
    .B(_2223_),
    .Y(_2225_)
);

XOR2X1 _23819_ (
    .A(_2222_),
    .B(_2225_),
    .Y(_2226_)
);

INVX1 _23820_ (
    .A(_2226_),
    .Y(_2227_)
);

OAI21X1 _23821_ (
    .A(_9153_),
    .B(_7225__bF$buf3),
    .C(_2227_),
    .Y(_2229_)
);

NAND3X1 _23822_ (
    .A(areg_29_bF$buf3),
    .B(breg[31]),
    .C(_2226_),
    .Y(_2230_)
);

AND2X2 _23823_ (
    .A(_2229_),
    .B(_2230_),
    .Y(_2231_)
);

OAI21X1 _23824_ (
    .A(_2191_),
    .B(_2189_),
    .C(_2187_),
    .Y(_2232_)
);

XOR2X1 _23825_ (
    .A(_2232_),
    .B(_2231_),
    .Y(_2233_)
);

XOR2X1 _23826_ (
    .A(_2233_),
    .B(_2219_),
    .Y(_2234_)
);

XNOR2X1 _23827_ (
    .A(_2215_),
    .B(_2234_),
    .Y(_2235_)
);

XNOR2X1 _23828_ (
    .A(_2213_),
    .B(_2235_),
    .Y(_0_[60])
);

AOI21X1 _23829_ (
    .A(_1993_),
    .B(_1986_),
    .C(_2209_),
    .Y(_2236_)
);

NOR2X1 _23830_ (
    .A(_2211_),
    .B(_2236_),
    .Y(_2237_)
);

NAND2X1 _23831_ (
    .A(_2234_),
    .B(_2215_),
    .Y(_2239_)
);

OAI21X1 _23832_ (
    .A(_2237_),
    .B(_2235_),
    .C(_2239_),
    .Y(_2240_)
);

INVX1 _23833_ (
    .A(_2192_),
    .Y(_2241_)
);

AOI22X1 _23834_ (
    .A(_2241_),
    .B(_2231_),
    .C(_2233_),
    .D(_2219_),
    .Y(_2242_)
);

NAND2X1 _23835_ (
    .A(_2225_),
    .B(_2222_),
    .Y(_2243_)
);

NAND2X1 _23836_ (
    .A(_2243_),
    .B(_2230_),
    .Y(_2244_)
);

AND2X2 _23837_ (
    .A(_2186_),
    .B(_2231_),
    .Y(_2245_)
);

NAND2X1 _23838_ (
    .A(areg_30_bF$buf5),
    .B(breg[31]),
    .Y(_2246_)
);

INVX1 _23839_ (
    .A(_2223_),
    .Y(_2247_)
);

OAI22X1 _23840_ (
    .A(_2139_),
    .B(_2179_),
    .C(_2247_),
    .D(_2224_),
    .Y(_2248_)
);

NOR2X1 _23841_ (
    .A(_6815__bF$buf3),
    .B(_8773_),
    .Y(_2250_)
);

XOR2X1 _23842_ (
    .A(_2248_),
    .B(_2250_),
    .Y(_2251_)
);

XNOR2X1 _23843_ (
    .A(_2251_),
    .B(_2246_),
    .Y(_2252_)
);

XOR2X1 _23844_ (
    .A(_2245_),
    .B(_2252_),
    .Y(_2253_)
);

XNOR2X1 _23845_ (
    .A(_2253_),
    .B(_2244_),
    .Y(_2254_)
);

XOR2X1 _23846_ (
    .A(_2242_),
    .B(_2254_),
    .Y(_2255_)
);

INVX2 _23847_ (
    .A(_2255_),
    .Y(_2256_)
);

XNOR2X1 _23848_ (
    .A(_2240_),
    .B(_2256_),
    .Y(_0_[61])
);

NOR2X1 _23849_ (
    .A(_2256_),
    .B(_2235_),
    .Y(_2257_)
);

NOR2X1 _23850_ (
    .A(_2254_),
    .B(_2242_),
    .Y(_2258_)
);

INVX1 _23851_ (
    .A(_2258_),
    .Y(_2260_)
);

OAI21X1 _23852_ (
    .A(_2256_),
    .B(_2239_),
    .C(_2260_),
    .Y(_2261_)
);

AOI21X1 _23853_ (
    .A(_2257_),
    .B(_2213_),
    .C(_2261_),
    .Y(_2262_)
);

NAND2X1 _23854_ (
    .A(_2252_),
    .B(_2245_),
    .Y(_2263_)
);

NAND2X1 _23855_ (
    .A(_2244_),
    .B(_2253_),
    .Y(_2264_)
);

NAND2X1 _23856_ (
    .A(_2263_),
    .B(_2264_),
    .Y(_2265_)
);

NAND2X1 _23857_ (
    .A(_2250_),
    .B(_2248_),
    .Y(_2266_)
);

NOR2X1 _23858_ (
    .A(_2250_),
    .B(_2248_),
    .Y(_2267_)
);

OAI21X1 _23859_ (
    .A(_2267_),
    .B(_2246_),
    .C(_2266_),
    .Y(_2268_)
);

NOR2X1 _23860_ (
    .A(_8773_),
    .B(_7225__bF$buf2),
    .Y(_2269_)
);

NAND2X1 _23861_ (
    .A(_2269_),
    .B(_2268_),
    .Y(_2271_)
);

INVX1 _23862_ (
    .A(_2271_),
    .Y(_2272_)
);

NOR2X1 _23863_ (
    .A(_2269_),
    .B(_2268_),
    .Y(_2273_)
);

NOR2X1 _23864_ (
    .A(_2273_),
    .B(_2272_),
    .Y(_2274_)
);

NOR2X1 _23865_ (
    .A(_2274_),
    .B(_2265_),
    .Y(_2275_)
);

AND2X2 _23866_ (
    .A(_2265_),
    .B(_2274_),
    .Y(_2276_)
);

NOR2X1 _23867_ (
    .A(_2275_),
    .B(_2276_),
    .Y(_2277_)
);

XNOR2X1 _23868_ (
    .A(_2262_),
    .B(_2277_),
    .Y(_0_[62])
);

OAI21X1 _23869_ (
    .A(_2236_),
    .B(_2211_),
    .C(_2257_),
    .Y(_2278_)
);

INVX1 _23870_ (
    .A(_2261_),
    .Y(_2279_)
);

INVX1 _23871_ (
    .A(_2277_),
    .Y(_2281_)
);

AOI21X1 _23872_ (
    .A(_2279_),
    .B(_2278_),
    .C(_2281_),
    .Y(_2282_)
);

OAI21X1 _23873_ (
    .A(_2282_),
    .B(_2276_),
    .C(_2271_),
    .Y(_2283_)
);

INVX1 _23874_ (
    .A(_2265_),
    .Y(_2284_)
);

OAI21X1 _23875_ (
    .A(_2262_),
    .B(_2284_),
    .C(_2272_),
    .Y(_2285_)
);

NAND2X1 _23876_ (
    .A(_2285_),
    .B(_2283_),
    .Y(_0_[63])
);

XNOR2X1 _23877_ (
    .A(_3231_),
    .B(_3055_),
    .Y(_0_[1])
);

NOR2X1 _23878_ (
    .A(_2551__bF$buf1),
    .B(_2376__bF$buf0),
    .Y(_0_[0])
);

XOR2X1 _23879_ (
    .A(_3263_),
    .B(_3252_),
    .Y(_0_[2])
);

XOR2X1 _23880_ (
    .A(_3285_),
    .B(_3274_),
    .Y(_0_[3])
);

XOR2X1 _23881_ (
    .A(_3307_),
    .B(_3296_),
    .Y(_0_[4])
);

BUFX2 _23882_ (
    .A(_11909_[0]),
    .Y(y[0])
);

BUFX2 _23883_ (
    .A(_11909_[1]),
    .Y(y[1])
);

BUFX2 _23884_ (
    .A(_11909_[2]),
    .Y(y[2])
);

BUFX2 _23885_ (
    .A(_11909_[3]),
    .Y(y[3])
);

BUFX2 _23886_ (
    .A(_11909_[4]),
    .Y(y[4])
);

BUFX2 _23887_ (
    .A(_11909_[5]),
    .Y(y[5])
);

BUFX2 _23888_ (
    .A(_11909_[6]),
    .Y(y[6])
);

BUFX2 _23889_ (
    .A(_11909_[7]),
    .Y(y[7])
);

BUFX2 _23890_ (
    .A(_11909_[8]),
    .Y(y[8])
);

BUFX2 _23891_ (
    .A(_11909_[9]),
    .Y(y[9])
);

BUFX2 _23892_ (
    .A(_11909_[10]),
    .Y(y[10])
);

BUFX2 _23893_ (
    .A(_11909_[11]),
    .Y(y[11])
);

BUFX2 _23894_ (
    .A(_11909_[12]),
    .Y(y[12])
);

BUFX2 _23895_ (
    .A(_11909_[13]),
    .Y(y[13])
);

BUFX2 _23896_ (
    .A(_11909_[14]),
    .Y(y[14])
);

BUFX2 _23897_ (
    .A(_11909_[15]),
    .Y(y[15])
);

BUFX2 _23898_ (
    .A(_11909_[16]),
    .Y(y[16])
);

BUFX2 _23899_ (
    .A(_11909_[17]),
    .Y(y[17])
);

BUFX2 _23900_ (
    .A(_11909_[18]),
    .Y(y[18])
);

BUFX2 _23901_ (
    .A(_11909_[19]),
    .Y(y[19])
);

BUFX2 _23902_ (
    .A(_11909_[20]),
    .Y(y[20])
);

BUFX2 _23903_ (
    .A(_11909_[21]),
    .Y(y[21])
);

BUFX2 _23904_ (
    .A(_11909_[22]),
    .Y(y[22])
);

BUFX2 _23905_ (
    .A(_11909_[23]),
    .Y(y[23])
);

BUFX2 _23906_ (
    .A(_11909_[24]),
    .Y(y[24])
);

BUFX2 _23907_ (
    .A(_11909_[25]),
    .Y(y[25])
);

BUFX2 _23908_ (
    .A(_11909_[26]),
    .Y(y[26])
);

BUFX2 _23909_ (
    .A(_11909_[27]),
    .Y(y[27])
);

BUFX2 _23910_ (
    .A(_11909_[28]),
    .Y(y[28])
);

BUFX2 _23911_ (
    .A(_11909_[29]),
    .Y(y[29])
);

BUFX2 _23912_ (
    .A(_11909_[30]),
    .Y(y[30])
);

BUFX2 _23913_ (
    .A(_11909_[31]),
    .Y(y[31])
);

BUFX2 _23914_ (
    .A(_11909_[32]),
    .Y(y[32])
);

BUFX2 _23915_ (
    .A(_11909_[33]),
    .Y(y[33])
);

BUFX2 _23916_ (
    .A(_11909_[34]),
    .Y(y[34])
);

BUFX2 _23917_ (
    .A(_11909_[35]),
    .Y(y[35])
);

BUFX2 _23918_ (
    .A(_11909_[36]),
    .Y(y[36])
);

BUFX2 _23919_ (
    .A(_11909_[37]),
    .Y(y[37])
);

BUFX2 _23920_ (
    .A(_11909_[38]),
    .Y(y[38])
);

BUFX2 _23921_ (
    .A(_11909_[39]),
    .Y(y[39])
);

BUFX2 _23922_ (
    .A(_11909_[40]),
    .Y(y[40])
);

BUFX2 _23923_ (
    .A(_11909_[41]),
    .Y(y[41])
);

BUFX2 _23924_ (
    .A(_11909_[42]),
    .Y(y[42])
);

BUFX2 _23925_ (
    .A(_11909_[43]),
    .Y(y[43])
);

BUFX2 _23926_ (
    .A(_11909_[44]),
    .Y(y[44])
);

BUFX2 _23927_ (
    .A(_11909_[45]),
    .Y(y[45])
);

BUFX2 _23928_ (
    .A(_11909_[46]),
    .Y(y[46])
);

BUFX2 _23929_ (
    .A(_11909_[47]),
    .Y(y[47])
);

BUFX2 _23930_ (
    .A(_11909_[48]),
    .Y(y[48])
);

BUFX2 _23931_ (
    .A(_11909_[49]),
    .Y(y[49])
);

BUFX2 _23932_ (
    .A(_11909_[50]),
    .Y(y[50])
);

BUFX2 _23933_ (
    .A(_11909_[51]),
    .Y(y[51])
);

BUFX2 _23934_ (
    .A(_11909_[52]),
    .Y(y[52])
);

BUFX2 _23935_ (
    .A(_11909_[53]),
    .Y(y[53])
);

BUFX2 _23936_ (
    .A(_11909_[54]),
    .Y(y[54])
);

BUFX2 _23937_ (
    .A(_11909_[55]),
    .Y(y[55])
);

BUFX2 _23938_ (
    .A(_11909_[56]),
    .Y(y[56])
);

BUFX2 _23939_ (
    .A(_11909_[57]),
    .Y(y[57])
);

BUFX2 _23940_ (
    .A(_11909_[58]),
    .Y(y[58])
);

BUFX2 _23941_ (
    .A(_11909_[59]),
    .Y(y[59])
);

BUFX2 _23942_ (
    .A(_11909_[60]),
    .Y(y[60])
);

BUFX2 _23943_ (
    .A(_11909_[61]),
    .Y(y[61])
);

BUFX2 _23944_ (
    .A(_11909_[62]),
    .Y(y[62])
);

BUFX2 _23945_ (
    .A(_11909_[63]),
    .Y(y[63])
);

DFFPOSX1 _23946_ (
    .CLK(clk_bF$buf10),
    .D(_0_[0]),
    .Q(_11909_[0])
);

DFFPOSX1 _23947_ (
    .CLK(clk_bF$buf9),
    .D(_0_[1]),
    .Q(_11909_[1])
);

DFFPOSX1 _23948_ (
    .CLK(clk_bF$buf8),
    .D(_0_[2]),
    .Q(_11909_[2])
);

DFFPOSX1 _23949_ (
    .CLK(clk_bF$buf7),
    .D(_0_[3]),
    .Q(_11909_[3])
);

DFFPOSX1 _23950_ (
    .CLK(clk_bF$buf6),
    .D(_0_[4]),
    .Q(_11909_[4])
);

DFFPOSX1 _23951_ (
    .CLK(clk_bF$buf5),
    .D(_0_[5]),
    .Q(_11909_[5])
);

DFFPOSX1 _23952_ (
    .CLK(clk_bF$buf4),
    .D(_0_[6]),
    .Q(_11909_[6])
);

DFFPOSX1 _23953_ (
    .CLK(clk_bF$buf3),
    .D(_0_[7]),
    .Q(_11909_[7])
);

DFFPOSX1 _23954_ (
    .CLK(clk_bF$buf2),
    .D(_0_[8]),
    .Q(_11909_[8])
);

DFFPOSX1 _23955_ (
    .CLK(clk_bF$buf1),
    .D(_0_[9]),
    .Q(_11909_[9])
);

DFFPOSX1 _23956_ (
    .CLK(clk_bF$buf0),
    .D(_0_[10]),
    .Q(_11909_[10])
);

DFFPOSX1 _23957_ (
    .CLK(clk_bF$buf10),
    .D(_0_[11]),
    .Q(_11909_[11])
);

DFFPOSX1 _23958_ (
    .CLK(clk_bF$buf9),
    .D(_0_[12]),
    .Q(_11909_[12])
);

DFFPOSX1 _23959_ (
    .CLK(clk_bF$buf8),
    .D(_0_[13]),
    .Q(_11909_[13])
);

DFFPOSX1 _23960_ (
    .CLK(clk_bF$buf7),
    .D(_0_[14]),
    .Q(_11909_[14])
);

DFFPOSX1 _23961_ (
    .CLK(clk_bF$buf6),
    .D(_0_[15]),
    .Q(_11909_[15])
);

DFFPOSX1 _23962_ (
    .CLK(clk_bF$buf5),
    .D(_0_[16]),
    .Q(_11909_[16])
);

DFFPOSX1 _23963_ (
    .CLK(clk_bF$buf4),
    .D(_0_[17]),
    .Q(_11909_[17])
);

DFFPOSX1 _23964_ (
    .CLK(clk_bF$buf3),
    .D(_0_[18]),
    .Q(_11909_[18])
);

DFFPOSX1 _23965_ (
    .CLK(clk_bF$buf2),
    .D(_0_[19]),
    .Q(_11909_[19])
);

DFFPOSX1 _23966_ (
    .CLK(clk_bF$buf1),
    .D(_0_[20]),
    .Q(_11909_[20])
);

DFFPOSX1 _23967_ (
    .CLK(clk_bF$buf0),
    .D(_0_[21]),
    .Q(_11909_[21])
);

DFFPOSX1 _23968_ (
    .CLK(clk_bF$buf10),
    .D(_0_[22]),
    .Q(_11909_[22])
);

DFFPOSX1 _23969_ (
    .CLK(clk_bF$buf9),
    .D(_0_[23]),
    .Q(_11909_[23])
);

DFFPOSX1 _23970_ (
    .CLK(clk_bF$buf8),
    .D(_0_[24]),
    .Q(_11909_[24])
);

DFFPOSX1 _23971_ (
    .CLK(clk_bF$buf7),
    .D(_0_[25]),
    .Q(_11909_[25])
);

DFFPOSX1 _23972_ (
    .CLK(clk_bF$buf6),
    .D(_0_[26]),
    .Q(_11909_[26])
);

DFFPOSX1 _23973_ (
    .CLK(clk_bF$buf5),
    .D(_0_[27]),
    .Q(_11909_[27])
);

DFFPOSX1 _23974_ (
    .CLK(clk_bF$buf4),
    .D(_0_[28]),
    .Q(_11909_[28])
);

DFFPOSX1 _23975_ (
    .CLK(clk_bF$buf3),
    .D(_0_[29]),
    .Q(_11909_[29])
);

DFFPOSX1 _23976_ (
    .CLK(clk_bF$buf2),
    .D(_0_[30]),
    .Q(_11909_[30])
);

DFFPOSX1 _23977_ (
    .CLK(clk_bF$buf1),
    .D(_0_[31]),
    .Q(_11909_[31])
);

DFFPOSX1 _23978_ (
    .CLK(clk_bF$buf0),
    .D(_0_[32]),
    .Q(_11909_[32])
);

DFFPOSX1 _23979_ (
    .CLK(clk_bF$buf10),
    .D(_0_[33]),
    .Q(_11909_[33])
);

DFFPOSX1 _23980_ (
    .CLK(clk_bF$buf9),
    .D(_0_[34]),
    .Q(_11909_[34])
);

DFFPOSX1 _23981_ (
    .CLK(clk_bF$buf8),
    .D(_0_[35]),
    .Q(_11909_[35])
);

DFFPOSX1 _23982_ (
    .CLK(clk_bF$buf7),
    .D(_0_[36]),
    .Q(_11909_[36])
);

DFFPOSX1 _23983_ (
    .CLK(clk_bF$buf6),
    .D(_0_[37]),
    .Q(_11909_[37])
);

DFFPOSX1 _23984_ (
    .CLK(clk_bF$buf5),
    .D(_0_[38]),
    .Q(_11909_[38])
);

DFFPOSX1 _23985_ (
    .CLK(clk_bF$buf4),
    .D(_0_[39]),
    .Q(_11909_[39])
);

DFFPOSX1 _23986_ (
    .CLK(clk_bF$buf3),
    .D(_0_[40]),
    .Q(_11909_[40])
);

DFFPOSX1 _23987_ (
    .CLK(clk_bF$buf2),
    .D(_0_[41]),
    .Q(_11909_[41])
);

DFFPOSX1 _23988_ (
    .CLK(clk_bF$buf1),
    .D(_0_[42]),
    .Q(_11909_[42])
);

DFFPOSX1 _23989_ (
    .CLK(clk_bF$buf0),
    .D(_0_[43]),
    .Q(_11909_[43])
);

DFFPOSX1 _23990_ (
    .CLK(clk_bF$buf10),
    .D(_0_[44]),
    .Q(_11909_[44])
);

DFFPOSX1 _23991_ (
    .CLK(clk_bF$buf9),
    .D(_0_[45]),
    .Q(_11909_[45])
);

DFFPOSX1 _23992_ (
    .CLK(clk_bF$buf8),
    .D(_0_[46]),
    .Q(_11909_[46])
);

DFFPOSX1 _23993_ (
    .CLK(clk_bF$buf7),
    .D(_0_[47]),
    .Q(_11909_[47])
);

DFFPOSX1 _23994_ (
    .CLK(clk_bF$buf6),
    .D(_0_[48]),
    .Q(_11909_[48])
);

DFFPOSX1 _23995_ (
    .CLK(clk_bF$buf5),
    .D(_0_[49]),
    .Q(_11909_[49])
);

DFFPOSX1 _23996_ (
    .CLK(clk_bF$buf4),
    .D(_0_[50]),
    .Q(_11909_[50])
);

DFFPOSX1 _23997_ (
    .CLK(clk_bF$buf3),
    .D(_0_[51]),
    .Q(_11909_[51])
);

DFFPOSX1 _23998_ (
    .CLK(clk_bF$buf2),
    .D(_0_[52]),
    .Q(_11909_[52])
);

DFFPOSX1 _23999_ (
    .CLK(clk_bF$buf1),
    .D(_0_[53]),
    .Q(_11909_[53])
);

DFFPOSX1 _24000_ (
    .CLK(clk_bF$buf0),
    .D(_0_[54]),
    .Q(_11909_[54])
);

DFFPOSX1 _24001_ (
    .CLK(clk_bF$buf10),
    .D(_0_[55]),
    .Q(_11909_[55])
);

DFFPOSX1 _24002_ (
    .CLK(clk_bF$buf9),
    .D(_0_[56]),
    .Q(_11909_[56])
);

DFFPOSX1 _24003_ (
    .CLK(clk_bF$buf8),
    .D(_0_[57]),
    .Q(_11909_[57])
);

DFFPOSX1 _24004_ (
    .CLK(clk_bF$buf7),
    .D(_0_[58]),
    .Q(_11909_[58])
);

DFFPOSX1 _24005_ (
    .CLK(clk_bF$buf6),
    .D(_0_[59]),
    .Q(_11909_[59])
);

DFFPOSX1 _24006_ (
    .CLK(clk_bF$buf5),
    .D(_0_[60]),
    .Q(_11909_[60])
);

DFFPOSX1 _24007_ (
    .CLK(clk_bF$buf4),
    .D(_0_[61]),
    .Q(_11909_[61])
);

DFFPOSX1 _24008_ (
    .CLK(clk_bF$buf3),
    .D(_0_[62]),
    .Q(_11909_[62])
);

DFFPOSX1 _24009_ (
    .CLK(clk_bF$buf2),
    .D(_0_[63]),
    .Q(_11909_[63])
);

DFFPOSX1 _24010_ (
    .CLK(clk_bF$buf1),
    .D(a[0]),
    .Q(areg[0])
);

DFFPOSX1 _24011_ (
    .CLK(clk_bF$buf0),
    .D(a[1]),
    .Q(areg[1])
);

DFFPOSX1 _24012_ (
    .CLK(clk_bF$buf10),
    .D(a[2]),
    .Q(areg[2])
);

DFFPOSX1 _24013_ (
    .CLK(clk_bF$buf9),
    .D(a[3]),
    .Q(areg[3])
);

DFFPOSX1 _24014_ (
    .CLK(clk_bF$buf8),
    .D(a[4]),
    .Q(areg[4])
);

DFFPOSX1 _24015_ (
    .CLK(clk_bF$buf7),
    .D(a[5]),
    .Q(areg[5])
);

DFFPOSX1 _24016_ (
    .CLK(clk_bF$buf6),
    .D(a[6]),
    .Q(areg[6])
);

DFFPOSX1 _24017_ (
    .CLK(clk_bF$buf5),
    .D(a[7]),
    .Q(areg[7])
);

DFFPOSX1 _24018_ (
    .CLK(clk_bF$buf4),
    .D(a[8]),
    .Q(areg[8])
);

DFFPOSX1 _24019_ (
    .CLK(clk_bF$buf3),
    .D(a[9]),
    .Q(areg[9])
);

DFFPOSX1 _24020_ (
    .CLK(clk_bF$buf2),
    .D(a[10]),
    .Q(areg[10])
);

DFFPOSX1 _24021_ (
    .CLK(clk_bF$buf1),
    .D(a[11]),
    .Q(areg[11])
);

DFFPOSX1 _24022_ (
    .CLK(clk_bF$buf0),
    .D(a[12]),
    .Q(areg[12])
);

DFFPOSX1 _24023_ (
    .CLK(clk_bF$buf10),
    .D(a[13]),
    .Q(areg[13])
);

DFFPOSX1 _24024_ (
    .CLK(clk_bF$buf9),
    .D(a[14]),
    .Q(areg[14])
);

DFFPOSX1 _24025_ (
    .CLK(clk_bF$buf8),
    .D(a[15]),
    .Q(areg[15])
);

DFFPOSX1 _24026_ (
    .CLK(clk_bF$buf7),
    .D(a[16]),
    .Q(areg[16])
);

DFFPOSX1 _24027_ (
    .CLK(clk_bF$buf6),
    .D(a[17]),
    .Q(areg[17])
);

DFFPOSX1 _24028_ (
    .CLK(clk_bF$buf5),
    .D(a[18]),
    .Q(areg[18])
);

DFFPOSX1 _24029_ (
    .CLK(clk_bF$buf4),
    .D(a[19]),
    .Q(areg[19])
);

DFFPOSX1 _24030_ (
    .CLK(clk_bF$buf3),
    .D(a[20]),
    .Q(areg[20])
);

DFFPOSX1 _24031_ (
    .CLK(clk_bF$buf2),
    .D(a[21]),
    .Q(areg[21])
);

DFFPOSX1 _24032_ (
    .CLK(clk_bF$buf1),
    .D(a[22]),
    .Q(areg[22])
);

DFFPOSX1 _24033_ (
    .CLK(clk_bF$buf0),
    .D(a[23]),
    .Q(areg[23])
);

DFFPOSX1 _24034_ (
    .CLK(clk_bF$buf10),
    .D(a[24]),
    .Q(areg[24])
);

DFFPOSX1 _24035_ (
    .CLK(clk_bF$buf9),
    .D(a[25]),
    .Q(areg[25])
);

DFFPOSX1 _24036_ (
    .CLK(clk_bF$buf8),
    .D(a[26]),
    .Q(areg[26])
);

DFFPOSX1 _24037_ (
    .CLK(clk_bF$buf7),
    .D(a[27]),
    .Q(areg[27])
);

DFFPOSX1 _24038_ (
    .CLK(clk_bF$buf6),
    .D(a[28]),
    .Q(areg[28])
);

DFFPOSX1 _24039_ (
    .CLK(clk_bF$buf5),
    .D(a[29]),
    .Q(areg[29])
);

DFFPOSX1 _24040_ (
    .CLK(clk_bF$buf4),
    .D(a[30]),
    .Q(areg[30])
);

DFFPOSX1 _24041_ (
    .CLK(clk_bF$buf3),
    .D(a[31]),
    .Q(areg[31])
);

DFFPOSX1 _24042_ (
    .CLK(clk_bF$buf2),
    .D(b[0]),
    .Q(breg[0])
);

DFFPOSX1 _24043_ (
    .CLK(clk_bF$buf1),
    .D(b[1]),
    .Q(breg[1])
);

DFFPOSX1 _24044_ (
    .CLK(clk_bF$buf0),
    .D(b[2]),
    .Q(breg[2])
);

DFFPOSX1 _24045_ (
    .CLK(clk_bF$buf10),
    .D(b[3]),
    .Q(breg[3])
);

DFFPOSX1 _24046_ (
    .CLK(clk_bF$buf9),
    .D(b[4]),
    .Q(breg[4])
);

DFFPOSX1 _24047_ (
    .CLK(clk_bF$buf8),
    .D(b[5]),
    .Q(breg[5])
);

DFFPOSX1 _24048_ (
    .CLK(clk_bF$buf7),
    .D(b[6]),
    .Q(breg[6])
);

DFFPOSX1 _24049_ (
    .CLK(clk_bF$buf6),
    .D(b[7]),
    .Q(breg[7])
);

DFFPOSX1 _24050_ (
    .CLK(clk_bF$buf5),
    .D(b[8]),
    .Q(breg[8])
);

DFFPOSX1 _24051_ (
    .CLK(clk_bF$buf4),
    .D(b[9]),
    .Q(breg[9])
);

DFFPOSX1 _24052_ (
    .CLK(clk_bF$buf3),
    .D(b[10]),
    .Q(breg[10])
);

DFFPOSX1 _24053_ (
    .CLK(clk_bF$buf2),
    .D(b[11]),
    .Q(breg[11])
);

DFFPOSX1 _24054_ (
    .CLK(clk_bF$buf1),
    .D(b[12]),
    .Q(breg[12])
);

DFFPOSX1 _24055_ (
    .CLK(clk_bF$buf0),
    .D(b[13]),
    .Q(breg[13])
);

DFFPOSX1 _24056_ (
    .CLK(clk_bF$buf10),
    .D(b[14]),
    .Q(breg[14])
);

DFFPOSX1 _24057_ (
    .CLK(clk_bF$buf9),
    .D(b[15]),
    .Q(breg[15])
);

DFFPOSX1 _24058_ (
    .CLK(clk_bF$buf8),
    .D(b[16]),
    .Q(breg[16])
);

DFFPOSX1 _24059_ (
    .CLK(clk_bF$buf7),
    .D(b[17]),
    .Q(breg[17])
);

DFFPOSX1 _24060_ (
    .CLK(clk_bF$buf6),
    .D(b[18]),
    .Q(breg[18])
);

DFFPOSX1 _24061_ (
    .CLK(clk_bF$buf5),
    .D(b[19]),
    .Q(breg[19])
);

DFFPOSX1 _24062_ (
    .CLK(clk_bF$buf4),
    .D(b[20]),
    .Q(breg[20])
);

DFFPOSX1 _24063_ (
    .CLK(clk_bF$buf3),
    .D(b[21]),
    .Q(breg[21])
);

DFFPOSX1 _24064_ (
    .CLK(clk_bF$buf2),
    .D(b[22]),
    .Q(breg[22])
);

DFFPOSX1 _24065_ (
    .CLK(clk_bF$buf1),
    .D(b[23]),
    .Q(breg[23])
);

DFFPOSX1 _24066_ (
    .CLK(clk_bF$buf0),
    .D(b[24]),
    .Q(breg[24])
);

DFFPOSX1 _24067_ (
    .CLK(clk_bF$buf10),
    .D(b[25]),
    .Q(breg[25])
);

DFFPOSX1 _24068_ (
    .CLK(clk_bF$buf9),
    .D(b[26]),
    .Q(breg[26])
);

DFFPOSX1 _24069_ (
    .CLK(clk_bF$buf8),
    .D(b[27]),
    .Q(breg[27])
);

DFFPOSX1 _24070_ (
    .CLK(clk_bF$buf7),
    .D(b[28]),
    .Q(breg[28])
);

DFFPOSX1 _24071_ (
    .CLK(clk_bF$buf6),
    .D(b[29]),
    .Q(breg[29])
);

DFFPOSX1 _24072_ (
    .CLK(clk_bF$buf5),
    .D(b[30]),
    .Q(breg[30])
);

DFFPOSX1 _24073_ (
    .CLK(clk_bF$buf4),
    .D(b[31]),
    .Q(breg[31])
);

endmodule
