/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module multiplier(
    inout vdd,
    inout gnd,
    input [15:0] a,
    input [15:0] b,
    input clk,
    output [31:0] y
);

wire [15:0] a ;
wire [15:0] b ;
wire _1677_ ;
wire _1257_ ;
wire [31:0] y ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _2712_ ;
wire _2521_ ;
wire _2101_ ;
wire _703_ ;
wire _1389_ ;
wire _2750_ ;
wire _2330_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _1198_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2424_ ;
wire _2004_ ;
wire _606_ ;
wire _2653_ ;
wire _2233_ ;
wire _1924_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _2462_ ;
wire _2042_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2518_ ;
wire _2691_ ;
wire _2271_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _2080_ ;
wire _929_ ;
wire _509_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2556_ ;
wire _2136_ ;
wire _1827_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _2594_ ;
wire _2174_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2459_ ;
wire _2039_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _1768_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire areg_7_bF$buf0 ;
wire areg_7_bF$buf1 ;
wire areg_7_bF$buf2 ;
wire areg_7_bF$buf3 ;
wire _16_ ;
wire _2803_ ;
wire _1195_ ;
wire _2612_ ;
wire _54_ ;
wire _2421_ ;
wire _2001_ ;
wire _603_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _1921_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _92_ ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2515_ ;
wire _870_ ;
wire _450_ ;
wire _2744_ ;
wire _2324_ ;
wire _926_ ;
wire _506_ ;
wire _2553_ ;
wire _2133_ ;
wire _1824_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _2782_ ;
wire _2362_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2418_ ;
wire _2591_ ;
wire _2171_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _1918_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2456_ ;
wire _2036_ ;
wire breg_5_bF$buf0 ;
wire breg_5_bF$buf1 ;
wire breg_5_bF$buf2 ;
wire breg_5_bF$buf3 ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _2494_ ;
wire _2074_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _1192_ ;
wire _2397_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _2703_ ;
wire _1095_ ;
wire _2512_ ;
wire _2741_ ;
wire _2321_ ;
wire _7_ ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _2550_ ;
wire _2130_ ;
wire _1821_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2415_ ;
wire areg_2_bF$buf0 ;
wire areg_2_bF$buf1 ;
wire areg_2_bF$buf2 ;
wire areg_2_bF$buf3 ;
wire areg_2_bF$buf4 ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _1915_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _2453_ ;
wire _2033_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _2509_ ;
wire _2682_ ;
wire _2262_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _2491_ ;
wire _2071_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2547_ ;
wire _2127_ ;
wire _1818_ ;
wire _729_ ;
wire _309_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _2394_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _1092_ ;
wire _2297_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _2603_ ;
wire _45_ ;
wire _2412_ ;
wire _2641_ ;
wire _2221_ ;
wire _1912_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _2450_ ;
wire _2030_ ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _2506_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _2544_ ;
wire _2124_ ;
wire _1815_ ;
wire _726_ ;
wire _306_ ;
wire _2773_ ;
wire _2353_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2409_ ;
wire _2582_ ;
wire _2162_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _2391_ ;
wire _1909_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2447_ ;
wire _2027_ ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _2294_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2579_ ;
wire _2159_ ;
wire [31:0] _1_ ;
wire _1183_ ;
wire _2388_ ;
wire breg_14_bF$buf0 ;
wire breg_14_bF$buf1 ;
wire breg_14_bF$buf2 ;
wire breg_14_bF$buf3 ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _2197_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _2503_ ;
wire _2732_ ;
wire _2312_ ;
wire _914_ ;
wire _2541_ ;
wire _2121_ ;
wire _1812_ ;
wire _723_ ;
wire _303_ ;
wire _2770_ ;
wire _2350_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2406_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _1906_ ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2444_ ;
wire _2024_ ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire _2673_ ;
wire _2253_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _2482_ ;
wire _2062_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2538_ ;
wire _2118_ ;
wire _2291_ ;
wire _1809_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2576_ ;
wire _2156_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _2385_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _2194_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2479_ ;
wire _2059_ ;
wire _1083_ ;
wire _2288_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2500_ ;
wire _2097_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _2403_ ;
wire _2632_ ;
wire _2212_ ;
wire _1903_ ;
wire _814_ ;
wire _74_ ;
wire _2441_ ;
wire _2021_ ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _2670_ ;
wire _2250_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2535_ ;
wire _2115_ ;
wire _1806_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _2764_ ;
wire _2344_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _2573_ ;
wire _2153_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _2382_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2438_ ;
wire _2018_ ;
wire _2191_ ;
wire _1709_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _1938_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2476_ ;
wire _2056_ ;
wire _1747_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _2285_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _2094_ ;
wire areg_11_bF$buf0 ;
wire areg_11_bF$buf1 ;
wire areg_11_bF$buf2 ;
wire areg_11_bF$buf3 ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire _2799_ ;
wire _2379_ ;
wire _2188_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2400_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _1900_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _2723_ ;
wire _2303_ ;
wire _905_ ;
wire _2532_ ;
wire _2112_ ;
wire _1803_ ;
wire _714_ ;
wire breg_7_bF$buf0 ;
wire breg_7_bF$buf1 ;
wire breg_7_bF$buf2 ;
wire breg_7_bF$buf3 ;
wire _2761_ ;
wire _2341_ ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2570_ ;
wire _2150_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2435_ ;
wire _2015_ ;
wire _1706_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _2473_ ;
wire _2053_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2529_ ;
wire _2109_ ;
wire _2282_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _2091_ ;
wire _1609_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2567_ ;
wire _2147_ ;
wire _1838_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _2796_ ;
wire _2376_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _2185_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire _2699_ ;
wire _2279_ ;
wire _2088_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire areg_4_bF$buf0 ;
wire areg_4_bF$buf1 ;
wire areg_4_bF$buf2 ;
wire areg_4_bF$buf3 ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _1800_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _2623_ ;
wire _2203_ ;
wire _805_ ;
wire _65_ ;
wire _2432_ ;
wire _2012_ ;
wire _1703_ ;
wire _614_ ;
wire _2661_ ;
wire _2241_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _2470_ ;
wire _2050_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2526_ ;
wire _2106_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _2564_ ;
wire _2144_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _2793_ ;
wire _2373_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2429_ ;
wire _2009_ ;
wire _2182_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _1929_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2467_ ;
wire _2047_ ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _2085_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _24_ ;
wire _2811_ ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _2523_ ;
wire _2103_ ;
wire _705_ ;
wire _2752_ ;
wire _2332_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _2561_ ;
wire _2141_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _2790_ ;
wire _2370_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2426_ ;
wire _2006_ ;
wire _608_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _1926_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _2464_ ;
wire _2044_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _2693_ ;
wire _2273_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _2082_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2558_ ;
wire _2138_ ;
wire _1829_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _2711_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2520_ ;
wire _2100_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _56_ ;
wire _2423_ ;
wire _2003_ ;
wire _605_ ;
wire _2652_ ;
wire _2232_ ;
wire _1923_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _2461_ ;
wire _2041_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2517_ ;
wire _2690_ ;
wire _2270_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _928_ ;
wire _508_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2555_ ;
wire _2135_ ;
wire _1826_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _2784_ ;
wire _2364_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _2593_ ;
wire _2173_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2458_ ;
wire _2038_ ;
wire _1729_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _1767_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire breg_11_bF$buf0 ;
wire breg_11_bF$buf1 ;
wire breg_11_bF$buf2 ;
wire breg_11_bF$buf3 ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _2802_ ;
wire _1194_ ;
wire _2399_ ;
wire _2611_ ;
wire _53_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2420_ ;
wire _2000_ ;
wire _602_ ;
wire [15:0] breg ;
wire _1288_ ;
wire _199_ ;
wire _1920_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _2514_ ;
wire _2743_ ;
wire _2323_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire _2552_ ;
wire _2132_ ;
wire _1823_ ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _2781_ ;
wire _2361_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2417_ ;
wire _2590_ ;
wire _2170_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire areg_13_bF$buf0 ;
wire areg_13_bF$buf1 ;
wire areg_13_bF$buf2 ;
wire areg_13_bF$buf3 ;
wire _1917_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2455_ ;
wire _2035_ ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _2493_ ;
wire _2073_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2549_ ;
wire _2129_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _2396_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire breg_9_bF$buf0 ;
wire breg_9_bF$buf1 ;
wire breg_9_bF$buf2 ;
wire breg_9_bF$buf3 ;
wire _1285_ ;
wire _196_ ;
wire _2702_ ;
wire _1094_ ;
wire _2299_ ;
wire _2511_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire [15:0] areg ;
wire _1188_ ;
wire _1820_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2414_ ;
wire _2643_ ;
wire _2223_ ;
wire _1914_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _2452_ ;
wire _2032_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _2508_ ;
wire _2681_ ;
wire _2261_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _2490_ ;
wire _2070_ ;
wire _919_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2546_ ;
wire _2126_ ;
wire _1817_ ;
wire _728_ ;
wire _308_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _2393_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2449_ ;
wire _2029_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _1758_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _2296_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _2602_ ;
wire _2199_ ;
wire _44_ ;
wire _2411_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _1911_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _2505_ ;
wire breg_4_bF$buf0 ;
wire breg_4_bF$buf1 ;
wire breg_4_bF$buf2 ;
wire breg_4_bF$buf3 ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _916_ ;
wire _2543_ ;
wire _2123_ ;
wire _1814_ ;
wire _725_ ;
wire _305_ ;
wire _2772_ ;
wire _2352_ ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2408_ ;
wire _2581_ ;
wire _2161_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _2390_ ;
wire _1908_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _2293_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2578_ ;
wire _2158_ ;
wire [15:0] _0_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _2387_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _2196_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _2502_ ;
wire _2099_ ;
wire _2731_ ;
wire _2311_ ;
wire _913_ ;
wire _1599_ ;
wire _1179_ ;
wire _2540_ ;
wire _2120_ ;
wire _1811_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2405_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _1905_ ;
wire _816_ ;
wire _76_ ;
wire _2443_ ;
wire _2023_ ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire _2672_ ;
wire _2252_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _2481_ ;
wire _2061_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2537_ ;
wire _2117_ ;
wire _2290_ ;
wire _1808_ ;
wire _719_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2575_ ;
wire _2155_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _2384_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _2193_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2478_ ;
wire _2058_ ;
wire _1749_ ;
wire _1329_ ;
wire _1082_ ;
wire _2287_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _2096_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _35_ ;
wire _2402_ ;
wire _2631_ ;
wire _2211_ ;
wire _1902_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _2440_ ;
wire _2020_ ;
wire _1711_ ;
wire _622_ ;
wire _202_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2534_ ;
wire _2114_ ;
wire _1805_ ;
wire _716_ ;
wire _2763_ ;
wire _2343_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2572_ ;
wire _2152_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _2381_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2437_ ;
wire _2017_ ;
wire _2190_ ;
wire _1708_ ;
wire breg_13_bF$buf0 ;
wire breg_13_bF$buf1 ;
wire breg_13_bF$buf2 ;
wire breg_13_bF$buf3 ;
wire _619_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _1937_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2475_ ;
wire _2055_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _2284_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _2093_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2569_ ;
wire _2149_ ;
wire _1593_ ;
wire _1173_ ;
wire _2798_ ;
wire _2378_ ;
wire _1649_ ;
wire _1229_ ;
wire _2187_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _2722_ ;
wire _2302_ ;
wire areg_15_bF$buf0 ;
wire areg_15_bF$buf1 ;
wire areg_15_bF$buf2 ;
wire areg_15_bF$buf3 ;
wire _904_ ;
wire _2531_ ;
wire _2111_ ;
wire _1802_ ;
wire _713_ ;
wire _1399_ ;
wire _2760_ ;
wire _2340_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire [31:0] _2816_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2434_ ;
wire _2014_ ;
wire _1705_ ;
wire _616_ ;
wire _2663_ ;
wire _2243_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _2472_ ;
wire _2052_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2528_ ;
wire _2108_ ;
wire _2281_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _2090_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2566_ ;
wire _2146_ ;
wire _1837_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _2795_ ;
wire _2375_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _2184_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2469_ ;
wire _2049_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2087_ ;
wire _1778_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _2813_ ;
wire _2622_ ;
wire _2202_ ;
wire _804_ ;
wire _64_ ;
wire _2431_ ;
wire _2011_ ;
wire _1702_ ;
wire _613_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire areg_8_bF$buf0 ;
wire areg_8_bF$buf1 ;
wire _2525_ ;
wire areg_8_bF$buf2 ;
wire _2105_ ;
wire areg_8_bF$buf3 ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2754_ ;
wire _2334_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _2563_ ;
wire _2143_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire areg_10_bF$buf0 ;
wire areg_10_bF$buf1 ;
wire areg_10_bF$buf2 ;
wire areg_10_bF$buf3 ;
wire _2792_ ;
wire _2372_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2428_ ;
wire _2008_ ;
wire _2181_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _1928_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _2466_ ;
wire _2046_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _2084_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _2713_ ;
wire _2522_ ;
wire _2102_ ;
wire _704_ ;
wire _2751_ ;
wire _2331_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _1199_ ;
wire _2560_ ;
wire _2140_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2425_ ;
wire _2005_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _1925_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _2463_ ;
wire _2043_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2519_ ;
wire _2692_ ;
wire _2272_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _2081_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2557_ ;
wire _2137_ ;
wire _1828_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire areg_3_bF$buf0 ;
wire areg_3_bF$buf1 ;
wire areg_3_bF$buf2 ;
wire areg_3_bF$buf3 ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _1196_ ;
wire _2613_ ;
wire _55_ ;
wire _2422_ ;
wire _2002_ ;
wire _604_ ;
wire _2651_ ;
wire _2231_ ;
wire _1922_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _93_ ;
wire _1099_ ;
wire _2460_ ;
wire _2040_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2516_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _2554_ ;
wire _2134_ ;
wire _1825_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _2783_ ;
wire _2363_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2419_ ;
wire _2592_ ;
wire _2172_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _1919_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2457_ ;
wire _2037_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _14_ ;
wire _2801_ ;
wire _1193_ ;
wire _2398_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _90_ ;
wire _1096_ ;
wire _2513_ ;
wire _2742_ ;
wire _2322_ ;
wire breg_15_bF$buf0 ;
wire breg_15_bF$buf1 ;
wire breg_15_bF$buf2 ;
wire breg_15_bF$buf3 ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _2551_ ;
wire _2131_ ;
wire _1822_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _2780_ ;
wire _2360_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2416_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _1916_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _2454_ ;
wire _2034_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _2683_ ;
wire _2263_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _2492_ ;
wire _2072_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2548_ ;
wire _2128_ ;
wire _1819_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _2395_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _2701_ ;
wire _1093_ ;
wire _2298_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2510_ ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _46_ ;
wire _2413_ ;
wire _2642_ ;
wire _2222_ ;
wire _1913_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _2451_ ;
wire _2031_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _2507_ ;
wire _2680_ ;
wire _2260_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _918_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2545_ ;
wire _2125_ ;
wire _1816_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _2774_ ;
wire _2354_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _2583_ ;
wire _2163_ ;
wire breg_10_bF$buf0 ;
wire breg_10_bF$buf1 ;
wire breg_10_bF$buf2 ;
wire breg_10_bF$buf3 ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _2392_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2448_ ;
wire _2028_ ;
wire _1719_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _1757_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _2295_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _2389_ ;
wire _2601_ ;
wire _2198_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2410_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _1910_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire _630_ ;
wire _210_ ;
wire _2504_ ;
wire _2733_ ;
wire _2313_ ;
wire _915_ ;
wire _2542_ ;
wire _2122_ ;
wire _1813_ ;
wire _724_ ;
wire _304_ ;
wire _2771_ ;
wire _2351_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2407_ ;
wire _2580_ ;
wire _2160_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _1907_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _2483_ ;
wire _2063_ ;
wire breg_8_bF$buf0 ;
wire breg_8_bF$buf1 ;
wire breg_8_bF$buf2 ;
wire breg_8_bF$buf3 ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2539_ ;
wire _2119_ ;
wire _2292_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _1619_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2577_ ;
wire _2157_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _2386_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _2195_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _1084_ ;
wire _2289_ ;
wire _2501_ ;
wire _2098_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _1810_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2404_ ;
wire _2633_ ;
wire _2213_ ;
wire _1904_ ;
wire _815_ ;
wire _75_ ;
wire _2442_ ;
wire _2022_ ;
wire _1713_ ;
wire _624_ ;
wire _204_ ;
wire areg_5_bF$buf0 ;
wire areg_5_bF$buf1 ;
wire areg_5_bF$buf2 ;
wire areg_5_bF$buf3 ;
wire _2671_ ;
wire _2251_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _2480_ ;
wire _2060_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2536_ ;
wire _2116_ ;
wire _1807_ ;
wire _718_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _2574_ ;
wire _2154_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _2383_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2439_ ;
wire _2019_ ;
wire _2192_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _1939_ ;
wire _1519_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2477_ ;
wire _2057_ ;
wire _1748_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _2286_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _2095_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire breg_3_bF$buf0 ;
wire breg_3_bF$buf1 ;
wire breg_3_bF$buf2 ;
wire breg_3_bF$buf3 ;
wire _2189_ ;
wire _34_ ;
wire _2401_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _1901_ ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _906_ ;
wire _2533_ ;
wire _2113_ ;
wire _1804_ ;
wire _715_ ;
wire _2762_ ;
wire _2342_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2571_ ;
wire _2151_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _2380_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2436_ ;
wire _2016_ ;
wire _1707_ ;
wire _618_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _2474_ ;
wire _2054_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _2283_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _2092_ ;
wire areg_0_bF$buf0 ;
wire areg_0_bF$buf1 ;
wire areg_0_bF$buf2 ;
wire areg_0_bF$buf3 ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2568_ ;
wire _2148_ ;
wire _1839_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _2797_ ;
wire _2377_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _2186_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _2089_ ;
wire _2721_ ;
wire _2301_ ;
wire _903_ ;
wire _1589_ ;
wire _1169_ ;
wire _2530_ ;
wire _2110_ ;
wire _1801_ ;
wire _712_ ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _806_ ;
wire _66_ ;
wire _2433_ ;
wire _2013_ ;
wire _1704_ ;
wire _615_ ;
wire _2662_ ;
wire _2242_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _2471_ ;
wire _2051_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2527_ ;
wire _2107_ ;
wire _2280_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2565_ ;
wire _2145_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _2794_ ;
wire _2374_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _2183_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2468_ ;
wire _2048_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _2086_ ;
wire _1777_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _2812_ ;
wire _2621_ ;
wire _2201_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _2430_ ;
wire _2010_ ;
wire _1701_ ;
wire _612_ ;
wire _1298_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire breg_12_bF$buf0 ;
wire breg_12_bF$buf1 ;
wire breg_12_bF$buf2 ;
wire breg_12_bF$buf3 ;
wire _650_ ;
wire _230_ ;
wire _2524_ ;
wire _2104_ ;
wire _706_ ;
wire _2753_ ;
wire _2333_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _2562_ ;
wire _2142_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _2791_ ;
wire _2371_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2427_ ;
wire _2007_ ;
wire _2180_ ;
wire _609_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _1927_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2465_ ;
wire _2045_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _2694_ ;
wire _2274_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _2083_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2559_ ;
wire _2139_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _1639_ ;
wire _1219_ ;
wire areg_14_bF$buf0 ;
wire areg_14_bF$buf1 ;
wire areg_14_bF$buf2 ;
wire areg_14_bF$buf3 ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf0)
);

BUFX2 BUFX2_insert103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf1)
);

BUFX2 BUFX2_insert102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf2)
);

BUFX2 BUFX2_insert101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf3)
);

BUFX2 BUFX2_insert100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf0)
);

BUFX2 BUFX2_insert99 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf1)
);

BUFX2 BUFX2_insert98 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf2)
);

BUFX2 BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf3)
);

BUFX2 BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf0)
);

BUFX2 BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf1)
);

BUFX2 BUFX2_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf2)
);

BUFX2 BUFX2_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf3)
);

BUFX2 BUFX2_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(breg_8_bF$buf0)
);

BUFX2 BUFX2_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(breg_8_bF$buf1)
);

BUFX2 BUFX2_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(breg_8_bF$buf2)
);

BUFX2 BUFX2_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(breg_8_bF$buf3)
);

BUFX2 BUFX2_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf0)
);

BUFX2 BUFX2_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf1)
);

BUFX2 BUFX2_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf2)
);

BUFX2 BUFX2_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf3)
);

BUFX2 BUFX2_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf0)
);

BUFX2 BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf1)
);

BUFX2 BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf2)
);

BUFX2 BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf3)
);

BUFX2 BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf0)
);

BUFX2 BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf1)
);

BUFX2 BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf2)
);

BUFX2 BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf3)
);

BUFX2 BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf4)
);

BUFX2 BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf0)
);

BUFX2 BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf1)
);

BUFX2 BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf2)
);

BUFX2 BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf3)
);

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf0)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf1)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf2)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf3)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf0)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf1)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf2)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf3)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf0)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf1)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf2)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf3)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf0)
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf1)
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf2)
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf3)
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf0)
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf1)
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf2)
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf3)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf0)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf1)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf2)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf3)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf0)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf1)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf2)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf3)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf0)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf1)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf2)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf3)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf0)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf1)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf2)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf3)
);

CLKBUF1 CLKBUF1_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf0)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf3)
);

INVX8 _2817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .Y(_2437_)
);

INVX4 _2818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(_2447_)
);

NOR2X1 _2819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2447_),
    .Y(_0_[0])
);

NAND3X1 _2820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_2_bF$buf4),
    .C(_0_[0]),
    .Y(_2468_)
);

INVX4 _2821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .Y(_2479_)
);

NAND2X1 _2822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[2]),
    .Y(_2490_)
);

OAI21X1 _2823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2479_),
    .C(_2490_),
    .Y(_2501_)
);

NAND2X1 _2824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2501_),
    .B(_2468_),
    .Y(_2512_)
);

INVX8 _2825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(_2523_)
);

INVX4 _2826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(_2534_)
);

NOR2X1 _2827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2534_),
    .Y(_2545_)
);

OAI21X1 _2828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2447_),
    .C(_2545_),
    .Y(_2556_)
);

XOR2X1 _2829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2512_),
    .B(_2556_),
    .Y(_1_[2])
);

NAND3X1 _2830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_0_[0]),
    .B(_2545_),
    .C(_2512_),
    .Y(_2587_)
);

INVX4 _2831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(_2597_)
);

NOR2X1 _2832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2523_),
    .Y(_2598_)
);

NAND2X1 _2833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_3_bF$buf3),
    .Y(_2609_)
);

NAND2X1 _2834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[1]),
    .Y(_2620_)
);

NAND2X1 _2835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_3_bF$buf3),
    .Y(_2631_)
);

NAND2X1 _2836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg_3_bF$buf2),
    .Y(_2642_)
);

OAI21X1 _2837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2534_),
    .C(_2642_),
    .Y(_2653_)
);

OAI21X1 _2838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2620_),
    .B(_2631_),
    .C(_2653_),
    .Y(_2664_)
);

XOR2X1 _2839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2664_),
    .B(_2609_),
    .Y(_2675_)
);

INVX1 _2840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .Y(_2686_)
);

OAI21X1 _2841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2512_),
    .B(_2686_),
    .C(_2468_),
    .Y(_2697_)
);

NOR2X1 _2842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2675_),
    .B(_2697_),
    .Y(_2708_)
);

AND2X2 _2843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2697_),
    .B(_2675_),
    .Y(_2729_)
);

NOR2X1 _2844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .B(_2729_),
    .Y(_2730_)
);

XNOR2X1 _2845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2730_),
    .B(_2598_),
    .Y(_2741_)
);

XOR2X1 _2846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2741_),
    .B(_2587_),
    .Y(_1_[3])
);

NOR2X1 _2847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2587_),
    .B(_2741_),
    .Y(_2761_)
);

INVX1 _2848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .Y(_2772_)
);

INVX1 _2849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2729_),
    .Y(_2783_)
);

OAI21X1 _2850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2708_),
    .B(_2772_),
    .C(_2783_),
    .Y(_2794_)
);

INVX1 _2851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2794_),
    .Y(_2805_)
);

NAND2X1 _2852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[1]),
    .Y(_2_)
);

NAND2X1 _2853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_4_bF$buf3),
    .Y(_13_)
);

INVX4 _2854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .Y(_24_)
);

INVX4 _2855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .Y(_35_)
);

OAI22X1 _2856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_35_),
    .C(_2523_),
    .D(_24_),
    .Y(_46_)
);

OAI21X1 _2857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_13_),
    .C(_46_),
    .Y(_57_)
);

NOR2X1 _2858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2620_),
    .B(_2631_),
    .Y(_68_)
);

NOR2X1 _2859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2609_),
    .B(_2664_),
    .Y(_79_)
);

INVX1 _2860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .Y(_90_)
);

NOR2X1 _2861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2534_),
    .B(_90_),
    .Y(_101_)
);

NAND2X1 _2862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_4_bF$buf3),
    .Y(_112_)
);

INVX4 _2863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .Y(_122_)
);

OAI22X1 _2864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_122_),
    .C(_2597_),
    .D(_2479_),
    .Y(_143_)
);

OAI21X1 _2865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2490_),
    .B(_112_),
    .C(_143_),
    .Y(_154_)
);

XNOR2X1 _2866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_101_),
    .Y(_155_)
);

OAI21X1 _2867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_79_),
    .C(_155_),
    .Y(_166_)
);

NOR2X1 _2868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_68_),
    .B(_79_),
    .Y(_177_)
);

INVX1 _2869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .Y(_188_)
);

XNOR2X1 _2870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_188_),
    .Y(_199_)
);

NAND2X1 _2871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_177_),
    .Y(_210_)
);

NAND2X1 _2872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_210_),
    .Y(_221_)
);

XNOR2X1 _2873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_57_),
    .Y(_232_)
);

NOR2X1 _2874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2805_),
    .B(_232_),
    .Y(_243_)
);

INVX2 _2875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_57_),
    .Y(_254_)
);

XNOR2X1 _2876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_254_),
    .Y(_265_)
);

NOR2X1 _2877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2794_),
    .B(_265_),
    .Y(_276_)
);

NOR2X1 _2878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_243_),
    .Y(_287_)
);

XOR2X1 _2879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_2761_),
    .Y(_1_[4])
);

NOR2X1 _2880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_13_),
    .Y(_307_)
);

NOR2X1 _2881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_177_),
    .Y(_318_)
);

AOI21X1 _2882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_210_),
    .C(_318_),
    .Y(_329_)
);

INVX1 _2883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .Y(_340_)
);

NAND2X1 _2884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .B(breg_4_bF$buf1),
    .Y(_351_)
);

NAND2X1 _2885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_5_bF$buf3),
    .Y(_362_)
);

NAND2X1 _2886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_4_bF$buf1),
    .Y(_373_)
);

XOR2X1 _2887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_373_),
    .Y(_384_)
);

XNOR2X1 _2888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_351_),
    .Y(_405_)
);

INVX2 _2889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .Y(_406_)
);

NOR2X1 _2890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2490_),
    .B(_112_),
    .Y(_417_)
);

AOI21X1 _2891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_143_),
    .C(_417_),
    .Y(_428_)
);

INVX1 _2892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .Y(_439_)
);

NOR2X1 _2893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_90_),
    .Y(_450_)
);

NAND2X1 _2894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg_5_bF$buf3),
    .Y(_461_)
);

XOR2X1 _2895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_461_),
    .Y(_472_)
);

NAND2X1 _2896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(_472_),
    .Y(_483_)
);

INVX1 _2897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .Y(_493_)
);

NOR2X1 _2898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_461_),
    .Y(_504_)
);

AND2X2 _2899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_461_),
    .Y(_515_)
);

OAI21X1 _2900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_504_),
    .C(_493_),
    .Y(_526_)
);

NAND3X1 _2901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(_483_),
    .C(_439_),
    .Y(_537_)
);

NAND2X1 _2902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_5_bF$buf2),
    .Y(_548_)
);

INVX4 _2903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .Y(_559_)
);

OAI21X1 _2904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_559_),
    .C(_2631_),
    .Y(_570_)
);

OAI21X1 _2905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2642_),
    .B(_548_),
    .C(_570_),
    .Y(_581_)
);

NOR2X1 _2906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_581_),
    .Y(_602_)
);

NOR2X1 _2907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(_472_),
    .Y(_613_)
);

OAI21X1 _2908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_602_),
    .C(_428_),
    .Y(_614_)
);

NAND2X1 _2909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_537_),
    .B(_614_),
    .Y(_625_)
);

NOR2X1 _2910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_625_),
    .Y(_636_)
);

INVX1 _2911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .Y(_647_)
);

NOR3X1 _2912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_428_),
    .C(_613_),
    .Y(_658_)
);

AOI21X1 _2913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_526_),
    .B(_483_),
    .C(_439_),
    .Y(_669_)
);

OAI21X1 _2914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_669_),
    .C(_406_),
    .Y(_680_)
);

NAND3X1 _2915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_680_),
    .C(_647_),
    .Y(_690_)
);

INVX1 _2916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .Y(_701_)
);

OAI21X1 _2917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_636_),
    .C(_329_),
    .Y(_712_)
);

NAND3X1 _2918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_712_),
    .C(_690_),
    .Y(_723_)
);

INVX2 _2919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .Y(_734_)
);

NOR3X1 _2920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_329_),
    .C(_701_),
    .Y(_745_)
);

AOI21X1 _2921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .B(_647_),
    .C(_340_),
    .Y(_756_)
);

OAI21X1 _2922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_745_),
    .C(_734_),
    .Y(_767_)
);

NAND2X1 _2923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_767_),
    .Y(_778_)
);

NAND2X1 _2924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2761_),
    .B(_287_),
    .Y(_789_)
);

OAI21X1 _2925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2805_),
    .B(_232_),
    .C(_789_),
    .Y(_800_)
);

XNOR2X1 _2926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_800_),
    .B(_778_),
    .Y(_1_[5])
);

OR2X2 _2927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .B(_778_),
    .Y(_821_)
);

NAND3X1 _2928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_723_),
    .C(_767_),
    .Y(_832_)
);

OAI21X1 _2929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_734_),
    .C(_690_),
    .Y(_843_)
);

NOR2X1 _2930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_559_),
    .Y(_863_)
);

NAND3X1 _2931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .B(breg_4_bF$buf0),
    .C(_384_),
    .Y(_864_)
);

OAI21X1 _2932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_373_),
    .C(_864_),
    .Y(_875_)
);

XNOR2X1 _2933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_863_),
    .Y(_886_)
);

OAI21X1 _2934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_669_),
    .C(_537_),
    .Y(_897_)
);

NAND2X1 _2935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[6]),
    .Y(_908_)
);

NAND2X1 _2936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_5_bF$buf2),
    .Y(_919_)
);

NOR2X1 _2937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_919_),
    .Y(_930_)
);

AOI22X1 _2938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_4_bF$buf0),
    .C(breg[1]),
    .D(areg_5_bF$buf1),
    .Y(_941_)
);

OAI21X1 _2939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(_941_),
    .C(_908_),
    .Y(_952_)
);

NOR2X1 _2940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_941_),
    .B(_930_),
    .Y(_963_)
);

NAND3X1 _2941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[6]),
    .C(_963_),
    .Y(_974_)
);

NAND2X1 _2942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .B(_974_),
    .Y(_985_)
);

AOI21X1 _2943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_450_),
    .B(_570_),
    .C(_504_),
    .Y(_996_)
);

NAND2X1 _2944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_3_bF$buf1),
    .Y(_1007_)
);

NAND2X1 _2945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[6]),
    .Y(_1018_)
);

NOR2X1 _2946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_1018_),
    .Y(_1029_)
);

AND2X2 _2947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_1018_),
    .Y(_1039_)
);

NOR3X1 _2948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .B(_1029_),
    .C(_1039_),
    .Y(_1050_)
);

INVX2 _2949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .Y(_1061_)
);

OR2X2 _2950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_1018_),
    .Y(_1072_)
);

INVX4 _2951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(_1083_)
);

OAI21X1 _2952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_1083_),
    .C(_112_),
    .Y(_1094_)
);

AOI21X1 _2953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1094_),
    .B(_1072_),
    .C(_1061_),
    .Y(_1115_)
);

NOR3X1 _2954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1115_),
    .B(_996_),
    .C(_1050_),
    .Y(_1126_)
);

INVX1 _2955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .Y(_1127_)
);

NAND3X1 _2956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1061_),
    .B(_1094_),
    .C(_1072_),
    .Y(_1138_)
);

OAI21X1 _2957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1039_),
    .B(_1029_),
    .C(_1007_),
    .Y(_1149_)
);

AOI21X1 _2958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1138_),
    .C(_1127_),
    .Y(_1160_)
);

NOR3X1 _2959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1160_),
    .B(_1126_),
    .C(_985_),
    .Y(_1171_)
);

XNOR2X1 _2960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .B(_908_),
    .Y(_1182_)
);

NAND3X1 _2961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1138_),
    .C(_1127_),
    .Y(_1193_)
);

OAI21X1 _2962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1050_),
    .B(_1115_),
    .C(_996_),
    .Y(_1203_)
);

AOI21X1 _2963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1203_),
    .B(_1193_),
    .C(_1182_),
    .Y(_1214_)
);

OAI21X1 _2964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1214_),
    .C(_897_),
    .Y(_1225_)
);

AOI21X1 _2965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_614_),
    .C(_658_),
    .Y(_1236_)
);

NAND3X1 _2966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1182_),
    .B(_1203_),
    .C(_1193_),
    .Y(_1247_)
);

OAI21X1 _2967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1160_),
    .B(_1126_),
    .C(_985_),
    .Y(_1258_)
);

NAND3X1 _2968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1258_),
    .C(_1236_),
    .Y(_1269_)
);

AOI21X1 _2969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(_1225_),
    .C(_886_),
    .Y(_1280_)
);

INVX1 _2970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1280_),
    .Y(_1291_)
);

NOR3X1 _2971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1214_),
    .C(_1236_),
    .Y(_1302_)
);

AOI21X1 _2972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1258_),
    .C(_897_),
    .Y(_1313_)
);

OAI21X1 _2973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1302_),
    .B(_1313_),
    .C(_886_),
    .Y(_1324_)
);

NAND3X1 _2974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1291_),
    .B(_1324_),
    .C(_843_),
    .Y(_1335_)
);

AOI21X1 _2975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_307_),
    .B(_712_),
    .C(_745_),
    .Y(_1346_)
);

INVX2 _2976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .Y(_1356_)
);

OAI21X1 _2977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(_1280_),
    .C(_1346_),
    .Y(_1367_)
);

NAND3X1 _2978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1335_),
    .C(_832_),
    .Y(_1378_)
);

INVX1 _2979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .Y(_1399_)
);

NAND3X1 _2980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_734_),
    .B(_712_),
    .C(_690_),
    .Y(_1400_)
);

OAI21X1 _2981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_745_),
    .C(_307_),
    .Y(_1411_)
);

AOI21X1 _2982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1400_),
    .B(_1411_),
    .C(_1399_),
    .Y(_1422_)
);

OAI21X1 _2983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(_1280_),
    .C(_843_),
    .Y(_1433_)
);

NAND3X1 _2984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1291_),
    .B(_1324_),
    .C(_1346_),
    .Y(_1444_)
);

NAND3X1 _2985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1444_),
    .C(_1422_),
    .Y(_1455_)
);

AOI21X1 _2986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1378_),
    .B(_1455_),
    .C(_821_),
    .Y(_1466_)
);

NOR2X1 _2987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_789_),
    .Y(_1477_)
);

NAND3X1 _2988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1335_),
    .C(_1422_),
    .Y(_1487_)
);

NAND3X1 _2989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1444_),
    .C(_832_),
    .Y(_1498_)
);

AOI21X1 _2990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1487_),
    .C(_1477_),
    .Y(_1509_)
);

NOR2X1 _2991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1509_),
    .B(_1466_),
    .Y(_1_[6])
);

NAND3X1 _2992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1487_),
    .C(_1477_),
    .Y(_1530_)
);

NOR3X1 _2993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1346_),
    .B(_1280_),
    .C(_1356_),
    .Y(_1541_)
);

NAND2X1 _2994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_875_),
    .Y(_1552_)
);

INVX2 _2995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .Y(_1563_)
);

NAND3X1 _2996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1258_),
    .C(_897_),
    .Y(_1574_)
);

OAI21X1 _2997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_886_),
    .C(_1574_),
    .Y(_1585_)
);

NAND2X1 _2998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_7_bF$buf3),
    .Y(_1596_)
);

NOR2X1 _2999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_1596_),
    .Y(_1607_)
);

INVX2 _3000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .Y(_1617_)
);

NAND2X1 _3001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_7_bF$buf2),
    .Y(_1628_)
);

OAI21X1 _3002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_1083_),
    .C(_1628_),
    .Y(_1639_)
);

AND2X2 _3003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_1639_),
    .Y(_1650_)
);

OAI21X1 _3004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_373_),
    .B(_919_),
    .C(_974_),
    .Y(_1661_)
);

XOR2X1 _3005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1650_),
    .Y(_1672_)
);

OAI21X1 _3006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .B(_1160_),
    .C(_1193_),
    .Y(_1683_)
);

INVX4 _3007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(_1694_)
);

NOR2X1 _3008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2534_),
    .B(_1694_),
    .Y(_1705_)
);

INVX1 _3009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .Y(_1725_)
);

XOR2X1 _3010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_13_),
    .B(_919_),
    .Y(_1736_)
);

XNOR2X1 _3011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1736_),
    .B(_1725_),
    .Y(_1737_)
);

OAI21X1 _3012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1039_),
    .B(_1007_),
    .C(_1072_),
    .Y(_1748_)
);

NAND2X1 _3013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_4_bF$buf3),
    .Y(_1759_)
);

INVX2 _3014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1759_),
    .Y(_1770_)
);

AND2X2 _3015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_5_bF$buf0),
    .Y(_1781_)
);

AND2X2 _3016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg_7_bF$buf3),
    .Y(_1792_)
);

NAND2X1 _3017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1781_),
    .B(_1792_),
    .Y(_1802_)
);

INVX4 _3018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .Y(_1813_)
);

OAI21X1 _3019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_1813_),
    .C(_548_),
    .Y(_1824_)
);

NAND3X1 _3020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(_1824_),
    .C(_1802_),
    .Y(_1835_)
);

NAND2X1 _3021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_7_bF$buf1),
    .Y(_1846_)
);

NOR2X1 _3022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_1846_),
    .Y(_1856_)
);

AOI21X1 _3023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg_7_bF$buf0),
    .C(_1781_),
    .Y(_1867_)
);

OAI21X1 _3024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1856_),
    .C(_1759_),
    .Y(_1878_)
);

NAND3X1 _3025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1748_),
    .B(_1835_),
    .C(_1878_),
    .Y(_1889_)
);

AOI21X1 _3026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1061_),
    .B(_1094_),
    .C(_1029_),
    .Y(_1900_)
);

OAI21X1 _3027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_559_),
    .C(_1792_),
    .Y(_1911_)
);

OAI21X1 _3028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_1813_),
    .C(_1781_),
    .Y(_1921_)
);

AOI21X1 _3029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1911_),
    .B(_1921_),
    .C(_1759_),
    .Y(_1932_)
);

AOI21X1 _3030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_1802_),
    .C(_1770_),
    .Y(_1943_)
);

OAI21X1 _3031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_1943_),
    .C(_1900_),
    .Y(_1954_)
);

NAND3X1 _3032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1889_),
    .B(_1954_),
    .C(_1737_),
    .Y(_1965_)
);

XNOR2X1 _3033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1736_),
    .B(_1705_),
    .Y(_1976_)
);

NOR3X1 _3034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1943_),
    .B(_1900_),
    .C(_1932_),
    .Y(_1986_)
);

AOI21X1 _3035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(_1878_),
    .C(_1748_),
    .Y(_1997_)
);

OAI21X1 _3036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1986_),
    .B(_1997_),
    .C(_1976_),
    .Y(_2008_)
);

NAND3X1 _3037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1965_),
    .B(_2008_),
    .C(_1683_),
    .Y(_2019_)
);

AOI21X1 _3038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1203_),
    .B(_1182_),
    .C(_1126_),
    .Y(_2029_)
);

OAI21X1 _3039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_1943_),
    .C(_1748_),
    .Y(_2040_)
);

NAND3X1 _3040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .B(_1835_),
    .C(_1878_),
    .Y(_2051_)
);

AOI21X1 _3041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2040_),
    .B(_2051_),
    .C(_1976_),
    .Y(_2061_)
);

AOI21X1 _3042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(_1889_),
    .C(_1737_),
    .Y(_2072_)
);

OAI21X1 _3043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2072_),
    .C(_2029_),
    .Y(_2081_)
);

NAND3X1 _3044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_2081_),
    .C(_2019_),
    .Y(_2082_)
);

XNOR2X1 _3045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1650_),
    .Y(_2083_)
);

NOR3X1 _3046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2072_),
    .C(_2029_),
    .Y(_2084_)
);

AOI21X1 _3047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_1965_),
    .C(_1683_),
    .Y(_2085_)
);

OAI21X1 _3048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2084_),
    .B(_2085_),
    .C(_2083_),
    .Y(_2086_)
);

NAND3X1 _3049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2082_),
    .B(_2086_),
    .C(_1585_),
    .Y(_2087_)
);

INVX1 _3050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .Y(_2088_)
);

OAI21X1 _3051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1214_),
    .C(_1236_),
    .Y(_2089_)
);

AOI21X1 _3052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2088_),
    .C(_1302_),
    .Y(_2090_)
);

NOR3X1 _3053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2083_),
    .C(_2084_),
    .Y(_2091_)
);

AOI21X1 _3054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2081_),
    .B(_2019_),
    .C(_1672_),
    .Y(_2092_)
);

OAI21X1 _3055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2092_),
    .C(_2090_),
    .Y(_2093_)
);

NAND3X1 _3056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1563_),
    .B(_2093_),
    .C(_2087_),
    .Y(_2094_)
);

NOR3X1 _3057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2092_),
    .C(_2090_),
    .Y(_2095_)
);

AOI21X1 _3058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2082_),
    .B(_2086_),
    .C(_1585_),
    .Y(_2096_)
);

OAI21X1 _3059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2095_),
    .B(_2096_),
    .C(_1552_),
    .Y(_2097_)
);

NAND3X1 _3060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .B(_1541_),
    .C(_2097_),
    .Y(_2098_)
);

NAND3X1 _3061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_2093_),
    .C(_2087_),
    .Y(_2099_)
);

OAI21X1 _3062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2095_),
    .B(_2096_),
    .C(_1563_),
    .Y(_2100_)
);

NAND3X1 _3063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_1335_),
    .C(_2100_),
    .Y(_2101_)
);

NAND3X1 _3064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2098_),
    .B(_1487_),
    .C(_2101_),
    .Y(_2102_)
);

AOI21X1 _3065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1433_),
    .B(_1444_),
    .C(_832_),
    .Y(_2103_)
);

NAND3X1 _3066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .B(_1335_),
    .C(_2097_),
    .Y(_2104_)
);

NAND3X1 _3067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_1541_),
    .C(_2100_),
    .Y(_2105_)
);

NAND3X1 _3068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2103_),
    .B(_2104_),
    .C(_2105_),
    .Y(_2106_)
);

AOI21X1 _3069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2106_),
    .B(_2102_),
    .C(_1530_),
    .Y(_2107_)
);

NAND3X1 _3070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2103_),
    .B(_2098_),
    .C(_2101_),
    .Y(_2108_)
);

NAND3X1 _3071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2104_),
    .B(_1487_),
    .C(_2105_),
    .Y(_2109_)
);

AOI21X1 _3072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2108_),
    .B(_2109_),
    .C(_1466_),
    .Y(_2110_)
);

NOR2X1 _3073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2110_),
    .Y(_1_[7])
);

AOI21X1 _3074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2104_),
    .B(_2105_),
    .C(_1487_),
    .Y(_2111_)
);

OAI21X1 _3075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_1552_),
    .C(_2087_),
    .Y(_2112_)
);

NAND2X1 _3076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1650_),
    .B(_1661_),
    .Y(_2113_)
);

OAI21X1 _3077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2083_),
    .C(_2019_),
    .Y(_2114_)
);

NAND2X1 _3078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_8_bF$buf3),
    .Y(_2115_)
);

INVX8 _3079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .Y(_2116_)
);

NAND2X1 _3080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_7_bF$buf1),
    .Y(_2117_)
);

OAI21X1 _3081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2116_),
    .C(_2117_),
    .Y(_2118_)
);

OAI21X1 _3082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1628_),
    .B(_2115_),
    .C(_2118_),
    .Y(_2119_)
);

OAI21X1 _3083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_1813_),
    .C(_2119_),
    .Y(_2120_)
);

NOR2X1 _3084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_1813_),
    .Y(_2121_)
);

NOR2X1 _3085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1628_),
    .B(_2115_),
    .Y(_2122_)
);

INVX2 _3086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .Y(_2123_)
);

NAND3X1 _3087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2121_),
    .B(_2118_),
    .C(_2123_),
    .Y(_2124_)
);

NOR2X1 _3088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_13_),
    .B(_919_),
    .Y(_2125_)
);

INVX2 _3089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .Y(_2126_)
);

OAI21X1 _3090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2126_),
    .C(_13_),
    .Y(_2127_)
);

AOI21X1 _3091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .B(_2127_),
    .C(_2125_),
    .Y(_2128_)
);

INVX1 _3092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2128_),
    .Y(_2129_)
);

NAND3X1 _3093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2124_),
    .B(_2120_),
    .C(_2129_),
    .Y(_2130_)
);

AOI21X1 _3094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2118_),
    .B(_2123_),
    .C(_2121_),
    .Y(_2131_)
);

INVX1 _3095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2121_),
    .Y(_2132_)
);

NOR2X1 _3096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2132_),
    .B(_2119_),
    .Y(_2133_)
);

OAI21X1 _3097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_2131_),
    .C(_2128_),
    .Y(_2134_)
);

NAND3X1 _3098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_2130_),
    .C(_2134_),
    .Y(_2135_)
);

NAND3X1 _3099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2128_),
    .B(_2124_),
    .C(_2120_),
    .Y(_2136_)
);

OAI21X1 _3100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2133_),
    .B(_2131_),
    .C(_2129_),
    .Y(_2137_)
);

NAND3X1 _3101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_2136_),
    .C(_2137_),
    .Y(_2138_)
);

NAND2X1 _3102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2135_),
    .B(_2138_),
    .Y(_2139_)
);

OAI21X1 _3103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1976_),
    .B(_1997_),
    .C(_1889_),
    .Y(_2140_)
);

NAND2X1 _3104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg[6]),
    .Y(_2141_)
);

INVX1 _3105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .Y(_2142_)
);

NAND2X1 _3106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_5_bF$buf3),
    .Y(_2143_)
);

NAND2X1 _3107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_4_bF$buf3),
    .Y(_2144_)
);

OR2X2 _3108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .B(_2144_),
    .Y(_2145_)
);

OAI21X1 _3109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_35_),
    .C(_2143_),
    .Y(_2146_)
);

NAND3X1 _3110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2146_),
    .C(_2145_),
    .Y(_2147_)
);

NOR2X1 _3111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .B(_2144_),
    .Y(_2148_)
);

AND2X2 _3112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .B(_2144_),
    .Y(_2149_)
);

OAI21X1 _3113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2149_),
    .B(_2148_),
    .C(_2141_),
    .Y(_2150_)
);

AND2X2 _3114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2147_),
    .B(_2150_),
    .Y(_2151_)
);

OAI21X1 _3115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1759_),
    .C(_1802_),
    .Y(_2152_)
);

NAND2X1 _3116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_5_bF$buf3),
    .Y(_2153_)
);

INVX2 _3117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2153_),
    .Y(_2154_)
);

AND2X2 _3118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg[6]),
    .Y(_2155_)
);

AND2X2 _3119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg_8_bF$buf3),
    .Y(_2156_)
);

NAND2X1 _3120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2155_),
    .B(_2156_),
    .Y(_2157_)
);

INVX4 _3121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf2),
    .Y(_2158_)
);

NAND2X1 _3122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg[6]),
    .Y(_2159_)
);

OAI21X1 _3123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2158_),
    .C(_2159_),
    .Y(_2160_)
);

NAND3X1 _3124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(_2160_),
    .C(_2157_),
    .Y(_2161_)
);

NAND2X1 _3125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg_8_bF$buf1),
    .Y(_2162_)
);

NOR2X1 _3126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2159_),
    .B(_2162_),
    .Y(_2163_)
);

NOR2X1 _3127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2155_),
    .B(_2156_),
    .Y(_2164_)
);

OAI21X1 _3128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2163_),
    .C(_2153_),
    .Y(_2165_)
);

NAND3X1 _3129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2152_),
    .C(_2165_),
    .Y(_2166_)
);

AOI21X1 _3130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(_1824_),
    .C(_1856_),
    .Y(_2167_)
);

OAI21X1 _3131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_1083_),
    .C(_2156_),
    .Y(_2168_)
);

OAI21X1 _3132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2158_),
    .C(_2155_),
    .Y(_2169_)
);

AOI21X1 _3133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2169_),
    .C(_2153_),
    .Y(_2170_)
);

AOI21X1 _3134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2157_),
    .C(_2154_),
    .Y(_2171_)
);

OAI21X1 _3135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .B(_2171_),
    .C(_2167_),
    .Y(_2172_)
);

NAND3X1 _3136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2151_),
    .B(_2166_),
    .C(_2172_),
    .Y(_2173_)
);

NAND2X1 _3137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2150_),
    .B(_2147_),
    .Y(_2174_)
);

NOR3X1 _3138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2167_),
    .C(_2170_),
    .Y(_2175_)
);

AOI21X1 _3139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2165_),
    .C(_2152_),
    .Y(_2176_)
);

OAI21X1 _3140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2175_),
    .B(_2176_),
    .C(_2174_),
    .Y(_2177_)
);

NAND3X1 _3141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2177_),
    .C(_2140_),
    .Y(_2178_)
);

AOI21X1 _3142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(_1737_),
    .C(_1986_),
    .Y(_2179_)
);

OAI21X1 _3143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .B(_2171_),
    .C(_2152_),
    .Y(_2180_)
);

NAND3X1 _3144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2161_),
    .C(_2165_),
    .Y(_2181_)
);

AOI21X1 _3145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2180_),
    .B(_2181_),
    .C(_2174_),
    .Y(_2182_)
);

AOI21X1 _3146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2166_),
    .C(_2151_),
    .Y(_2183_)
);

OAI21X1 _3147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2183_),
    .B(_2182_),
    .C(_2179_),
    .Y(_2184_)
);

NAND3X1 _3148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2178_),
    .C(_2139_),
    .Y(_2185_)
);

NAND3X1 _3149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_2130_),
    .C(_2134_),
    .Y(_2186_)
);

NAND3X1 _3150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_2136_),
    .C(_2137_),
    .Y(_2187_)
);

NAND2X1 _3151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2186_),
    .B(_2187_),
    .Y(_2188_)
);

NOR3X1 _3152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2183_),
    .C(_2179_),
    .Y(_2189_)
);

AOI21X1 _3153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2177_),
    .C(_2140_),
    .Y(_2190_)
);

OAI21X1 _3154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2189_),
    .B(_2190_),
    .C(_2188_),
    .Y(_2191_)
);

AOI21X1 _3155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2191_),
    .C(_2114_),
    .Y(_2192_)
);

AOI21X1 _3156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_2081_),
    .C(_2084_),
    .Y(_2193_)
);

OAI21X1 _3157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2183_),
    .B(_2182_),
    .C(_2140_),
    .Y(_2194_)
);

NAND3X1 _3158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2177_),
    .C(_2179_),
    .Y(_2195_)
);

AOI21X1 _3159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2194_),
    .B(_2195_),
    .C(_2188_),
    .Y(_2196_)
);

AOI21X1 _3160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2178_),
    .C(_2139_),
    .Y(_2197_)
);

NOR3X1 _3161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .B(_2197_),
    .C(_2193_),
    .Y(_2198_)
);

OAI21X1 _3162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2192_),
    .C(_2113_),
    .Y(_2199_)
);

INVX2 _3163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2113_),
    .Y(_2200_)
);

OAI21X1 _3164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2196_),
    .B(_2197_),
    .C(_2193_),
    .Y(_2201_)
);

NAND3X1 _3165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2114_),
    .B(_2185_),
    .C(_2191_),
    .Y(_2202_)
);

NAND3X1 _3166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .B(_2201_),
    .C(_2202_),
    .Y(_2203_)
);

NAND3X1 _3167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2203_),
    .B(_2199_),
    .C(_2112_),
    .Y(_2204_)
);

AOI21X1 _3168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1563_),
    .B(_2093_),
    .C(_2095_),
    .Y(_2205_)
);

AOI21X1 _3169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2201_),
    .B(_2202_),
    .C(_2200_),
    .Y(_2206_)
);

NOR3X1 _3170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2192_),
    .B(_2113_),
    .C(_2198_),
    .Y(_2207_)
);

OAI21X1 _3171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2206_),
    .C(_2205_),
    .Y(_2208_)
);

NAND3X1 _3172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2204_),
    .B(_2208_),
    .C(_2098_),
    .Y(_2209_)
);

AOI21X1 _3173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_2100_),
    .C(_1335_),
    .Y(_2210_)
);

OAI21X1 _3174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2206_),
    .C(_2112_),
    .Y(_2211_)
);

NAND3X1 _3175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .B(_2203_),
    .C(_2205_),
    .Y(_2212_)
);

NAND3X1 _3176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2212_),
    .B(_2211_),
    .C(_2210_),
    .Y(_2213_)
);

AOI21X1 _3177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2213_),
    .C(_2111_),
    .Y(_2214_)
);

AOI21X1 _3178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2212_),
    .B(_2211_),
    .C(_2210_),
    .Y(_2215_)
);

AOI21X1 _3179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2204_),
    .B(_2208_),
    .C(_2098_),
    .Y(_2216_)
);

NOR3X1 _3180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2108_),
    .B(_2216_),
    .C(_2215_),
    .Y(_2217_)
);

NOR2X1 _3181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2214_),
    .B(_2217_),
    .Y(_2218_)
);

XNOR2X1 _3182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .B(_2107_),
    .Y(_1_[8])
);

NAND3X1 _3183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2108_),
    .B(_2109_),
    .C(_1466_),
    .Y(_2219_)
);

OAI21X1 _3184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2215_),
    .B(_2216_),
    .C(_2111_),
    .Y(_2220_)
);

OAI21X1 _3185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2218_),
    .B(_2219_),
    .C(_2220_),
    .Y(_2221_)
);

AOI21X1 _3186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(_2212_),
    .C(_2098_),
    .Y(_2222_)
);

NOR3X1 _3187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2206_),
    .C(_2205_),
    .Y(_2223_)
);

OAI21X1 _3188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2192_),
    .B(_2113_),
    .C(_2202_),
    .Y(_2224_)
);

NOR2X1 _3189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2158_),
    .Y(_2225_)
);

NAND2X1 _3190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2130_),
    .B(_2186_),
    .Y(_2226_)
);

XOR2X1 _3191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2225_),
    .Y(_2227_)
);

OAI21X1 _3192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2188_),
    .C(_2178_),
    .Y(_2228_)
);

OAI21X1 _3193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2119_),
    .B(_2132_),
    .C(_2123_),
    .Y(_2229_)
);

INVX1 _3194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .Y(_2230_)
);

NAND2X1 _3195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[9]),
    .Y(_2231_)
);

NAND2X1 _3196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_8_bF$buf1),
    .Y(_2232_)
);

NOR2X1 _3197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2117_),
    .B(_2232_),
    .Y(_2233_)
);

NAND2X1 _3198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_7_bF$buf0),
    .Y(_2234_)
);

AND2X2 _3199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2234_),
    .Y(_2235_)
);

OAI21X1 _3200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2233_),
    .C(_2231_),
    .Y(_2236_)
);

INVX1 _3201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .Y(_2237_)
);

OR2X2 _3202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2234_),
    .Y(_2238_)
);

INVX8 _3203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .Y(_2239_)
);

OAI21X1 _3204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2239_),
    .C(_2115_),
    .Y(_2240_)
);

NAND3X1 _3205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .B(_2240_),
    .C(_2238_),
    .Y(_2241_)
);

OAI21X1 _3206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2149_),
    .B(_2141_),
    .C(_2145_),
    .Y(_2242_)
);

NAND3X1 _3207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2242_),
    .B(_2241_),
    .C(_2236_),
    .Y(_2243_)
);

AOI21X1 _3208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2238_),
    .C(_2237_),
    .Y(_2244_)
);

NOR3X1 _3209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2233_),
    .C(_2235_),
    .Y(_2245_)
);

AOI21X1 _3210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2146_),
    .C(_2148_),
    .Y(_2246_)
);

OAI21X1 _3211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2245_),
    .B(_2244_),
    .C(_2246_),
    .Y(_2247_)
);

NAND3X1 _3212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .B(_2247_),
    .C(_2230_),
    .Y(_2248_)
);

NAND3X1 _3213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .B(_2236_),
    .C(_2241_),
    .Y(_2249_)
);

OAI21X1 _3214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2245_),
    .B(_2244_),
    .C(_2242_),
    .Y(_2250_)
);

NAND3X1 _3215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2249_),
    .C(_2250_),
    .Y(_2251_)
);

NAND2X1 _3216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2248_),
    .Y(_2252_)
);

OAI21X1 _3217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .B(_2174_),
    .C(_2166_),
    .Y(_2253_)
);

NOR2X1 _3218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_1694_),
    .Y(_2254_)
);

AND2X2 _3219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_4_bF$buf2),
    .Y(_2255_)
);

AND2X2 _3220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_5_bF$buf2),
    .Y(_2256_)
);

AOI22X1 _3221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_5_bF$buf1),
    .C(areg_4_bF$buf1),
    .D(breg_5_bF$buf1),
    .Y(_2257_)
);

AOI21X1 _3222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2255_),
    .B(_2256_),
    .C(_2257_),
    .Y(_2258_)
);

XOR2X1 _3223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2254_),
    .Y(_2259_)
);

OAI21X1 _3224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2153_),
    .C(_2157_),
    .Y(_2260_)
);

NAND2X1 _3225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg[6]),
    .Y(_2261_)
);

INVX2 _3226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .Y(_2262_)
);

AND2X2 _3227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_7_bF$buf3),
    .Y(_2263_)
);

AND2X2 _3228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg_9_bF$buf3),
    .Y(_2264_)
);

NAND2X1 _3229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2264_),
    .Y(_2265_)
);

INVX8 _3230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf2),
    .Y(_2266_)
);

OAI21X1 _3231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2266_),
    .C(_1846_),
    .Y(_2267_)
);

NAND3X1 _3232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2267_),
    .C(_2265_),
    .Y(_2268_)
);

NAND2X1 _3233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg_9_bF$buf1),
    .Y(_2269_)
);

NOR2X1 _3234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1846_),
    .B(_2269_),
    .Y(_2270_)
);

NOR2X1 _3235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2264_),
    .Y(_2271_)
);

OAI21X1 _3236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .B(_2270_),
    .C(_2261_),
    .Y(_2272_)
);

NAND3X1 _3237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2268_),
    .B(_2260_),
    .C(_2272_),
    .Y(_2273_)
);

AOI21X1 _3238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(_2160_),
    .C(_2163_),
    .Y(_2274_)
);

OAI21X1 _3239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_1813_),
    .C(_2264_),
    .Y(_2275_)
);

OAI21X1 _3240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2266_),
    .C(_2263_),
    .Y(_2276_)
);

AOI21X1 _3241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2275_),
    .B(_2276_),
    .C(_2261_),
    .Y(_2277_)
);

AOI21X1 _3242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2267_),
    .B(_2265_),
    .C(_2262_),
    .Y(_2278_)
);

OAI21X1 _3243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2277_),
    .B(_2278_),
    .C(_2274_),
    .Y(_2279_)
);

NAND3X1 _3244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2259_),
    .B(_2279_),
    .C(_2273_),
    .Y(_2280_)
);

XNOR2X1 _3245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2254_),
    .Y(_2281_)
);

OAI21X1 _3246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2277_),
    .B(_2278_),
    .C(_2260_),
    .Y(_2282_)
);

NAND3X1 _3247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2274_),
    .B(_2268_),
    .C(_2272_),
    .Y(_2283_)
);

NAND3X1 _3248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2281_),
    .B(_2282_),
    .C(_2283_),
    .Y(_2284_)
);

NAND3X1 _3249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2280_),
    .B(_2284_),
    .C(_2253_),
    .Y(_2285_)
);

AOI21X1 _3250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2151_),
    .C(_2175_),
    .Y(_2286_)
);

AOI21X1 _3251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2282_),
    .B(_2283_),
    .C(_2281_),
    .Y(_2287_)
);

AOI21X1 _3252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2279_),
    .B(_2273_),
    .C(_2259_),
    .Y(_2288_)
);

OAI21X1 _3253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2287_),
    .C(_2286_),
    .Y(_2289_)
);

NAND3X1 _3254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .B(_2285_),
    .C(_2289_),
    .Y(_2290_)
);

AND2X2 _3255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2248_),
    .B(_2251_),
    .Y(_2291_)
);

OAI21X1 _3256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2287_),
    .C(_2253_),
    .Y(_2292_)
);

NAND3X1 _3257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2284_),
    .B(_2280_),
    .C(_2286_),
    .Y(_2293_)
);

NAND3X1 _3258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2292_),
    .C(_2291_),
    .Y(_2294_)
);

NAND3X1 _3259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2290_),
    .B(_2294_),
    .C(_2228_),
    .Y(_2295_)
);

AOI21X1 _3260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2139_),
    .B(_2184_),
    .C(_2189_),
    .Y(_2296_)
);

AOI21X1 _3261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2292_),
    .C(_2291_),
    .Y(_2297_)
);

AOI21X1 _3262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2285_),
    .B(_2289_),
    .C(_2252_),
    .Y(_2298_)
);

OAI21X1 _3263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2297_),
    .B(_2298_),
    .C(_2296_),
    .Y(_2299_)
);

NAND3X1 _3264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2299_),
    .C(_2295_),
    .Y(_2300_)
);

XNOR2X1 _3265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2225_),
    .Y(_2301_)
);

NOR3X1 _3266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2297_),
    .B(_2298_),
    .C(_2296_),
    .Y(_2302_)
);

AOI21X1 _3267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2290_),
    .B(_2294_),
    .C(_2228_),
    .Y(_2303_)
);

OAI21X1 _3268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2303_),
    .C(_2301_),
    .Y(_2304_)
);

NAND3X1 _3269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2224_),
    .C(_2304_),
    .Y(_2305_)
);

AOI21X1 _3270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .B(_2201_),
    .C(_2198_),
    .Y(_2306_)
);

NOR3X1 _3271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2301_),
    .B(_2303_),
    .C(_2302_),
    .Y(_2307_)
);

AOI21X1 _3272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2299_),
    .B(_2295_),
    .C(_2227_),
    .Y(_2308_)
);

OAI21X1 _3273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2308_),
    .C(_2306_),
    .Y(_2309_)
);

NAND3X1 _3274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2309_),
    .C(_2223_),
    .Y(_2310_)
);

NOR3X1 _3275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2306_),
    .B(_2308_),
    .C(_2307_),
    .Y(_2311_)
);

AOI21X1 _3276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2304_),
    .C(_2224_),
    .Y(_2312_)
);

OAI21X1 _3277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2312_),
    .C(_2204_),
    .Y(_2313_)
);

NAND3X1 _3278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2222_),
    .B(_2313_),
    .C(_2310_),
    .Y(_2314_)
);

NAND3X1 _3279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2204_),
    .B(_2208_),
    .C(_2210_),
    .Y(_2315_)
);

NAND3X1 _3280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2309_),
    .C(_2204_),
    .Y(_2316_)
);

OAI21X1 _3281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2312_),
    .C(_2223_),
    .Y(_2317_)
);

NAND3X1 _3282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2317_),
    .C(_2315_),
    .Y(_2318_)
);

NAND2X1 _3283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2314_),
    .Y(_2319_)
);

XNOR2X1 _3284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(_2319_),
    .Y(_1_[9])
);

OAI21X1 _3285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2215_),
    .B(_2216_),
    .C(_2108_),
    .Y(_2320_)
);

NAND3X1 _3286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2213_),
    .C(_2111_),
    .Y(_2321_)
);

AOI21X1 _3287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2321_),
    .B(_2320_),
    .C(_2219_),
    .Y(_2322_)
);

AND2X2 _3288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2318_),
    .Y(_2323_)
);

NAND2X1 _3289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2220_),
    .Y(_2324_)
);

AOI22X1 _3290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2324_),
    .C(_2322_),
    .D(_2323_),
    .Y(_2325_)
);

NAND2X1 _3291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2225_),
    .B(_2226_),
    .Y(_2326_)
);

INVX2 _3292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2326_),
    .Y(_2327_)
);

OAI21X1 _3293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .B(_2301_),
    .C(_2295_),
    .Y(_2328_)
);

NAND2X1 _3294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_10_bF$buf3),
    .Y(_2329_)
);

NAND2X1 _3295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_10_bF$buf2),
    .Y(_2330_)
);

OAI21X1 _3296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2266_),
    .C(_2330_),
    .Y(_2331_)
);

OAI21X1 _3297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_2329_),
    .C(_2331_),
    .Y(_2332_)
);

INVX2 _3298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .Y(_2333_)
);

NAND2X1 _3299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .B(_2247_),
    .Y(_2334_)
);

OAI21X1 _3300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2334_),
    .B(_2230_),
    .C(_2243_),
    .Y(_2335_)
);

XNOR2X1 _3301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2335_),
    .B(_2333_),
    .Y(_2336_)
);

INVX2 _3302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .Y(_2337_)
);

AOI21X1 _3303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2284_),
    .B(_2280_),
    .C(_2253_),
    .Y(_2338_)
);

OAI21X1 _3304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .B(_2338_),
    .C(_2285_),
    .Y(_2339_)
);

OAI21X1 _3305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2231_),
    .C(_2238_),
    .Y(_2340_)
);

INVX1 _3306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .Y(_2341_)
);

INVX4 _3307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(_2342_)
);

NOR2X1 _3308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2534_),
    .B(_2342_),
    .Y(_2343_)
);

INVX1 _3309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2232_),
    .Y(_2344_)
);

NAND2X1 _3310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_7_bF$buf2),
    .Y(_2345_)
);

INVX1 _3311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .Y(_2346_)
);

NAND2X1 _3312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2344_),
    .B(_2346_),
    .Y(_2347_)
);

OAI21X1 _3313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_2239_),
    .C(_2232_),
    .Y(_2348_)
);

NAND3X1 _3314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2343_),
    .B(_2348_),
    .C(_2347_),
    .Y(_2349_)
);

NAND2X1 _3315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .B(areg_8_bF$buf0),
    .Y(_2350_)
);

OAI21X1 _3316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2350_),
    .C(_2348_),
    .Y(_2351_)
);

OAI21X1 _3317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2534_),
    .B(_2342_),
    .C(_2351_),
    .Y(_2352_)
);

INVX1 _3318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .Y(_2353_)
);

NAND2X1 _3319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf0),
    .B(areg_5_bF$buf0),
    .Y(_2354_)
);

OAI22X1 _3320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .B(_2354_),
    .C(_2353_),
    .D(_2257_),
    .Y(_2355_)
);

NAND3X1 _3321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2355_),
    .C(_2352_),
    .Y(_2356_)
);

INVX1 _3322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2343_),
    .Y(_2357_)
);

OAI21X1 _3323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2116_),
    .C(_2346_),
    .Y(_2358_)
);

OAI21X1 _3324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_2239_),
    .C(_2344_),
    .Y(_2359_)
);

AOI21X1 _3325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2358_),
    .B(_2359_),
    .C(_2357_),
    .Y(_2360_)
);

AOI21X1 _3326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2348_),
    .B(_2347_),
    .C(_2343_),
    .Y(_2361_)
);

AOI22X1 _3327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2255_),
    .B(_2256_),
    .C(_2258_),
    .D(_2254_),
    .Y(_2362_)
);

OAI21X1 _3328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2361_),
    .C(_2362_),
    .Y(_2363_)
);

NAND3X1 _3329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .B(_2356_),
    .C(_2363_),
    .Y(_2364_)
);

NAND3X1 _3330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .B(_2349_),
    .C(_2352_),
    .Y(_2365_)
);

OAI21X1 _3331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2361_),
    .C(_2355_),
    .Y(_2366_)
);

NAND3X1 _3332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2365_),
    .C(_2366_),
    .Y(_2367_)
);

NAND2X1 _3333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2367_),
    .Y(_2368_)
);

AOI21X1 _3334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2268_),
    .B(_2272_),
    .C(_2260_),
    .Y(_2369_)
);

OAI21X1 _3335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2369_),
    .B(_2281_),
    .C(_2273_),
    .Y(_2370_)
);

NOR2X1 _3336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_1694_),
    .Y(_2371_)
);

NAND2X1 _3337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_5_bF$buf3),
    .Y(_2372_)
);

NAND2X1 _3338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg[6]),
    .Y(_2373_)
);

OAI21X1 _3339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_1083_),
    .C(_2354_),
    .Y(_2374_)
);

OAI21X1 _3340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .B(_2373_),
    .C(_2374_),
    .Y(_2375_)
);

XNOR2X1 _3341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2375_),
    .B(_2371_),
    .Y(_2376_)
);

OAI21X1 _3342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .B(_2261_),
    .C(_2265_),
    .Y(_2377_)
);

NAND2X1 _3343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_7_bF$buf2),
    .Y(_2378_)
);

INVX2 _3344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .Y(_2379_)
);

AND2X2 _3345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_10_bF$buf3),
    .Y(_2380_)
);

NAND2X1 _3346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(_2380_),
    .Y(_2381_)
);

AOI22X1 _3347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg_10_bF$buf2),
    .C(areg_2_bF$buf3),
    .D(breg_8_bF$buf0),
    .Y(_2382_)
);

INVX2 _3348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2382_),
    .Y(_2383_)
);

NAND3X1 _3349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2383_),
    .C(_2381_),
    .Y(_2384_)
);

NAND2X1 _3350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_10_bF$buf1),
    .Y(_2385_)
);

NOR2X1 _3351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2162_),
    .B(_2385_),
    .Y(_2386_)
);

OAI21X1 _3352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2382_),
    .C(_2378_),
    .Y(_2387_)
);

NAND3X1 _3353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_2384_),
    .C(_2377_),
    .Y(_2388_)
);

AOI21X1 _3354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2267_),
    .C(_2270_),
    .Y(_2389_)
);

NOR3X1 _3355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .B(_2382_),
    .C(_2386_),
    .Y(_2390_)
);

AOI21X1 _3356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2381_),
    .C(_2379_),
    .Y(_2391_)
);

OAI21X1 _3357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2390_),
    .C(_2389_),
    .Y(_2392_)
);

NAND3X1 _3358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2388_),
    .B(_2392_),
    .C(_2376_),
    .Y(_2393_)
);

INVX1 _3359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .Y(_2394_)
);

XNOR2X1 _3360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2375_),
    .B(_2394_),
    .Y(_2395_)
);

OAI21X1 _3361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2390_),
    .C(_2377_),
    .Y(_2396_)
);

NAND3X1 _3362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2389_),
    .B(_2387_),
    .C(_2384_),
    .Y(_2397_)
);

NAND3X1 _3363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2396_),
    .B(_2397_),
    .C(_2395_),
    .Y(_2398_)
);

NAND3X1 _3364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2393_),
    .B(_2398_),
    .C(_2370_),
    .Y(_2399_)
);

NOR3X1 _3365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .B(_2274_),
    .C(_2277_),
    .Y(_2400_)
);

AOI21X1 _3366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2279_),
    .B(_2259_),
    .C(_2400_),
    .Y(_2401_)
);

AOI21X1 _3367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2396_),
    .C(_2395_),
    .Y(_2402_)
);

AOI21X1 _3368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2388_),
    .C(_2376_),
    .Y(_2403_)
);

OAI21X1 _3369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .B(_2402_),
    .C(_2401_),
    .Y(_2404_)
);

NAND3X1 _3370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2399_),
    .B(_2404_),
    .C(_2368_),
    .Y(_2405_)
);

NAND3X1 _3371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2356_),
    .C(_2363_),
    .Y(_2406_)
);

NAND3X1 _3372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .B(_2365_),
    .C(_2366_),
    .Y(_2407_)
);

NAND2X1 _3373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2406_),
    .B(_2407_),
    .Y(_2408_)
);

OAI21X1 _3374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .B(_2402_),
    .C(_2370_),
    .Y(_2409_)
);

NAND3X1 _3375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2393_),
    .C(_2401_),
    .Y(_2410_)
);

NAND3X1 _3376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2409_),
    .C(_2408_),
    .Y(_2411_)
);

NAND3X1 _3377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2411_),
    .C(_2339_),
    .Y(_2412_)
);

NOR3X1 _3378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2287_),
    .C(_2286_),
    .Y(_2413_)
);

AOI21X1 _3379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .B(_2289_),
    .C(_2413_),
    .Y(_2414_)
);

AOI21X1 _3380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2409_),
    .C(_2408_),
    .Y(_2415_)
);

AOI21X1 _3381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2399_),
    .B(_2404_),
    .C(_2368_),
    .Y(_2416_)
);

OAI21X1 _3382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2416_),
    .C(_2414_),
    .Y(_2417_)
);

NAND3X1 _3383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2412_),
    .C(_2417_),
    .Y(_2418_)
);

OAI21X1 _3384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2416_),
    .C(_2339_),
    .Y(_2419_)
);

NAND3X1 _3385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2411_),
    .C(_2414_),
    .Y(_2420_)
);

NAND3X1 _3386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2419_),
    .C(_2420_),
    .Y(_2421_)
);

NAND3X1 _3387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2418_),
    .B(_2421_),
    .C(_2328_),
    .Y(_2422_)
);

AOI21X1 _3388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2299_),
    .C(_2302_),
    .Y(_2423_)
);

AOI21X1 _3389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .B(_2420_),
    .C(_2336_),
    .Y(_2424_)
);

AOI21X1 _3390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2412_),
    .B(_2417_),
    .C(_2337_),
    .Y(_2425_)
);

OAI21X1 _3391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2425_),
    .C(_2423_),
    .Y(_2426_)
);

NAND3X1 _3392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2422_),
    .C(_2426_),
    .Y(_2427_)
);

OAI21X1 _3393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2425_),
    .C(_2328_),
    .Y(_2428_)
);

NAND3X1 _3394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2418_),
    .B(_2421_),
    .C(_2423_),
    .Y(_2429_)
);

NAND3X1 _3395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2326_),
    .B(_2428_),
    .C(_2429_),
    .Y(_2430_)
);

NAND3X1 _3396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2427_),
    .C(_2430_),
    .Y(_2431_)
);

NAND3X1 _3397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2326_),
    .B(_2422_),
    .C(_2426_),
    .Y(_2432_)
);

NAND3X1 _3398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2428_),
    .C(_2429_),
    .Y(_2433_)
);

NAND3X1 _3399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2432_),
    .C(_2433_),
    .Y(_2434_)
);

NAND3X1 _3400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2310_),
    .B(_2431_),
    .C(_2434_),
    .Y(_2435_)
);

NOR3X1 _3401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2204_),
    .B(_2312_),
    .C(_2311_),
    .Y(_2436_)
);

NAND3X1 _3402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2427_),
    .C(_2430_),
    .Y(_2438_)
);

NAND3X1 _3403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2432_),
    .C(_2433_),
    .Y(_2439_)
);

NAND3X1 _3404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2438_),
    .C(_2439_),
    .Y(_2440_)
);

NAND2X1 _3405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2440_),
    .Y(_2441_)
);

XNOR2X1 _3406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2441_),
    .Y(_1_[10])
);

NAND2X1 _3407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2434_),
    .Y(_2442_)
);

OR2X2 _3408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_2310_),
    .Y(_2443_)
);

AND2X2 _3409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2440_),
    .Y(_2444_)
);

OAI21X1 _3410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2444_),
    .C(_2443_),
    .Y(_2445_)
);

AOI21X1 _3411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .B(_2433_),
    .C(_2305_),
    .Y(_2446_)
);

AOI21X1 _3412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2418_),
    .B(_2421_),
    .C(_2328_),
    .Y(_2448_)
);

OAI21X1 _3413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2448_),
    .B(_2326_),
    .C(_2422_),
    .Y(_2449_)
);

NAND2X1 _3414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2333_),
    .B(_2335_),
    .Y(_2450_)
);

INVX2 _3415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2450_),
    .Y(_2451_)
);

AOI21X1 _3416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2411_),
    .C(_2339_),
    .Y(_2452_)
);

OAI21X1 _3417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_2336_),
    .C(_2412_),
    .Y(_2453_)
);

INVX2 _3418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .Y(_2454_)
);

NOR2X1 _3419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2454_),
    .Y(_2455_)
);

INVX1 _3420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .Y(_2456_)
);

NAND2X1 _3421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_11_bF$buf3),
    .Y(_2457_)
);

INVX4 _3422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .Y(_2458_)
);

NAND2X1 _3423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_10_bF$buf1),
    .Y(_2459_)
);

OAI21X1 _3424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2458_),
    .C(_2459_),
    .Y(_2460_)
);

OAI21X1 _3425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2330_),
    .B(_2457_),
    .C(_2460_),
    .Y(_2461_)
);

XNOR2X1 _3426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(_2456_),
    .Y(_2462_)
);

OAI21X1 _3427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_2329_),
    .C(_2462_),
    .Y(_2463_)
);

NOR2X1 _3428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_2329_),
    .Y(_2464_)
);

INVX1 _3429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2464_),
    .Y(_2465_)
);

NOR2X1 _3430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .B(_2462_),
    .Y(_2466_)
);

INVX2 _3431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .Y(_2467_)
);

NAND2X1 _3432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2463_),
    .B(_2467_),
    .Y(_2469_)
);

AND2X2 _3433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2406_),
    .B(_2356_),
    .Y(_2470_)
);

XOR2X1 _3434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2470_),
    .Y(_2471_)
);

AOI21X1 _3435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2393_),
    .C(_2370_),
    .Y(_2472_)
);

OAI21X1 _3436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2408_),
    .B(_2472_),
    .C(_2399_),
    .Y(_2473_)
);

OAI21X1 _3437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2357_),
    .C(_2347_),
    .Y(_2474_)
);

INVX2 _3438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .Y(_2475_)
);

NOR2X1 _3439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2342_),
    .Y(_2476_)
);

AND2X2 _3440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_8_bF$buf3),
    .Y(_2477_)
);

NAND2X1 _3441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2346_),
    .Y(_2478_)
);

OAI21X1 _3442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_2239_),
    .C(_2350_),
    .Y(_2480_)
);

NAND3X1 _3443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .B(_2480_),
    .C(_2478_),
    .Y(_2481_)
);

NAND2X1 _3444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_8_bF$buf2),
    .Y(_2482_)
);

OAI21X1 _3445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .B(_2482_),
    .C(_2480_),
    .Y(_2483_)
);

OAI21X1 _3446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2342_),
    .C(_2483_),
    .Y(_2484_)
);

NAND2X1 _3447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg[6]),
    .Y(_2485_)
);

NOR2X1 _3448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2354_),
    .B(_2485_),
    .Y(_2486_)
);

AOI21X1 _3449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .B(_2374_),
    .C(_2486_),
    .Y(_2487_)
);

INVX2 _3450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2487_),
    .Y(_2488_)
);

NAND3X1 _3451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .B(_2484_),
    .C(_2488_),
    .Y(_2489_)
);

INVX1 _3452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2476_),
    .Y(_2491_)
);

NOR2X1 _3453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2491_),
    .B(_2483_),
    .Y(_2492_)
);

AOI21X1 _3454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .B(_2478_),
    .C(_2476_),
    .Y(_2493_)
);

OAI21X1 _3455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2493_),
    .C(_2487_),
    .Y(_2494_)
);

NAND3X1 _3456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2489_),
    .C(_2494_),
    .Y(_2495_)
);

NAND3X1 _3457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2487_),
    .B(_2481_),
    .C(_2484_),
    .Y(_2496_)
);

OAI21X1 _3458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2493_),
    .C(_2488_),
    .Y(_2497_)
);

NAND3X1 _3459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2496_),
    .C(_2497_),
    .Y(_2498_)
);

NAND2X1 _3460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .B(_2498_),
    .Y(_2499_)
);

AOI21X1 _3461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_2384_),
    .C(_2377_),
    .Y(_2500_)
);

OAI21X1 _3462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2395_),
    .B(_2500_),
    .C(_2388_),
    .Y(_2502_)
);

NAND2X1 _3463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg[6]),
    .Y(_2503_)
);

INVX2 _3464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2503_),
    .Y(_2504_)
);

NAND2X1 _3465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_7_bF$buf1),
    .Y(_2505_)
);

OAI21X1 _3466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_1813_),
    .C(_2373_),
    .Y(_2506_)
);

OAI21X1 _3467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2485_),
    .B(_2505_),
    .C(_2506_),
    .Y(_2507_)
);

XNOR2X1 _3468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2504_),
    .Y(_2508_)
);

OAI21X1 _3469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .B(_2382_),
    .C(_2381_),
    .Y(_2509_)
);

NAND2X1 _3470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_8_bF$buf3),
    .Y(_2510_)
);

INVX2 _3471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .Y(_2511_)
);

AND2X2 _3472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_9_bF$buf3),
    .Y(_2513_)
);

AND2X2 _3473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg_11_bF$buf3),
    .Y(_2514_)
);

NAND2X1 _3474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2514_),
    .Y(_2515_)
);

NAND2X1 _3475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg_11_bF$buf2),
    .Y(_2516_)
);

OAI21X1 _3476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2266_),
    .C(_2516_),
    .Y(_2517_)
);

NAND3X1 _3477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_2517_),
    .C(_2515_),
    .Y(_2518_)
);

NAND2X1 _3478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_11_bF$buf1),
    .Y(_2519_)
);

NOR2X1 _3479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .B(_2519_),
    .Y(_2520_)
);

NOR2X1 _3480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2514_),
    .Y(_2521_)
);

OAI21X1 _3481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2521_),
    .B(_2520_),
    .C(_2510_),
    .Y(_2522_)
);

NAND3X1 _3482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2509_),
    .B(_2518_),
    .C(_2522_),
    .Y(_2524_)
);

AOI21X1 _3483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2383_),
    .C(_2386_),
    .Y(_2525_)
);

OAI21X1 _3484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2266_),
    .C(_2514_),
    .Y(_2526_)
);

INVX4 _3485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .Y(_2527_)
);

OAI21X1 _3486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2527_),
    .C(_2513_),
    .Y(_2528_)
);

AOI21X1 _3487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2526_),
    .B(_2528_),
    .C(_2510_),
    .Y(_2529_)
);

AOI21X1 _3488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2517_),
    .B(_2515_),
    .C(_2511_),
    .Y(_2530_)
);

OAI21X1 _3489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2529_),
    .B(_2530_),
    .C(_2525_),
    .Y(_2531_)
);

NAND3X1 _3490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2524_),
    .B(_2531_),
    .C(_2508_),
    .Y(_2532_)
);

XNOR2X1 _3491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2507_),
    .B(_2503_),
    .Y(_2533_)
);

NOR3X1 _3492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2525_),
    .C(_2529_),
    .Y(_2535_)
);

AOI21X1 _3493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2518_),
    .B(_2522_),
    .C(_2509_),
    .Y(_2536_)
);

OAI21X1 _3494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2535_),
    .B(_2536_),
    .C(_2533_),
    .Y(_2537_)
);

NAND3X1 _3495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2532_),
    .C(_2537_),
    .Y(_2538_)
);

NOR3X1 _3496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2389_),
    .C(_2391_),
    .Y(_2539_)
);

AOI21X1 _3497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2376_),
    .C(_2539_),
    .Y(_2540_)
);

OAI21X1 _3498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2529_),
    .B(_2530_),
    .C(_2509_),
    .Y(_2541_)
);

NAND3X1 _3499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2525_),
    .B(_2518_),
    .C(_2522_),
    .Y(_2542_)
);

AOI21X1 _3500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2541_),
    .B(_2542_),
    .C(_2533_),
    .Y(_2543_)
);

AOI21X1 _3501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2531_),
    .B(_2524_),
    .C(_2508_),
    .Y(_2544_)
);

OAI21X1 _3502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_2544_),
    .C(_2540_),
    .Y(_2546_)
);

NAND3X1 _3503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2538_),
    .C(_2499_),
    .Y(_2547_)
);

NAND3X1 _3504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2489_),
    .C(_2494_),
    .Y(_2548_)
);

NAND3X1 _3505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2496_),
    .C(_2497_),
    .Y(_2549_)
);

NAND2X1 _3506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2548_),
    .B(_2549_),
    .Y(_2550_)
);

NOR3X1 _3507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_2544_),
    .C(_2540_),
    .Y(_2551_)
);

AOI21X1 _3508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2537_),
    .C(_2502_),
    .Y(_2552_)
);

OAI21X1 _3509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_2552_),
    .C(_2550_),
    .Y(_2553_)
);

NAND3X1 _3510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2473_),
    .C(_2553_),
    .Y(_2554_)
);

NOR3X1 _3511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .B(_2402_),
    .C(_2401_),
    .Y(_2555_)
);

AOI21X1 _3512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_2368_),
    .C(_2555_),
    .Y(_2557_)
);

OAI21X1 _3513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_2544_),
    .C(_2502_),
    .Y(_2558_)
);

NAND3X1 _3514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_2532_),
    .C(_2537_),
    .Y(_2559_)
);

AOI21X1 _3515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2559_),
    .C(_2550_),
    .Y(_2560_)
);

AOI21X1 _3516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2538_),
    .C(_2499_),
    .Y(_2561_)
);

OAI21X1 _3517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2561_),
    .C(_2557_),
    .Y(_2562_)
);

NAND3X1 _3518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2471_),
    .B(_2562_),
    .C(_2554_),
    .Y(_2563_)
);

XNOR2X1 _3519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2470_),
    .Y(_2564_)
);

OAI21X1 _3520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2561_),
    .C(_2473_),
    .Y(_2565_)
);

NAND3X1 _3521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2557_),
    .B(_2547_),
    .C(_2553_),
    .Y(_2566_)
);

NAND3X1 _3522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2565_),
    .C(_2566_),
    .Y(_2567_)
);

NAND3X1 _3523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2453_),
    .B(_2563_),
    .C(_2567_),
    .Y(_2568_)
);

NOR3X1 _3524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2416_),
    .C(_2414_),
    .Y(_2569_)
);

AOI21X1 _3525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2417_),
    .C(_2569_),
    .Y(_2570_)
);

AOI21X1 _3526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2565_),
    .B(_2566_),
    .C(_2564_),
    .Y(_2571_)
);

AOI21X1 _3527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .B(_2554_),
    .C(_2471_),
    .Y(_2572_)
);

OAI21X1 _3528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2572_),
    .C(_2570_),
    .Y(_2573_)
);

NAND3X1 _3529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2568_),
    .C(_2573_),
    .Y(_2574_)
);

NOR3X1 _3530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2572_),
    .C(_2570_),
    .Y(_2575_)
);

AOI21X1 _3531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2567_),
    .B(_2563_),
    .C(_2453_),
    .Y(_2576_)
);

OAI21X1 _3532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2575_),
    .B(_2576_),
    .C(_2450_),
    .Y(_2577_)
);

NAND3X1 _3533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .B(_2574_),
    .C(_2577_),
    .Y(_2578_)
);

NOR3X1 _3534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2425_),
    .C(_2423_),
    .Y(_2579_)
);

AOI21X1 _3535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2426_),
    .C(_2579_),
    .Y(_2580_)
);

OAI21X1 _3536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2572_),
    .C(_2453_),
    .Y(_2581_)
);

NAND3X1 _3537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2563_),
    .B(_2567_),
    .C(_2570_),
    .Y(_2582_)
);

AOI21X1 _3538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2582_),
    .B(_2581_),
    .C(_2450_),
    .Y(_2583_)
);

AOI21X1 _3539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2568_),
    .B(_2573_),
    .C(_2451_),
    .Y(_2584_)
);

OAI21X1 _3540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2580_),
    .Y(_2585_)
);

NAND3X1 _3541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2446_),
    .B(_2585_),
    .C(_2578_),
    .Y(_2586_)
);

OAI21X1 _3542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2449_),
    .Y(_2588_)
);

NAND3X1 _3543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2580_),
    .B(_2574_),
    .C(_2577_),
    .Y(_2589_)
);

NAND3X1 _3544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2588_),
    .C(_2589_),
    .Y(_2590_)
);

NAND2X1 _3545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2590_),
    .Y(_2591_)
);

XNOR2X1 _3546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2591_),
    .Y(_1_[11])
);

NOR2X1 _3547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2310_),
    .B(_2442_),
    .Y(_2592_)
);

INVX1 _3548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2593_)
);

AOI21X1 _3549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2592_),
    .B(_2590_),
    .C(_2593_),
    .Y(_2594_)
);

NAND3X1 _3550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2590_),
    .C(_2441_),
    .Y(_2595_)
);

OAI21X1 _3551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2595_),
    .C(_2594_),
    .Y(_2596_)
);

NOR3X1 _3552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2580_),
    .Y(_2599_)
);

OAI21X1 _3553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2576_),
    .B(_2450_),
    .C(_2568_),
    .Y(_2600_)
);

NOR2X1 _3554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .B(_2469_),
    .Y(_2601_)
);

AOI21X1 _3555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2553_),
    .C(_2473_),
    .Y(_2602_)
);

OAI21X1 _3556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2602_),
    .B(_2564_),
    .C(_2554_),
    .Y(_2603_)
);

NOR2X1 _3557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2527_),
    .Y(_2604_)
);

NOR2X1 _3558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2330_),
    .B(_2457_),
    .Y(_2605_)
);

AOI21X1 _3559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2460_),
    .C(_2605_),
    .Y(_2606_)
);

INVX1 _3560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .Y(_2607_)
);

INVX4 _3561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(_2608_)
);

NOR2X1 _3562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2608_),
    .Y(_2610_)
);

NAND2X1 _3563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_10_bF$buf0),
    .Y(_2611_)
);

NOR2X1 _3564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_2611_),
    .Y(_2612_)
);

INVX1 _3565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2612_),
    .Y(_2613_)
);

INVX4 _3566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .Y(_2614_)
);

OAI21X1 _3567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2614_),
    .C(_2457_),
    .Y(_2615_)
);

NAND3X1 _3568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2615_),
    .C(_2613_),
    .Y(_2616_)
);

NAND2X1 _3569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_11_bF$buf1),
    .Y(_2617_)
);

OAI21X1 _3570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_2617_),
    .C(_2615_),
    .Y(_2618_)
);

OAI21X1 _3571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2608_),
    .C(_2618_),
    .Y(_2619_)
);

NAND3X1 _3572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2616_),
    .B(_2619_),
    .C(_2607_),
    .Y(_2621_)
);

INVX1 _3573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .Y(_2622_)
);

NOR2X1 _3574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2622_),
    .B(_2618_),
    .Y(_2623_)
);

AOI21X1 _3575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2615_),
    .B(_2613_),
    .C(_2610_),
    .Y(_2624_)
);

OAI21X1 _3576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2624_),
    .C(_2606_),
    .Y(_2625_)
);

NAND3X1 _3577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2621_),
    .C(_2625_),
    .Y(_2626_)
);

INVX1 _3578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .Y(_2627_)
);

OAI21X1 _3579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2624_),
    .C(_2607_),
    .Y(_2628_)
);

NAND3X1 _3580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(_2616_),
    .C(_2619_),
    .Y(_2629_)
);

NAND3X1 _3581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2627_),
    .B(_2629_),
    .C(_2628_),
    .Y(_2630_)
);

AOI21X1 _3582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2481_),
    .B(_2484_),
    .C(_2488_),
    .Y(_2632_)
);

OAI21X1 _3583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2632_),
    .B(_2475_),
    .C(_2489_),
    .Y(_2633_)
);

NAND3X1 _3584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2633_),
    .B(_2626_),
    .C(_2630_),
    .Y(_2634_)
);

AOI21X1 _3585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2629_),
    .B(_2628_),
    .C(_2627_),
    .Y(_2635_)
);

AOI21X1 _3586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2625_),
    .C(_2604_),
    .Y(_2636_)
);

NOR3X1 _3587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2493_),
    .B(_2487_),
    .C(_2492_),
    .Y(_2637_)
);

AOI21X1 _3588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2494_),
    .C(_2637_),
    .Y(_2638_)
);

OAI21X1 _3589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2635_),
    .C(_2638_),
    .Y(_2639_)
);

NAND3X1 _3590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2634_),
    .C(_2639_),
    .Y(_2640_)
);

NAND3X1 _3591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(_2630_),
    .C(_2638_),
    .Y(_2641_)
);

OAI21X1 _3592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2635_),
    .C(_2633_),
    .Y(_2643_)
);

NAND3X1 _3593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .B(_2641_),
    .C(_2643_),
    .Y(_2644_)
);

NAND2X1 _3594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2640_),
    .B(_2644_),
    .Y(_2645_)
);

OAI21X1 _3595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .B(_2550_),
    .C(_2538_),
    .Y(_2646_)
);

OAI21X1 _3596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2491_),
    .C(_2478_),
    .Y(_2647_)
);

NAND2X1 _3597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg[9]),
    .Y(_2648_)
);

AND2X2 _3598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg_7_bF$buf1),
    .Y(_2649_)
);

OAI21X1 _3599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_2116_),
    .C(_2649_),
    .Y(_2650_)
);

OAI21X1 _3600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2239_),
    .C(_2477_),
    .Y(_2651_)
);

AOI21X1 _3601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2650_),
    .B(_2651_),
    .C(_2648_),
    .Y(_2652_)
);

INVX1 _3602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .Y(_2654_)
);

NAND2X1 _3603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2649_),
    .Y(_2655_)
);

OAI21X1 _3604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2239_),
    .C(_2482_),
    .Y(_2656_)
);

AOI21X1 _3605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2656_),
    .B(_2655_),
    .C(_2654_),
    .Y(_2657_)
);

NAND2X1 _3606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_7_bF$buf0),
    .Y(_2658_)
);

NOR2X1 _3607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2658_),
    .Y(_2659_)
);

AOI21X1 _3608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(_2506_),
    .C(_2659_),
    .Y(_2660_)
);

OAI21X1 _3609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2657_),
    .C(_2660_),
    .Y(_2661_)
);

NAND3X1 _3610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2654_),
    .B(_2656_),
    .C(_2655_),
    .Y(_2662_)
);

NAND3X1 _3611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2648_),
    .B(_2650_),
    .C(_2651_),
    .Y(_2663_)
);

AND2X2 _3612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2658_),
    .Y(_2665_)
);

OAI22X1 _3613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2485_),
    .B(_2505_),
    .C(_2665_),
    .D(_2503_),
    .Y(_2666_)
);

NAND3X1 _3614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2662_),
    .B(_2663_),
    .C(_2666_),
    .Y(_2667_)
);

NAND3X1 _3615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .B(_2667_),
    .C(_2661_),
    .Y(_2668_)
);

INVX1 _3616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .Y(_2669_)
);

AOI21X1 _3617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2662_),
    .B(_2663_),
    .C(_2666_),
    .Y(_2670_)
);

NOR3X1 _3618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2657_),
    .B(_2660_),
    .C(_2652_),
    .Y(_2671_)
);

OAI21X1 _3619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2671_),
    .B(_2670_),
    .C(_2669_),
    .Y(_2672_)
);

AND2X2 _3620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .B(_2668_),
    .Y(_2673_)
);

OAI21X1 _3621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2533_),
    .B(_2536_),
    .C(_2524_),
    .Y(_2674_)
);

NAND2X1 _3622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg[6]),
    .Y(_2676_)
);

INVX2 _3623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .Y(_2677_)
);

NAND2X1 _3624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_8_bF$buf2),
    .Y(_2678_)
);

OAI21X1 _3625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_2158_),
    .C(_2505_),
    .Y(_2679_)
);

OAI21X1 _3626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2678_),
    .C(_2679_),
    .Y(_2680_)
);

XNOR2X1 _3627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .B(_2677_),
    .Y(_2681_)
);

OAI21X1 _3628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2521_),
    .B(_2510_),
    .C(_2515_),
    .Y(_2682_)
);

NAND2X1 _3629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_9_bF$buf2),
    .Y(_2683_)
);

INVX2 _3630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2683_),
    .Y(_2684_)
);

AND2X2 _3631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg_12_bF$buf3),
    .Y(_2685_)
);

NAND2X1 _3632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .B(_2685_),
    .Y(_2687_)
);

NAND2X1 _3633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg_12_bF$buf2),
    .Y(_2688_)
);

OAI21X1 _3634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2454_),
    .C(_2688_),
    .Y(_2689_)
);

NAND3X1 _3635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2689_),
    .C(_2687_),
    .Y(_2690_)
);

NOR2X1 _3636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2688_),
    .Y(_2691_)
);

NOR2X1 _3637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .B(_2685_),
    .Y(_2692_)
);

OAI21X1 _3638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2691_),
    .C(_2683_),
    .Y(_2693_)
);

NAND3X1 _3639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2690_),
    .B(_2693_),
    .C(_2682_),
    .Y(_2694_)
);

AOI21X1 _3640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2511_),
    .B(_2517_),
    .C(_2520_),
    .Y(_2695_)
);

OAI21X1 _3641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2454_),
    .C(_2685_),
    .Y(_2696_)
);

INVX2 _3642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .Y(_2698_)
);

OAI21X1 _3643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2698_),
    .C(_2380_),
    .Y(_2699_)
);

AOI21X1 _3644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2696_),
    .B(_2699_),
    .C(_2683_),
    .Y(_2700_)
);

AOI21X1 _3645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_2687_),
    .C(_2684_),
    .Y(_2701_)
);

OAI21X1 _3646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2701_),
    .C(_2695_),
    .Y(_2702_)
);

NAND3X1 _3647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2702_),
    .B(_2694_),
    .C(_2681_),
    .Y(_2703_)
);

XNOR2X1 _3648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .B(_2676_),
    .Y(_2704_)
);

OAI21X1 _3649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_2701_),
    .C(_2682_),
    .Y(_2705_)
);

NAND3X1 _3650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2695_),
    .B(_2690_),
    .C(_2693_),
    .Y(_2706_)
);

NAND3X1 _3651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2706_),
    .C(_2704_),
    .Y(_2707_)
);

NAND3X1 _3652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2707_),
    .C(_2674_),
    .Y(_2709_)
);

AOI21X1 _3653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2531_),
    .B(_2508_),
    .C(_2535_),
    .Y(_2710_)
);

AOI21X1 _3654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2706_),
    .C(_2704_),
    .Y(_2711_)
);

AOI21X1 _3655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2702_),
    .B(_2694_),
    .C(_2681_),
    .Y(_2712_)
);

OAI21X1 _3656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2711_),
    .C(_2710_),
    .Y(_2713_)
);

NAND3X1 _3657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2709_),
    .B(_2713_),
    .C(_2673_),
    .Y(_2714_)
);

NAND2X1 _3658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2668_),
    .B(_2672_),
    .Y(_2715_)
);

OAI21X1 _3659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2711_),
    .C(_2674_),
    .Y(_2716_)
);

NAND3X1 _3660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2707_),
    .C(_2710_),
    .Y(_2717_)
);

NAND3X1 _3661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2715_),
    .B(_2717_),
    .C(_2716_),
    .Y(_2718_)
);

NAND3X1 _3662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_2718_),
    .C(_2646_),
    .Y(_2719_)
);

AOI21X1 _3663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2499_),
    .C(_2551_),
    .Y(_2720_)
);

AOI21X1 _3664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2717_),
    .B(_2716_),
    .C(_2715_),
    .Y(_2721_)
);

AOI21X1 _3665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2709_),
    .B(_2713_),
    .C(_2673_),
    .Y(_2722_)
);

OAI21X1 _3666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2721_),
    .C(_2720_),
    .Y(_2723_)
);

NAND3X1 _3667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2719_),
    .B(_2723_),
    .C(_2645_),
    .Y(_2724_)
);

NAND3X1 _3668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .B(_2634_),
    .C(_2639_),
    .Y(_2725_)
);

NAND3X1 _3669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2641_),
    .C(_2643_),
    .Y(_2726_)
);

NAND2X1 _3670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .B(_2726_),
    .Y(_2727_)
);

NOR3X1 _3671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2721_),
    .C(_2720_),
    .Y(_2728_)
);

AOI21X1 _3672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2718_),
    .B(_2714_),
    .C(_2646_),
    .Y(_2731_)
);

OAI21X1 _3673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2728_),
    .B(_2731_),
    .C(_2727_),
    .Y(_2732_)
);

NAND3X1 _3674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2724_),
    .B(_2603_),
    .C(_2732_),
    .Y(_2733_)
);

NOR3X1 _3675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .B(_2561_),
    .C(_2557_),
    .Y(_2734_)
);

AOI21X1 _3676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .B(_2471_),
    .C(_2734_),
    .Y(_2735_)
);

OAI21X1 _3677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2721_),
    .C(_2646_),
    .Y(_2736_)
);

NAND3X1 _3678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2718_),
    .B(_2714_),
    .C(_2720_),
    .Y(_2737_)
);

AOI21X1 _3679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2737_),
    .C(_2727_),
    .Y(_2738_)
);

AOI21X1 _3680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2723_),
    .B(_2719_),
    .C(_2645_),
    .Y(_2739_)
);

OAI21X1 _3681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .B(_2738_),
    .C(_2735_),
    .Y(_2740_)
);

NAND3X1 _3682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2601_),
    .B(_2740_),
    .C(_2733_),
    .Y(_2742_)
);

INVX2 _3683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2601_),
    .Y(_2743_)
);

NOR3X1 _3684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .B(_2738_),
    .C(_2735_),
    .Y(_2744_)
);

AOI21X1 _3685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2724_),
    .B(_2732_),
    .C(_2603_),
    .Y(_2745_)
);

OAI21X1 _3686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_),
    .B(_2745_),
    .C(_2743_),
    .Y(_2746_)
);

NAND3X1 _3687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2600_),
    .B(_2742_),
    .C(_2746_),
    .Y(_2747_)
);

AOI21X1 _3688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2573_),
    .C(_2575_),
    .Y(_2748_)
);

OAI21X1 _3689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .B(_2738_),
    .C(_2603_),
    .Y(_2749_)
);

NAND3X1 _3690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2724_),
    .B(_2735_),
    .C(_2732_),
    .Y(_2750_)
);

AOI21X1 _3691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2749_),
    .B(_2750_),
    .C(_2743_),
    .Y(_2751_)
);

AOI21X1 _3692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2740_),
    .B(_2733_),
    .C(_2601_),
    .Y(_2752_)
);

OAI21X1 _3693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2751_),
    .B(_2752_),
    .C(_2748_),
    .Y(_2753_)
);

NAND3X1 _3694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2747_),
    .B(_2753_),
    .C(_2599_),
    .Y(_2754_)
);

OAI21X1 _3695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2751_),
    .B(_2752_),
    .C(_2600_),
    .Y(_2755_)
);

NAND3X1 _3696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2742_),
    .B(_2748_),
    .C(_2746_),
    .Y(_2756_)
);

NAND3X1 _3697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2755_),
    .B(_2756_),
    .C(_2578_),
    .Y(_2757_)
);

NAND2X1 _3698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2754_),
    .Y(_2758_)
);

XNOR2X1 _3699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(_2758_),
    .Y(_1_[12])
);

OAI21X1 _3700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2214_),
    .C(_2107_),
    .Y(_2759_)
);

NAND2X1 _3701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2324_),
    .Y(_2760_)
);

OAI21X1 _3702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2759_),
    .B(_2319_),
    .C(_2760_),
    .Y(_2762_)
);

OAI21X1 _3703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .B(_2443_),
    .C(_2586_),
    .Y(_2763_)
);

NOR2X1 _3704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .B(_2591_),
    .Y(_2764_)
);

AOI21X1 _3705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .B(_2762_),
    .C(_2763_),
    .Y(_2765_)
);

OAI21X1 _3706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2765_),
    .B(_2758_),
    .C(_2754_),
    .Y(_2766_)
);

NOR3X1 _3707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2751_),
    .B(_2752_),
    .C(_2748_),
    .Y(_2767_)
);

OAI21X1 _3708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2745_),
    .B(_2743_),
    .C(_2733_),
    .Y(_2768_)
);

NAND2X1 _3709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2634_),
    .B(_2725_),
    .Y(_2769_)
);

OAI21X1 _3710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .B(_2731_),
    .C(_2719_),
    .Y(_2770_)
);

AND2X2 _3711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(_2621_),
    .Y(_2771_)
);

NOR2X1 _3712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .B(_2608_),
    .Y(_2773_)
);

NAND2X1 _3713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .B(_2773_),
    .Y(_2774_)
);

NAND2X1 _3714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg[12]),
    .Y(_2775_)
);

OAI21X1 _3715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_2698_),
    .C(_2775_),
    .Y(_2776_)
);

NAND2X1 _3716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2776_),
    .B(_2774_),
    .Y(_2777_)
);

INVX1 _3717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2777_),
    .Y(_2778_)
);

AOI21X1 _3718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2615_),
    .C(_2612_),
    .Y(_2779_)
);

INVX1 _3719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .Y(_2780_)
);

INVX2 _3720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .Y(_2781_)
);

NOR2X1 _3721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2781_),
    .Y(_2782_)
);

NAND2X1 _3722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_10_bF$buf2),
    .Y(_2784_)
);

NOR2X1 _3723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2617_),
    .B(_2784_),
    .Y(_2785_)
);

INVX1 _3724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2785_),
    .Y(_2786_)
);

OAI21X1 _3725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_2614_),
    .C(_2617_),
    .Y(_2787_)
);

NAND3X1 _3726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2782_),
    .B(_2787_),
    .C(_2786_),
    .Y(_2788_)
);

NAND2X1 _3727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_11_bF$buf0),
    .Y(_2789_)
);

OAI21X1 _3728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .B(_2789_),
    .C(_2787_),
    .Y(_2790_)
);

OAI21X1 _3729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2781_),
    .C(_2790_),
    .Y(_2791_)
);

NAND3X1 _3730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2788_),
    .B(_2791_),
    .C(_2780_),
    .Y(_2792_)
);

INVX1 _3731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2782_),
    .Y(_2793_)
);

NOR2X1 _3732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2793_),
    .B(_2790_),
    .Y(_2795_)
);

AOI21X1 _3733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2787_),
    .B(_2786_),
    .C(_2782_),
    .Y(_2796_)
);

OAI21X1 _3734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2795_),
    .B(_2796_),
    .C(_2779_),
    .Y(_2797_)
);

NAND3X1 _3735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2778_),
    .B(_2792_),
    .C(_2797_),
    .Y(_2798_)
);

OAI21X1 _3736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2795_),
    .B(_2796_),
    .C(_2780_),
    .Y(_2799_)
);

NAND3X1 _3737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .B(_2788_),
    .C(_2791_),
    .Y(_2800_)
);

NAND3X1 _3738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2777_),
    .B(_2800_),
    .C(_2799_),
    .Y(_2801_)
);

OAI21X1 _3739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .B(_2670_),
    .C(_2667_),
    .Y(_2802_)
);

NAND3X1 _3740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2802_),
    .B(_2798_),
    .C(_2801_),
    .Y(_2803_)
);

AOI21X1 _3741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .B(_2799_),
    .C(_2777_),
    .Y(_2804_)
);

AOI21X1 _3742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_2797_),
    .C(_2778_),
    .Y(_2806_)
);

AOI21X1 _3743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2647_),
    .C(_2671_),
    .Y(_2807_)
);

OAI21X1 _3744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2804_),
    .B(_2806_),
    .C(_2807_),
    .Y(_2808_)
);

NAND3X1 _3745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2771_),
    .B(_2803_),
    .C(_2808_),
    .Y(_2809_)
);

NAND2X1 _3746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2626_),
    .Y(_2810_)
);

NAND3X1 _3747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .B(_2798_),
    .C(_2801_),
    .Y(_2811_)
);

OAI21X1 _3748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2804_),
    .B(_2806_),
    .C(_2802_),
    .Y(_2812_)
);

NAND3X1 _3749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(_2811_),
    .C(_2812_),
    .Y(_2813_)
);

NAND2X1 _3750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2809_),
    .B(_2813_),
    .Y(_2814_)
);

AOI21X1 _3751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2707_),
    .C(_2674_),
    .Y(_2815_)
);

OAI21X1 _3752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2815_),
    .B(_2715_),
    .C(_2709_),
    .Y(_3_)
);

NAND2X1 _3753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2662_),
    .Y(_4_)
);

NAND2X1 _3754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg[9]),
    .Y(_5_)
);

AND2X2 _3755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_7_bF$buf0),
    .Y(_6_)
);

OAI21X1 _3756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2116_),
    .C(_6_),
    .Y(_7_)
);

AND2X2 _3757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf0),
    .B(areg_8_bF$buf1),
    .Y(_8_)
);

OAI21X1 _3758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_2239_),
    .C(_8_),
    .Y(_9_)
);

AOI21X1 _3759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_9_),
    .C(_5_),
    .Y(_10_)
);

INVX1 _3760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5_),
    .Y(_11_)
);

NAND2X1 _3761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(_8_),
    .Y(_12_)
);

OAI21X1 _3762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2116_),
    .C(_1596_),
    .Y(_14_)
);

AOI21X1 _3763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(_12_),
    .C(_11_),
    .Y(_15_)
);

NAND2X1 _3764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_8_bF$buf1),
    .Y(_16_)
);

NOR2X1 _3765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2505_),
    .B(_16_),
    .Y(_17_)
);

AOI21X1 _3766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2679_),
    .C(_17_),
    .Y(_18_)
);

OAI21X1 _3767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(_15_),
    .C(_18_),
    .Y(_19_)
);

NAND3X1 _3768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11_),
    .B(_14_),
    .C(_12_),
    .Y(_20_)
);

NAND3X1 _3769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5_),
    .B(_7_),
    .C(_9_),
    .Y(_21_)
);

AND2X2 _3770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2505_),
    .B(_16_),
    .Y(_22_)
);

OAI22X1 _3771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2678_),
    .C(_22_),
    .D(_2676_),
    .Y(_23_)
);

NAND3X1 _3772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_20_),
    .B(_21_),
    .C(_23_),
    .Y(_25_)
);

NAND3X1 _3773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_25_),
    .C(_19_),
    .Y(_26_)
);

INVX1 _3774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .Y(_27_)
);

AOI21X1 _3775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_20_),
    .B(_21_),
    .C(_23_),
    .Y(_28_)
);

NOR3X1 _3776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_15_),
    .B(_18_),
    .C(_10_),
    .Y(_29_)
);

OAI21X1 _3777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_28_),
    .C(_27_),
    .Y(_30_)
);

AND2X2 _3778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_26_),
    .Y(_31_)
);

AOI21X1 _3779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2690_),
    .B(_2693_),
    .C(_2682_),
    .Y(_32_)
);

OAI21X1 _3780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_32_),
    .C(_2694_),
    .Y(_33_)
);

NOR2X1 _3781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_1813_),
    .Y(_34_)
);

NAND2X1 _3782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_9_bF$buf1),
    .Y(_36_)
);

NAND2X1 _3783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_9_bF$buf0),
    .Y(_37_)
);

OAI21X1 _3784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2158_),
    .C(_37_),
    .Y(_38_)
);

OAI21X1 _3785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_16_),
    .B(_36_),
    .C(_38_),
    .Y(_39_)
);

XNOR2X1 _3786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_34_),
    .Y(_40_)
);

OAI21X1 _3787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2683_),
    .C(_2687_),
    .Y(_41_)
);

NAND2X1 _3788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_10_bF$buf3),
    .Y(_42_)
);

INVX2 _3789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .Y(_43_)
);

AND2X2 _3790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_13_bF$buf3),
    .Y(_44_)
);

NAND2X1 _3791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .B(_44_),
    .Y(_45_)
);

NAND2X1 _3792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg_13_bF$buf2),
    .Y(_47_)
);

OAI21X1 _3793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2527_),
    .C(_47_),
    .Y(_48_)
);

NAND3X1 _3794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_48_),
    .C(_45_),
    .Y(_49_)
);

NAND2X1 _3795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_13_bF$buf1),
    .Y(_50_)
);

NOR2X1 _3796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .B(_50_),
    .Y(_51_)
);

AND2X2 _3797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_47_),
    .Y(_52_)
);

OAI21X1 _3798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_52_),
    .B(_51_),
    .C(_42_),
    .Y(_53_)
);

NAND3X1 _3799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .C(_41_),
    .Y(_54_)
);

AOI21X1 _3800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2689_),
    .C(_2691_),
    .Y(_55_)
);

NOR3X1 _3801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_51_),
    .C(_52_),
    .Y(_56_)
);

AOI21X1 _3802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_48_),
    .B(_45_),
    .C(_43_),
    .Y(_58_)
);

OAI21X1 _3803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_58_),
    .C(_55_),
    .Y(_59_)
);

NAND3X1 _3804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_59_),
    .C(_40_),
    .Y(_60_)
);

INVX1 _3805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .Y(_61_)
);

XNOR2X1 _3806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_61_),
    .Y(_62_)
);

OAI21X1 _3807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .B(_58_),
    .C(_41_),
    .Y(_63_)
);

NAND3X1 _3808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_49_),
    .C(_53_),
    .Y(_64_)
);

NAND3X1 _3809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_64_),
    .B(_63_),
    .C(_62_),
    .Y(_65_)
);

NAND3X1 _3810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_65_),
    .C(_33_),
    .Y(_66_)
);

NOR3X1 _3811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_2695_),
    .C(_2700_),
    .Y(_67_)
);

AOI21X1 _3812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2702_),
    .B(_2681_),
    .C(_67_),
    .Y(_69_)
);

AOI21X1 _3813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_64_),
    .B(_63_),
    .C(_62_),
    .Y(_70_)
);

AOI21X1 _3814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_59_),
    .C(_40_),
    .Y(_71_)
);

OAI21X1 _3815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_70_),
    .C(_69_),
    .Y(_72_)
);

NAND3X1 _3816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_72_),
    .C(_31_),
    .Y(_73_)
);

NAND2X1 _3817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_26_),
    .B(_30_),
    .Y(_74_)
);

NOR3X1 _3818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_70_),
    .C(_69_),
    .Y(_75_)
);

AOI21X1 _3819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_65_),
    .C(_33_),
    .Y(_76_)
);

OAI21X1 _3820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_76_),
    .C(_74_),
    .Y(_77_)
);

NAND3X1 _3821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3_),
    .B(_73_),
    .C(_77_),
    .Y(_78_)
);

NOR3X1 _3822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2711_),
    .C(_2710_),
    .Y(_80_)
);

AOI21X1 _3823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2713_),
    .B(_2673_),
    .C(_80_),
    .Y(_81_)
);

OAI21X1 _3824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_71_),
    .B(_70_),
    .C(_33_),
    .Y(_82_)
);

NAND3X1 _3825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_65_),
    .C(_69_),
    .Y(_83_)
);

AOI21X1 _3826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_83_),
    .B(_82_),
    .C(_74_),
    .Y(_84_)
);

AOI21X1 _3827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_72_),
    .C(_31_),
    .Y(_85_)
);

OAI21X1 _3828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_84_),
    .C(_81_),
    .Y(_86_)
);

NAND3X1 _3829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_2814_),
    .C(_78_),
    .Y(_87_)
);

NAND3X1 _3830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2810_),
    .B(_2803_),
    .C(_2808_),
    .Y(_88_)
);

NAND3X1 _3831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2771_),
    .B(_2811_),
    .C(_2812_),
    .Y(_89_)
);

NAND2X1 _3832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_89_),
    .Y(_91_)
);

NOR3X1 _3833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_84_),
    .C(_81_),
    .Y(_92_)
);

AOI21X1 _3834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_77_),
    .C(_3_),
    .Y(_93_)
);

OAI21X1 _3835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_93_),
    .C(_91_),
    .Y(_94_)
);

NAND3X1 _3836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2770_),
    .B(_87_),
    .C(_94_),
    .Y(_95_)
);

AOI21X1 _3837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2723_),
    .B(_2645_),
    .C(_2728_),
    .Y(_96_)
);

OAI21X1 _3838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_85_),
    .B(_84_),
    .C(_3_),
    .Y(_97_)
);

NAND3X1 _3839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_73_),
    .B(_81_),
    .C(_77_),
    .Y(_98_)
);

AOI21X1 _3840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_98_),
    .C(_91_),
    .Y(_99_)
);

AOI21X1 _3841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_78_),
    .C(_2814_),
    .Y(_100_)
);

OAI21X1 _3842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_100_),
    .C(_96_),
    .Y(_102_)
);

NAND3X1 _3843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2769_),
    .B(_102_),
    .C(_95_),
    .Y(_103_)
);

INVX2 _3844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2769_),
    .Y(_104_)
);

NOR3X1 _3845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_96_),
    .C(_100_),
    .Y(_105_)
);

AOI21X1 _3846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_94_),
    .C(_2770_),
    .Y(_106_)
);

OAI21X1 _3847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_106_),
    .C(_104_),
    .Y(_107_)
);

NAND3X1 _3848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_103_),
    .B(_2768_),
    .C(_107_),
    .Y(_108_)
);

AOI21X1 _3849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2601_),
    .B(_2740_),
    .C(_2744_),
    .Y(_109_)
);

OAI21X1 _3850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_100_),
    .C(_2770_),
    .Y(_110_)
);

NAND3X1 _3851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_96_),
    .C(_94_),
    .Y(_111_)
);

AOI21X1 _3852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_110_),
    .B(_111_),
    .C(_104_),
    .Y(_113_)
);

AOI21X1 _3853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_95_),
    .C(_2769_),
    .Y(_114_)
);

OAI21X1 _3854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_114_),
    .C(_109_),
    .Y(_115_)
);

NAND3X1 _3855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_115_),
    .C(_2767_),
    .Y(_116_)
);

OAI21X1 _3856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_114_),
    .C(_2768_),
    .Y(_117_)
);

NAND3X1 _3857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_103_),
    .C(_107_),
    .Y(_118_)
);

NAND3X1 _3858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2747_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

NAND2X1 _3859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_116_),
    .Y(_120_)
);

XNOR2X1 _3860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2766_),
    .B(_120_),
    .Y(_1_[13])
);

NAND2X1 _3861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2754_),
    .B(_116_),
    .Y(_121_)
);

NAND2X1 _3862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_121_),
    .Y(_123_)
);

INVX1 _3863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .Y(_124_)
);

NOR2X1 _3864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(_120_),
    .Y(_125_)
);

AOI21X1 _3865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(_2596_),
    .C(_124_),
    .Y(_126_)
);

OAI21X1 _3866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_106_),
    .B(_104_),
    .C(_95_),
    .Y(_127_)
);

INVX2 _3867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2774_),
    .Y(_128_)
);

NAND2X1 _3868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2803_),
    .B(_88_),
    .Y(_129_)
);

XNOR2X1 _3869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_128_),
    .Y(_130_)
);

INVX2 _3870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .Y(_131_)
);

OAI21X1 _3871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_91_),
    .C(_78_),
    .Y(_132_)
);

NAND2X1 _3872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_2798_),
    .Y(_133_)
);

NAND2X1 _3873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .B(breg_13_bF$buf0),
    .Y(_134_)
);

NAND2X1 _3874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg[12]),
    .Y(_135_)
);

NAND2X1 _3875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_13_bF$buf2),
    .Y(_136_)
);

XOR2X1 _3876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_136_),
    .Y(_137_)
);

XNOR2X1 _3877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_134_),
    .Y(_138_)
);

AOI21X1 _3878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2782_),
    .B(_2787_),
    .C(_2785_),
    .Y(_139_)
);

INVX1 _3879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .Y(_140_)
);

NAND2X1 _3880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_14_bF$buf3),
    .Y(_141_)
);

INVX2 _3881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .Y(_142_)
);

AND2X2 _3882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .B(areg_11_bF$buf3),
    .Y(_144_)
);

AND2X2 _3883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_10_bF$buf1),
    .Y(_145_)
);

NAND2X1 _3884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_145_),
    .Y(_146_)
);

NAND2X1 _3885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_10_bF$buf0),
    .Y(_147_)
);

OAI21X1 _3886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_2458_),
    .C(_147_),
    .Y(_148_)
);

NAND3X1 _3887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_148_),
    .C(_146_),
    .Y(_149_)
);

NOR2X1 _3888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2789_),
    .B(_147_),
    .Y(_150_)
);

NOR2X1 _3889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_145_),
    .Y(_151_)
);

OAI21X1 _3890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_150_),
    .C(_141_),
    .Y(_152_)
);

NAND3X1 _3891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_149_),
    .B(_152_),
    .C(_140_),
    .Y(_153_)
);

NOR3X1 _3892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_150_),
    .C(_151_),
    .Y(_156_)
);

AOI21X1 _3893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_146_),
    .C(_142_),
    .Y(_157_)
);

OAI21X1 _3894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_157_),
    .C(_139_),
    .Y(_158_)
);

NAND3X1 _3895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_158_),
    .C(_153_),
    .Y(_159_)
);

XOR2X1 _3896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_134_),
    .Y(_160_)
);

OAI21X1 _3897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_156_),
    .B(_157_),
    .C(_140_),
    .Y(_161_)
);

NAND3X1 _3898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_139_),
    .B(_149_),
    .C(_152_),
    .Y(_162_)
);

NAND3X1 _3899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_161_),
    .C(_160_),
    .Y(_163_)
);

OAI21X1 _3900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_28_),
    .C(_25_),
    .Y(_164_)
);

AOI21X1 _3901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_159_),
    .C(_164_),
    .Y(_165_)
);

AOI21X1 _3902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_161_),
    .C(_160_),
    .Y(_167_)
);

AOI21X1 _3903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_153_),
    .C(_138_),
    .Y(_168_)
);

AOI21X1 _3904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_19_),
    .C(_29_),
    .Y(_169_)
);

NOR3X1 _3905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_169_),
    .C(_168_),
    .Y(_170_)
);

OAI21X1 _3906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_165_),
    .C(_133_),
    .Y(_171_)
);

AND2X2 _3907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2798_),
    .B(_2792_),
    .Y(_172_)
);

OAI21X1 _3908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_167_),
    .C(_169_),
    .Y(_173_)
);

NAND3X1 _3909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_164_),
    .C(_159_),
    .Y(_174_)
);

NAND3X1 _3910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_175_)
);

NAND2X1 _3911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_171_),
    .Y(_176_)
);

OAI21X1 _3912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_74_),
    .C(_66_),
    .Y(_178_)
);

NAND2X1 _3913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_20_),
    .Y(_179_)
);

INVX2 _3914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .Y(_180_)
);

NOR2X1 _3915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2342_),
    .Y(_181_)
);

NAND2X1 _3916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_8_bF$buf0),
    .Y(_182_)
);

INVX1 _3917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .Y(_183_)
);

NAND2X1 _3918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(_183_),
    .Y(_184_)
);

NAND2X1 _3919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_7_bF$buf3),
    .Y(_185_)
);

OAI21X1 _3920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_2116_),
    .C(_185_),
    .Y(_186_)
);

NAND3X1 _3921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_186_),
    .C(_184_),
    .Y(_187_)
);

OAI21X1 _3922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_182_),
    .C(_186_),
    .Y(_189_)
);

OAI21X1 _3923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2342_),
    .C(_189_),
    .Y(_190_)
);

NOR2X1 _3924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2678_),
    .B(_37_),
    .Y(_191_)
);

AOI21X1 _3925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(_38_),
    .C(_191_),
    .Y(_192_)
);

INVX2 _3926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .Y(_193_)
);

NAND3X1 _3927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_190_),
    .C(_193_),
    .Y(_194_)
);

INVX1 _3928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .Y(_195_)
);

NOR2X1 _3929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_189_),
    .Y(_196_)
);

AOI21X1 _3930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_186_),
    .B(_184_),
    .C(_181_),
    .Y(_197_)
);

OAI21X1 _3931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_197_),
    .C(_192_),
    .Y(_198_)
);

NAND3X1 _3932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_194_),
    .C(_198_),
    .Y(_200_)
);

NAND3X1 _3933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_192_),
    .B(_187_),
    .C(_190_),
    .Y(_201_)
);

OAI21X1 _3934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_197_),
    .C(_193_),
    .Y(_202_)
);

NAND3X1 _3935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_201_),
    .C(_202_),
    .Y(_203_)
);

NAND2X1 _3936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_203_),
    .Y(_204_)
);

AOI21X1 _3937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .C(_41_),
    .Y(_205_)
);

OAI21X1 _3938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_205_),
    .C(_54_),
    .Y(_206_)
);

NOR2X1 _3939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_2158_),
    .Y(_207_)
);

NAND2X1 _3940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_10_bF$buf2),
    .Y(_208_)
);

NAND2X1 _3941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_10_bF$buf1),
    .Y(_209_)
);

OAI21X1 _3942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2266_),
    .C(_209_),
    .Y(_211_)
);

OAI21X1 _3943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .B(_208_),
    .C(_211_),
    .Y(_212_)
);

XNOR2X1 _3944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_207_),
    .Y(_213_)
);

OAI21X1 _3945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_52_),
    .B(_42_),
    .C(_45_),
    .Y(_214_)
);

NAND2X1 _3946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_11_bF$buf3),
    .Y(_215_)
);

INVX2 _3947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .Y(_216_)
);

NAND2X1 _3948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_12_bF$buf0),
    .Y(_217_)
);

NAND2X1 _3949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg_14_bF$buf3),
    .Y(_218_)
);

OR2X2 _3950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_218_),
    .Y(_219_)
);

INVX4 _3951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf2),
    .Y(_220_)
);

OAI21X1 _3952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_220_),
    .C(_217_),
    .Y(_222_)
);

NAND3X1 _3953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_222_),
    .C(_219_),
    .Y(_223_)
);

NAND2X1 _3954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_14_bF$buf1),
    .Y(_224_)
);

NOR2X1 _3955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .B(_224_),
    .Y(_225_)
);

AND2X2 _3956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_218_),
    .Y(_226_)
);

OAI21X1 _3957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_225_),
    .C(_215_),
    .Y(_227_)
);

NAND3X1 _3958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_223_),
    .C(_227_),
    .Y(_228_)
);

AOI21X1 _3959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_48_),
    .C(_51_),
    .Y(_229_)
);

NAND3X1 _3960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg_14_bF$buf0),
    .C(_217_),
    .Y(_230_)
);

NAND3X1 _3961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_12_bF$buf3),
    .C(_218_),
    .Y(_231_)
);

AOI21X1 _3962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_231_),
    .C(_215_),
    .Y(_233_)
);

AOI21X1 _3963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_219_),
    .C(_216_),
    .Y(_234_)
);

OAI21X1 _3964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_233_),
    .C(_229_),
    .Y(_235_)
);

NAND3X1 _3965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_235_),
    .C(_213_),
    .Y(_236_)
);

INVX1 _3966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .Y(_237_)
);

XNOR2X1 _3967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_212_),
    .B(_237_),
    .Y(_238_)
);

NOR3X1 _3968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_233_),
    .B(_229_),
    .C(_234_),
    .Y(_239_)
);

AOI21X1 _3969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_223_),
    .C(_214_),
    .Y(_240_)
);

OAI21X1 _3970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(_240_),
    .C(_238_),
    .Y(_241_)
);

NAND3X1 _3971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_206_),
    .C(_241_),
    .Y(_242_)
);

NOR3X1 _3972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_55_),
    .C(_56_),
    .Y(_244_)
);

AOI21X1 _3973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_40_),
    .C(_244_),
    .Y(_245_)
);

OAI21X1 _3974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_233_),
    .C(_214_),
    .Y(_246_)
);

NAND3X1 _3975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_227_),
    .C(_223_),
    .Y(_247_)
);

AOI21X1 _3976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_246_),
    .C(_238_),
    .Y(_248_)
);

AOI21X1 _3977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_228_),
    .B(_235_),
    .C(_213_),
    .Y(_249_)
);

OAI21X1 _3978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_249_),
    .C(_245_),
    .Y(_250_)
);

NAND3X1 _3979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_242_),
    .B(_250_),
    .C(_204_),
    .Y(_251_)
);

NAND3X1 _3980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_194_),
    .C(_198_),
    .Y(_252_)
);

NAND3X1 _3981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .B(_201_),
    .C(_202_),
    .Y(_253_)
);

NAND2X1 _3982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_252_),
    .B(_253_),
    .Y(_255_)
);

OAI21X1 _3983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_249_),
    .C(_206_),
    .Y(_256_)
);

NAND3X1 _3984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_245_),
    .C(_241_),
    .Y(_257_)
);

NAND3X1 _3985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_258_)
);

NAND3X1 _3986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_251_),
    .C(_258_),
    .Y(_259_)
);

AOI21X1 _3987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .B(_31_),
    .C(_75_),
    .Y(_260_)
);

AOI21X1 _3988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_256_),
    .B(_257_),
    .C(_255_),
    .Y(_261_)
);

AOI21X1 _3989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_242_),
    .C(_204_),
    .Y(_262_)
);

OAI21X1 _3990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_262_),
    .C(_260_),
    .Y(_263_)
);

NAND3X1 _3991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_263_),
    .C(_176_),
    .Y(_264_)
);

NAND3X1 _3992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_174_),
    .C(_173_),
    .Y(_266_)
);

OAI21X1 _3993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_165_),
    .C(_172_),
    .Y(_267_)
);

NAND2X1 _3994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_267_),
    .Y(_268_)
);

OAI21X1 _3995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_262_),
    .C(_178_),
    .Y(_269_)
);

NAND3X1 _3996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_258_),
    .C(_260_),
    .Y(_270_)
);

NAND3X1 _3997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_270_),
    .C(_268_),
    .Y(_271_)
);

NAND3X1 _3998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_271_),
    .C(_132_),
    .Y(_272_)
);

AOI21X1 _3999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_2814_),
    .C(_92_),
    .Y(_273_)
);

AOI21X1 _4000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_270_),
    .C(_268_),
    .Y(_274_)
);

AOI21X1 _4001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_263_),
    .C(_176_),
    .Y(_275_)
);

OAI21X1 _4002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_275_),
    .C(_273_),
    .Y(_277_)
);

NAND3X1 _4003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_277_),
    .C(_131_),
    .Y(_278_)
);

NOR3X1 _4004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_275_),
    .C(_273_),
    .Y(_279_)
);

AOI21X1 _4005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_271_),
    .C(_132_),
    .Y(_280_)
);

OAI21X1 _4006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_279_),
    .B(_280_),
    .C(_130_),
    .Y(_281_)
);

NAND3X1 _4007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_127_),
    .C(_281_),
    .Y(_282_)
);

AOI21X1 _4008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2769_),
    .B(_102_),
    .C(_105_),
    .Y(_283_)
);

OAI21X1 _4009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_275_),
    .C(_132_),
    .Y(_284_)
);

NAND3X1 _4010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_271_),
    .C(_273_),
    .Y(_285_)
);

AOI21X1 _4011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_285_),
    .C(_130_),
    .Y(_286_)
);

AOI21X1 _4012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_272_),
    .C(_131_),
    .Y(_288_)
);

OAI21X1 _4013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_286_),
    .C(_283_),
    .Y(_289_)
);

NAND3X1 _4014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .B(_282_),
    .C(_108_),
    .Y(_290_)
);

NOR3X1 _4015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_109_),
    .C(_114_),
    .Y(_291_)
);

OAI21X1 _4016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_286_),
    .C(_127_),
    .Y(_292_)
);

NAND3X1 _4017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_283_),
    .C(_281_),
    .Y(_293_)
);

NAND3X1 _4018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_293_),
    .C(_291_),
    .Y(_294_)
);

NAND2X1 _4019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_290_),
    .B(_294_),
    .Y(_295_)
);

XNOR2X1 _4020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_295_),
    .Y(_1_[14])
);

NAND3X1 _4021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_289_),
    .C(_291_),
    .Y(_296_)
);

NAND3X1 _4022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_293_),
    .C(_108_),
    .Y(_297_)
);

NAND2X1 _4023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_296_),
    .Y(_298_)
);

OAI21X1 _4024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_298_),
    .C(_296_),
    .Y(_299_)
);

NAND2X1 _4025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_129_),
    .Y(_300_)
);

OAI21X1 _4026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_130_),
    .C(_272_),
    .Y(_301_)
);

NOR2X1 _4027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2523_),
    .B(_220_),
    .Y(_302_)
);

INVX2 _4028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .Y(_303_)
);

NAND3X1 _4029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .B(breg_13_bF$buf3),
    .C(_137_),
    .Y(_304_)
);

OAI21X1 _4030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_136_),
    .C(_304_),
    .Y(_305_)
);

OAI21X1 _4031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_165_),
    .C(_174_),
    .Y(_306_)
);

NAND2X1 _4032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .B(_306_),
    .Y(_308_)
);

OR2X2 _4033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_305_),
    .Y(_309_)
);

NAND3X1 _4034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_308_),
    .C(_309_),
    .Y(_310_)
);

AND2X2 _4035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_305_),
    .Y(_311_)
);

NOR2X1 _4036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .B(_306_),
    .Y(_312_)
);

OAI21X1 _4037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_312_),
    .C(_302_),
    .Y(_313_)
);

NAND2X1 _4038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_310_),
    .Y(_314_)
);

AOI21X1 _4039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_258_),
    .C(_178_),
    .Y(_315_)
);

OAI21X1 _4040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_315_),
    .C(_259_),
    .Y(_316_)
);

AND2X2 _4041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_153_),
    .Y(_317_)
);

NAND2X1 _4042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg[12]),
    .Y(_319_)
);

NAND2X1 _4043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_14_bF$buf2),
    .Y(_320_)
);

NOR2X1 _4044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_320_),
    .Y(_321_)
);

AOI22X1 _4045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_13_bF$buf1),
    .C(breg[1]),
    .D(areg_14_bF$buf1),
    .Y(_322_)
);

NOR2X1 _4046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_321_),
    .Y(_323_)
);

XNOR2X1 _4047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .B(_319_),
    .Y(_324_)
);

AOI21X1 _4048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_148_),
    .C(_150_),
    .Y(_325_)
);

INVX1 _4049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .Y(_326_)
);

AND2X2 _4050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_11_bF$buf2),
    .Y(_327_)
);

NAND2X1 _4051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_15_bF$buf3),
    .Y(_328_)
);

NAND2X1 _4052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_10_bF$buf3),
    .Y(_330_)
);

NOR2X1 _4053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_330_),
    .Y(_331_)
);

INVX1 _4054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_331_),
    .Y(_332_)
);

OAI21X1 _4055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_2614_),
    .C(_328_),
    .Y(_333_)
);

NAND3X1 _4056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_333_),
    .C(_332_),
    .Y(_334_)
);

NAND2X1 _4057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_15_bF$buf2),
    .Y(_335_)
);

OAI21X1 _4058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2330_),
    .B(_335_),
    .C(_333_),
    .Y(_336_)
);

OAI21X1 _4059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_2458_),
    .C(_336_),
    .Y(_337_)
);

NAND3X1 _4060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_337_),
    .C(_326_),
    .Y(_338_)
);

NAND2X1 _4061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_11_bF$buf1),
    .Y(_339_)
);

NOR2X1 _4062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_336_),
    .Y(_341_)
);

AOI21X1 _4063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_332_),
    .C(_327_),
    .Y(_342_)
);

OAI21X1 _4064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_342_),
    .C(_325_),
    .Y(_343_)
);

NAND3X1 _4065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_338_),
    .C(_343_),
    .Y(_344_)
);

OAI21X1 _4066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_322_),
    .C(_319_),
    .Y(_345_)
);

NAND3X1 _4067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg[12]),
    .C(_323_),
    .Y(_346_)
);

NAND2X1 _4068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_346_),
    .Y(_347_)
);

OAI21X1 _4069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_342_),
    .C(_326_),
    .Y(_348_)
);

NAND3X1 _4070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_334_),
    .C(_337_),
    .Y(_349_)
);

NAND3X1 _4071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_347_),
    .B(_349_),
    .C(_348_),
    .Y(_350_)
);

AOI21X1 _4072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_190_),
    .C(_193_),
    .Y(_352_)
);

OAI21X1 _4073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_180_),
    .C(_194_),
    .Y(_353_)
);

NAND3X1 _4074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_344_),
    .C(_350_),
    .Y(_354_)
);

AOI21X1 _4075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_348_),
    .C(_347_),
    .Y(_355_)
);

AOI21X1 _4076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_343_),
    .C(_324_),
    .Y(_356_)
);

NOR3X1 _4077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_192_),
    .C(_196_),
    .Y(_357_)
);

AOI21X1 _4078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_198_),
    .C(_357_),
    .Y(_358_)
);

OAI21X1 _4079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_356_),
    .C(_358_),
    .Y(_359_)
);

NAND3X1 _4080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_354_),
    .C(_359_),
    .Y(_360_)
);

NAND2X1 _4081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_159_),
    .Y(_361_)
);

NAND3X1 _4082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_350_),
    .C(_358_),
    .Y(_363_)
);

OAI21X1 _4083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_356_),
    .C(_353_),
    .Y(_364_)
);

NAND3X1 _4084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_363_),
    .C(_364_),
    .Y(_365_)
);

NAND2X1 _4085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_365_),
    .Y(_366_)
);

AOI21X1 _4086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_241_),
    .C(_206_),
    .Y(_367_)
);

OAI21X1 _4087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_367_),
    .C(_242_),
    .Y(_368_)
);

OAI21X1 _4088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_195_),
    .C(_184_),
    .Y(_369_)
);

INVX2 _4089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .Y(_370_)
);

NOR2X1 _4090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_2342_),
    .Y(_371_)
);

NAND2X1 _4091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf0),
    .B(areg_8_bF$buf3),
    .Y(_372_)
);

OR2X2 _4092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_372_),
    .Y(_374_)
);

OAI21X1 _4093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_2158_),
    .C(_182_),
    .Y(_375_)
);

NAND3X1 _4094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_375_),
    .C(_374_),
    .Y(_376_)
);

OAI21X1 _4095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_372_),
    .C(_375_),
    .Y(_377_)
);

OAI21X1 _4096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_2342_),
    .C(_377_),
    .Y(_378_)
);

NOR2X1 _4097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .B(_208_),
    .Y(_379_)
);

AOI21X1 _4098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_211_),
    .C(_379_),
    .Y(_380_)
);

INVX2 _4099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .Y(_381_)
);

NAND3X1 _4100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_378_),
    .C(_381_),
    .Y(_382_)
);

INVX1 _4101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .Y(_383_)
);

NOR2X1 _4102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_377_),
    .Y(_385_)
);

AOI21X1 _4103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_374_),
    .C(_371_),
    .Y(_386_)
);

OAI21X1 _4104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_386_),
    .C(_380_),
    .Y(_387_)
);

NAND3X1 _4105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_382_),
    .C(_387_),
    .Y(_388_)
);

NAND3X1 _4106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_380_),
    .C(_378_),
    .Y(_389_)
);

OAI21X1 _4107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_386_),
    .C(_381_),
    .Y(_390_)
);

NAND3X1 _4108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_389_),
    .C(_390_),
    .Y(_391_)
);

NAND2X1 _4109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .B(_391_),
    .Y(_392_)
);

OAI21X1 _4110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_240_),
    .C(_228_),
    .Y(_393_)
);

NOR2X1 _4111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_2266_),
    .Y(_394_)
);

NAND2X1 _4112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_11_bF$buf2),
    .Y(_395_)
);

OAI21X1 _4113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_2527_),
    .C(_208_),
    .Y(_396_)
);

OAI21X1 _4114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_395_),
    .C(_396_),
    .Y(_397_)
);

XNOR2X1 _4115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_394_),
    .Y(_398_)
);

OAI21X1 _4116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_215_),
    .C(_219_),
    .Y(_399_)
);

NAND2X1 _4117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_12_bF$buf2),
    .Y(_400_)
);

INVX2 _4118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .Y(_401_)
);

NAND2X1 _4119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_15_bF$buf3),
    .Y(_402_)
);

OR2X2 _4120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_402_),
    .Y(_403_)
);

AOI22X1 _4121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg_15_bF$buf2),
    .C(areg_2_bF$buf3),
    .D(breg_13_bF$buf2),
    .Y(_404_)
);

INVX2 _4122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .Y(_407_)
);

NAND3X1 _4123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_407_),
    .C(_403_),
    .Y(_408_)
);

NOR2X1 _4124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_402_),
    .Y(_409_)
);

OAI21X1 _4125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_404_),
    .C(_400_),
    .Y(_410_)
);

NAND3X1 _4126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_399_),
    .C(_408_),
    .Y(_411_)
);

AOI21X1 _4127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_216_),
    .B(_222_),
    .C(_225_),
    .Y(_412_)
);

NOR3X1 _4128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_404_),
    .C(_409_),
    .Y(_413_)
);

AOI21X1 _4129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .B(_403_),
    .C(_401_),
    .Y(_414_)
);

OAI21X1 _4130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_413_),
    .C(_412_),
    .Y(_415_)
);

NAND3X1 _4131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_411_),
    .B(_415_),
    .C(_398_),
    .Y(_416_)
);

INVX1 _4132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .Y(_418_)
);

XNOR2X1 _4133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_397_),
    .B(_418_),
    .Y(_419_)
);

OAI21X1 _4134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_413_),
    .C(_399_),
    .Y(_420_)
);

NAND3X1 _4135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_412_),
    .B(_410_),
    .C(_408_),
    .Y(_421_)
);

NAND3X1 _4136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_420_),
    .C(_419_),
    .Y(_422_)
);

NAND3X1 _4137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_422_),
    .C(_393_),
    .Y(_423_)
);

AOI21X1 _4138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_213_),
    .C(_239_),
    .Y(_424_)
);

AOI21X1 _4139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_420_),
    .C(_419_),
    .Y(_425_)
);

AOI21X1 _4140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_411_),
    .B(_415_),
    .C(_398_),
    .Y(_426_)
);

OAI21X1 _4141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_426_),
    .C(_424_),
    .Y(_427_)
);

NAND3X1 _4142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_427_),
    .C(_392_),
    .Y(_429_)
);

NAND3X1 _4143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_382_),
    .C(_387_),
    .Y(_430_)
);

NAND3X1 _4144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_389_),
    .C(_390_),
    .Y(_431_)
);

NAND2X1 _4145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_431_),
    .Y(_432_)
);

NOR3X1 _4146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_426_),
    .C(_424_),
    .Y(_433_)
);

AOI21X1 _4147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_422_),
    .C(_393_),
    .Y(_434_)
);

OAI21X1 _4148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_434_),
    .C(_432_),
    .Y(_435_)
);

NAND3X1 _4149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_368_),
    .C(_435_),
    .Y(_436_)
);

NOR3X1 _4150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_249_),
    .C(_245_),
    .Y(_437_)
);

AOI21X1 _4151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_204_),
    .C(_437_),
    .Y(_438_)
);

OAI21X1 _4152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_426_),
    .C(_393_),
    .Y(_440_)
);

NAND3X1 _4153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_422_),
    .C(_424_),
    .Y(_441_)
);

AOI21X1 _4154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_440_),
    .C(_432_),
    .Y(_442_)
);

AOI21X1 _4155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_427_),
    .C(_392_),
    .Y(_443_)
);

OAI21X1 _4156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_443_),
    .C(_438_),
    .Y(_444_)
);

NAND3X1 _4157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_436_),
    .C(_366_),
    .Y(_445_)
);

NAND3X1 _4158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_354_),
    .C(_359_),
    .Y(_446_)
);

NAND3X1 _4159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_363_),
    .C(_364_),
    .Y(_447_)
);

NAND2X1 _4160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_447_),
    .Y(_448_)
);

NOR3X1 _4161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_443_),
    .C(_438_),
    .Y(_449_)
);

AOI21X1 _4162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_435_),
    .C(_368_),
    .Y(_451_)
);

OAI21X1 _4163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_449_),
    .B(_451_),
    .C(_448_),
    .Y(_452_)
);

NAND3X1 _4164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_316_),
    .B(_445_),
    .C(_452_),
    .Y(_453_)
);

NOR3X1 _4165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_261_),
    .B(_262_),
    .C(_260_),
    .Y(_454_)
);

AOI21X1 _4166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_263_),
    .C(_454_),
    .Y(_455_)
);

OAI21X1 _4167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_442_),
    .B(_443_),
    .C(_368_),
    .Y(_456_)
);

NAND3X1 _4168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_438_),
    .C(_435_),
    .Y(_457_)
);

AOI21X1 _4169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_457_),
    .C(_448_),
    .Y(_458_)
);

AOI21X1 _4170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_436_),
    .C(_366_),
    .Y(_459_)
);

OAI21X1 _4171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_459_),
    .C(_455_),
    .Y(_460_)
);

NAND3X1 _4172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_460_),
    .C(_453_),
    .Y(_462_)
);

NAND3X1 _4173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_308_),
    .C(_309_),
    .Y(_463_)
);

OAI21X1 _4174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_312_),
    .C(_303_),
    .Y(_464_)
);

NAND2X1 _4175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_463_),
    .Y(_465_)
);

OAI21X1 _4176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_459_),
    .C(_316_),
    .Y(_466_)
);

NAND3X1 _4177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .B(_445_),
    .C(_452_),
    .Y(_467_)
);

NAND3X1 _4178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .B(_466_),
    .C(_467_),
    .Y(_468_)
);

NAND3X1 _4179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_301_),
    .B(_462_),
    .C(_468_),
    .Y(_469_)
);

AOI21X1 _4180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_131_),
    .C(_279_),
    .Y(_470_)
);

AOI21X1 _4181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_466_),
    .B(_467_),
    .C(_465_),
    .Y(_471_)
);

AOI21X1 _4182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_453_),
    .C(_314_),
    .Y(_473_)
);

OAI21X1 _4183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(_473_),
    .C(_470_),
    .Y(_474_)
);

NAND3X1 _4184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_469_),
    .C(_474_),
    .Y(_475_)
);

INVX2 _4185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .Y(_476_)
);

OAI21X1 _4186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(_473_),
    .C(_301_),
    .Y(_477_)
);

NAND3X1 _4187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_468_),
    .C(_470_),
    .Y(_478_)
);

NAND3X1 _4188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_478_),
    .C(_477_),
    .Y(_479_)
);

AOI21X1 _4189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_475_),
    .B(_479_),
    .C(_282_),
    .Y(_480_)
);

INVX1 _4190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .Y(_481_)
);

NAND3X1 _4191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_469_),
    .C(_474_),
    .Y(_482_)
);

NAND3X1 _4192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .B(_478_),
    .C(_477_),
    .Y(_484_)
);

AOI21X1 _4193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_484_),
    .C(_481_),
    .Y(_485_)
);

NOR2X1 _4194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_485_),
    .Y(_486_)
);

XOR2X1 _4195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_486_),
    .Y(_1_[15])
);

NAND3X1 _4196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_481_),
    .B(_482_),
    .C(_484_),
    .Y(_487_)
);

NAND3X1 _4197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_475_),
    .C(_479_),
    .Y(_488_)
);

NAND3X1 _4198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_295_),
    .C(_488_),
    .Y(_489_)
);

INVX1 _4199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .Y(_490_)
);

AOI21X1 _4200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_490_),
    .B(_488_),
    .C(_480_),
    .Y(_491_)
);

OAI21X1 _4201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_123_),
    .C(_491_),
    .Y(_492_)
);

AND2X2 _4202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2754_),
    .B(_2757_),
    .Y(_494_)
);

AND2X2 _4203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_119_),
    .Y(_495_)
);

NAND2X1 _4204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_494_),
    .B(_495_),
    .Y(_496_)
);

NOR2X1 _4205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_489_),
    .Y(_497_)
);

AOI21X1 _4206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(_497_),
    .C(_492_),
    .Y(_498_)
);

AOI21X1 _4207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_468_),
    .C(_301_),
    .Y(_499_)
);

OAI21X1 _4208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_499_),
    .B(_300_),
    .C(_469_),
    .Y(_500_)
);

OAI21X1 _4209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_312_),
    .B(_303_),
    .C(_308_),
    .Y(_501_)
);

INVX2 _4210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .Y(_502_)
);

AOI21X1 _4211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_452_),
    .C(_316_),
    .Y(_503_)
);

OAI21X1 _4212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_465_),
    .C(_453_),
    .Y(_505_)
);

OAI21X1 _4213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_320_),
    .C(_346_),
    .Y(_506_)
);

NAND2X1 _4214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_446_),
    .Y(_507_)
);

XOR2X1 _4215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .B(_506_),
    .Y(_508_)
);

INVX2 _4216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .Y(_509_)
);

OAI21X1 _4217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .B(_448_),
    .C(_436_),
    .Y(_510_)
);

NAND2X1 _4218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_344_),
    .Y(_511_)
);

NAND2X1 _4219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .B(breg_15_bF$buf1),
    .Y(_512_)
);

NAND2X1 _4220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_13_bF$buf0),
    .Y(_513_)
);

NOR2X1 _4221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_513_),
    .Y(_514_)
);

AOI22X1 _4222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_13_bF$buf3),
    .C(breg_4_bF$buf3),
    .D(areg[12]),
    .Y(_516_)
);

OAI21X1 _4223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_516_),
    .C(_512_),
    .Y(_517_)
);

INVX1 _4224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .Y(_518_)
);

NOR2X1 _4225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_514_),
    .Y(_519_)
);

NAND2X1 _4226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_519_),
    .Y(_520_)
);

AND2X2 _4227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_517_),
    .Y(_521_)
);

AOI21X1 _4228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_327_),
    .B(_333_),
    .C(_331_),
    .Y(_522_)
);

INVX1 _4229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .Y(_523_)
);

INVX1 _4230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .Y(_524_)
);

NOR2X1 _4231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_335_),
    .Y(_525_)
);

INVX1 _4232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .Y(_527_)
);

INVX4 _4233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf1),
    .Y(_528_)
);

NAND2X1 _4234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg_11_bF$buf0),
    .Y(_529_)
);

OAI21X1 _4235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2534_),
    .B(_528_),
    .C(_529_),
    .Y(_530_)
);

NAND3X1 _4236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_530_),
    .C(_527_),
    .Y(_531_)
);

AOI22X1 _4237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_15_bF$buf0),
    .C(breg_5_bF$buf0),
    .D(areg_11_bF$buf3),
    .Y(_532_)
);

OAI21X1 _4238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_525_),
    .B(_532_),
    .C(_320_),
    .Y(_533_)
);

NAND3X1 _4239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_531_),
    .C(_523_),
    .Y(_534_)
);

OAI21X1 _4240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_335_),
    .C(_530_),
    .Y(_535_)
);

NOR2X1 _4241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_535_),
    .Y(_536_)
);

INVX1 _4242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .Y(_538_)
);

OAI21X1 _4243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_538_),
    .C(_522_),
    .Y(_539_)
);

NAND3X1 _4244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_521_),
    .C(_539_),
    .Y(_540_)
);

NAND2X1 _4245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_517_),
    .B(_520_),
    .Y(_541_)
);

OAI21X1 _4246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_538_),
    .C(_523_),
    .Y(_542_)
);

NAND3X1 _4247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_533_),
    .C(_531_),
    .Y(_543_)
);

NAND3X1 _4248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_543_),
    .C(_542_),
    .Y(_544_)
);

AOI21X1 _4249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_378_),
    .C(_381_),
    .Y(_545_)
);

OAI21X1 _4250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_370_),
    .C(_382_),
    .Y(_546_)
);

NAND3X1 _4251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_544_),
    .C(_540_),
    .Y(_547_)
);

AOI21X1 _4252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_542_),
    .C(_541_),
    .Y(_549_)
);

AOI21X1 _4253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_539_),
    .C(_521_),
    .Y(_550_)
);

NOR3X1 _4254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_380_),
    .C(_385_),
    .Y(_551_)
);

AOI21X1 _4255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_387_),
    .C(_551_),
    .Y(_552_)
);

OAI21X1 _4256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_550_),
    .C(_552_),
    .Y(_553_)
);

NAND3X1 _4257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(_547_),
    .C(_553_),
    .Y(_554_)
);

AND2X2 _4258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_338_),
    .Y(_555_)
);

NAND3X1 _4259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .B(_540_),
    .C(_552_),
    .Y(_556_)
);

OAI21X1 _4260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_550_),
    .C(_546_),
    .Y(_557_)
);

NAND3X1 _4261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_556_),
    .C(_557_),
    .Y(_558_)
);

NAND2X1 _4262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_558_),
    .Y(_560_)
);

OAI21X1 _4263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_432_),
    .B(_434_),
    .C(_423_),
    .Y(_561_)
);

OAI21X1 _4264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_383_),
    .C(_374_),
    .Y(_562_)
);

NAND2X1 _4265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_10_bF$buf2),
    .Y(_563_)
);

INVX1 _4266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .Y(_564_)
);

NAND2X1 _4267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf3),
    .B(areg[9]),
    .Y(_565_)
);

NOR2X1 _4268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_182_),
    .B(_565_),
    .Y(_566_)
);

INVX1 _4269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .Y(_567_)
);

AOI22X1 _4270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf1),
    .B(areg[9]),
    .C(breg_8_bF$buf2),
    .D(areg_8_bF$buf2),
    .Y(_568_)
);

INVX1 _4271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .Y(_569_)
);

NAND3X1 _4272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(_569_),
    .C(_567_),
    .Y(_571_)
);

OAI21X1 _4273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_566_),
    .B(_568_),
    .C(_563_),
    .Y(_572_)
);

NOR2X1 _4274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_395_),
    .Y(_573_)
);

AOI21X1 _4275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_396_),
    .C(_573_),
    .Y(_574_)
);

INVX2 _4276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .Y(_575_)
);

NAND3X1 _4277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_571_),
    .C(_575_),
    .Y(_576_)
);

NOR3X1 _4278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_568_),
    .C(_566_),
    .Y(_577_)
);

INVX2 _4279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .Y(_578_)
);

OAI21X1 _4280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_577_),
    .C(_574_),
    .Y(_579_)
);

NAND3X1 _4281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_576_),
    .C(_579_),
    .Y(_580_)
);

INVX2 _4282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .Y(_582_)
);

NAND3X1 _4283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_574_),
    .C(_571_),
    .Y(_583_)
);

OAI21X1 _4284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_578_),
    .B(_577_),
    .C(_575_),
    .Y(_584_)
);

NAND3X1 _4285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_583_),
    .C(_584_),
    .Y(_585_)
);

NAND2X1 _4286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(_585_),
    .Y(_586_)
);

AOI21X1 _4287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_408_),
    .C(_399_),
    .Y(_587_)
);

OAI21X1 _4288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_587_),
    .C(_411_),
    .Y(_588_)
);

NAND2X1 _4289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_9_bF$buf3),
    .Y(_589_)
);

INVX1 _4290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .Y(_590_)
);

AND2X2 _4291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_10_bF$buf0),
    .Y(_591_)
);

AND2X2 _4292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_11_bF$buf1),
    .Y(_592_)
);

AOI22X1 _4293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_11_bF$buf0),
    .C(areg[6]),
    .D(breg_10_bF$buf3),
    .Y(_593_)
);

AOI21X1 _4294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_591_),
    .B(_592_),
    .C(_593_),
    .Y(_594_)
);

XNOR2X1 _4295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_590_),
    .Y(_595_)
);

OAI21X1 _4296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_404_),
    .C(_403_),
    .Y(_596_)
);

NAND2X1 _4297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_12_bF$buf1),
    .Y(_597_)
);

NAND2X1 _4298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_14_bF$buf3),
    .Y(_598_)
);

NOR2X1 _4299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_598_),
    .Y(_599_)
);

AOI22X1 _4300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_14_bF$buf2),
    .C(areg_3_bF$buf2),
    .D(breg_13_bF$buf1),
    .Y(_600_)
);

NOR3X1 _4301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(_600_),
    .C(_599_),
    .Y(_601_)
);

INVX2 _4302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .Y(_603_)
);

AND2X2 _4303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_14_bF$buf1),
    .Y(_604_)
);

NAND2X1 _4304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_604_),
    .Y(_605_)
);

INVX2 _4305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_600_),
    .Y(_606_)
);

AOI21X1 _4306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_606_),
    .B(_605_),
    .C(_603_),
    .Y(_607_)
);

OAI21X1 _4307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_601_),
    .C(_596_),
    .Y(_608_)
);

AOI21X1 _4308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_407_),
    .C(_409_),
    .Y(_609_)
);

NAND3X1 _4309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_606_),
    .C(_605_),
    .Y(_610_)
);

OAI21X1 _4310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_600_),
    .C(_597_),
    .Y(_611_)
);

NAND3X1 _4311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_609_),
    .C(_610_),
    .Y(_612_)
);

AOI21X1 _4312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_612_),
    .B(_608_),
    .C(_595_),
    .Y(_615_)
);

XNOR2X1 _4313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_589_),
    .Y(_616_)
);

NAND3X1 _4314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_596_),
    .C(_610_),
    .Y(_617_)
);

OAI21X1 _4315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_601_),
    .C(_609_),
    .Y(_618_)
);

AOI21X1 _4316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_618_),
    .C(_616_),
    .Y(_619_)
);

OAI21X1 _4317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_619_),
    .C(_588_),
    .Y(_620_)
);

NOR3X1 _4318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_412_),
    .C(_414_),
    .Y(_621_)
);

AOI21X1 _4319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_398_),
    .C(_621_),
    .Y(_622_)
);

NAND3X1 _4320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_616_),
    .B(_617_),
    .C(_618_),
    .Y(_623_)
);

NAND3X1 _4321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .B(_612_),
    .C(_608_),
    .Y(_624_)
);

NAND3X1 _4322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_623_),
    .C(_622_),
    .Y(_626_)
);

AOI21X1 _4323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_620_),
    .C(_586_),
    .Y(_627_)
);

NAND3X1 _4324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_576_),
    .C(_579_),
    .Y(_628_)
);

NAND3X1 _4325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_583_),
    .C(_584_),
    .Y(_629_)
);

NAND2X1 _4326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_629_),
    .Y(_630_)
);

NAND3X1 _4327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_623_),
    .C(_588_),
    .Y(_631_)
);

OAI21X1 _4328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_619_),
    .C(_622_),
    .Y(_632_)
);

AOI21X1 _4329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_632_),
    .C(_630_),
    .Y(_633_)
);

OAI21X1 _4330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_633_),
    .C(_561_),
    .Y(_634_)
);

AOI21X1 _4331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_392_),
    .C(_433_),
    .Y(_635_)
);

NAND3X1 _4332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_632_),
    .C(_630_),
    .Y(_637_)
);

NAND3X1 _4333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_626_),
    .C(_586_),
    .Y(_638_)
);

NAND3X1 _4334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_638_),
    .C(_635_),
    .Y(_639_)
);

AOI21X1 _4335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_639_),
    .C(_560_),
    .Y(_640_)
);

NAND3X1 _4336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_547_),
    .C(_553_),
    .Y(_641_)
);

NAND3X1 _4337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_511_),
    .B(_556_),
    .C(_557_),
    .Y(_642_)
);

NAND2X1 _4338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_642_),
    .Y(_643_)
);

NAND3X1 _4339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_638_),
    .C(_561_),
    .Y(_644_)
);

OAI21X1 _4340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_633_),
    .C(_635_),
    .Y(_645_)
);

AOI21X1 _4341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_644_),
    .C(_643_),
    .Y(_646_)
);

OAI21X1 _4342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_646_),
    .C(_510_),
    .Y(_648_)
);

AOI21X1 _4343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_366_),
    .C(_449_),
    .Y(_649_)
);

NAND3X1 _4344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_644_),
    .B(_645_),
    .C(_643_),
    .Y(_650_)
);

NOR3X1 _4345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_633_),
    .C(_635_),
    .Y(_651_)
);

AOI21X1 _4346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_638_),
    .C(_561_),
    .Y(_652_)
);

OAI21X1 _4347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(_652_),
    .C(_560_),
    .Y(_653_)
);

NAND3X1 _4348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_649_),
    .C(_653_),
    .Y(_654_)
);

AOI21X1 _4349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_654_),
    .C(_509_),
    .Y(_655_)
);

NAND3X1 _4350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_510_),
    .C(_653_),
    .Y(_656_)
);

OAI21X1 _4351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_646_),
    .C(_649_),
    .Y(_657_)
);

AOI21X1 _4352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_657_),
    .B(_656_),
    .C(_508_),
    .Y(_659_)
);

OAI21X1 _4353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_655_),
    .C(_505_),
    .Y(_660_)
);

NOR3X1 _4354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_459_),
    .C(_455_),
    .Y(_661_)
);

AOI21X1 _4355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_314_),
    .B(_460_),
    .C(_661_),
    .Y(_662_)
);

NAND3X1 _4356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_657_),
    .C(_656_),
    .Y(_663_)
);

NOR3X1 _4357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_646_),
    .C(_649_),
    .Y(_664_)
);

AOI21X1 _4358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_650_),
    .B(_653_),
    .C(_510_),
    .Y(_665_)
);

OAI21X1 _4359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_665_),
    .C(_509_),
    .Y(_666_)
);

NAND3X1 _4360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_662_),
    .C(_666_),
    .Y(_667_)
);

AOI21X1 _4361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_667_),
    .C(_502_),
    .Y(_668_)
);

NAND3X1 _4362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_505_),
    .C(_666_),
    .Y(_670_)
);

OAI21X1 _4363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_655_),
    .C(_662_),
    .Y(_671_)
);

AOI21X1 _4364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_670_),
    .C(_501_),
    .Y(_672_)
);

OAI21X1 _4365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(_672_),
    .C(_500_),
    .Y(_673_)
);

NOR3X1 _4366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_471_),
    .B(_473_),
    .C(_470_),
    .Y(_674_)
);

AOI21X1 _4367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_476_),
    .B(_474_),
    .C(_674_),
    .Y(_675_)
);

NAND3X1 _4368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_671_),
    .C(_670_),
    .Y(_676_)
);

NAND3X1 _4369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_660_),
    .C(_667_),
    .Y(_677_)
);

NAND3X1 _4370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_677_),
    .C(_675_),
    .Y(_678_)
);

AND2X2 _4371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_678_),
    .Y(_679_)
);

XOR2X1 _4372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_679_),
    .Y(_1_[16])
);

NAND3X1 _4373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .B(_676_),
    .C(_677_),
    .Y(_681_)
);

OAI21X1 _4374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_679_),
    .C(_681_),
    .Y(_682_)
);

AOI21X1 _4375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_666_),
    .C(_505_),
    .Y(_683_)
);

OAI21X1 _4376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_502_),
    .C(_670_),
    .Y(_684_)
);

NAND2X1 _4377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_507_),
    .Y(_685_)
);

INVX2 _4378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .Y(_686_)
);

OAI21X1 _4379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .B(_665_),
    .C(_656_),
    .Y(_687_)
);

OAI21X1 _4380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_513_),
    .C(_520_),
    .Y(_688_)
);

NAND2X1 _4381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_554_),
    .Y(_689_)
);

XOR2X1 _4382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_688_),
    .Y(_691_)
);

OAI21X1 _4383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_652_),
    .C(_644_),
    .Y(_692_)
);

AND2X2 _4384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_540_),
    .B(_534_),
    .Y(_693_)
);

AOI22X1 _4385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_13_bF$buf2),
    .C(breg_5_bF$buf3),
    .D(areg[12]),
    .Y(_694_)
);

NAND2X1 _4386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg[12]),
    .Y(_695_)
);

NAND2X1 _4387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_13_bF$buf1),
    .Y(_696_)
);

NOR2X1 _4388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_696_),
    .Y(_697_)
);

NOR2X1 _4389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_694_),
    .B(_697_),
    .Y(_698_)
);

OAI21X1 _4390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_532_),
    .B(_320_),
    .C(_527_),
    .Y(_699_)
);

NAND2X1 _4391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .B(areg_14_bF$buf0),
    .Y(_700_)
);

INVX2 _4392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .Y(_702_)
);

NAND2X1 _4393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_11_bF$buf2),
    .Y(_703_)
);

NAND2X1 _4394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_15_bF$buf3),
    .Y(_704_)
);

OR2X2 _4395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_704_),
    .Y(_705_)
);

OAI21X1 _4396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_528_),
    .C(_703_),
    .Y(_706_)
);

NAND3X1 _4397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_706_),
    .C(_705_),
    .Y(_707_)
);

NAND2X1 _4398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_15_bF$buf2),
    .Y(_708_)
);

NOR2X1 _4399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2617_),
    .B(_708_),
    .Y(_709_)
);

AND2X2 _4400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_704_),
    .Y(_710_)
);

OAI21X1 _4401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_709_),
    .C(_700_),
    .Y(_711_)
);

NAND3X1 _4402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_711_),
    .C(_699_),
    .Y(_713_)
);

AOI21X1 _4403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_530_),
    .C(_525_),
    .Y(_714_)
);

NOR3X1 _4404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_709_),
    .C(_710_),
    .Y(_715_)
);

AOI21X1 _4405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .B(_705_),
    .C(_702_),
    .Y(_716_)
);

OAI21X1 _4406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_716_),
    .C(_714_),
    .Y(_717_)
);

NAND3X1 _4407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .B(_717_),
    .C(_713_),
    .Y(_718_)
);

INVX1 _4408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_698_),
    .Y(_719_)
);

OAI21X1 _4409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_716_),
    .C(_699_),
    .Y(_720_)
);

NAND3X1 _4410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_711_),
    .C(_707_),
    .Y(_721_)
);

NAND3X1 _4411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_721_),
    .C(_720_),
    .Y(_722_)
);

AOI21X1 _4412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_571_),
    .C(_575_),
    .Y(_724_)
);

OAI21X1 _4413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_582_),
    .C(_576_),
    .Y(_725_)
);

NAND3X1 _4414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_722_),
    .C(_725_),
    .Y(_726_)
);

AOI21X1 _4415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_720_),
    .C(_719_),
    .Y(_727_)
);

AOI21X1 _4416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_717_),
    .B(_713_),
    .C(_698_),
    .Y(_728_)
);

NOR3X1 _4417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_574_),
    .C(_578_),
    .Y(_729_)
);

AOI21X1 _4418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_579_),
    .C(_729_),
    .Y(_730_)
);

OAI21X1 _4419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(_728_),
    .C(_730_),
    .Y(_731_)
);

NAND3X1 _4420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_731_),
    .C(_693_),
    .Y(_732_)
);

NAND2X1 _4421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_540_),
    .Y(_733_)
);

NAND3X1 _4422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_722_),
    .C(_730_),
    .Y(_735_)
);

OAI21X1 _4423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .B(_727_),
    .C(_725_),
    .Y(_736_)
);

NAND3X1 _4424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_736_),
    .C(_735_),
    .Y(_737_)
);

NAND2X1 _4425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_737_),
    .B(_732_),
    .Y(_738_)
);

AOI21X1 _4426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_623_),
    .C(_588_),
    .Y(_739_)
);

OAI21X1 _4427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_739_),
    .C(_631_),
    .Y(_740_)
);

OAI21X1 _4428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_568_),
    .C(_567_),
    .Y(_741_)
);

NAND2X1 _4429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_10_bF$buf1),
    .Y(_742_)
);

INVX1 _4430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .Y(_743_)
);

AND2X2 _4431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf1),
    .B(areg[9]),
    .Y(_744_)
);

AND2X2 _4432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf1),
    .B(breg_9_bF$buf2),
    .Y(_746_)
);

NAND2X1 _4433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_746_),
    .Y(_747_)
);

OAI21X1 _4434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_2266_),
    .C(_565_),
    .Y(_748_)
);

NAND3X1 _4435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_748_),
    .C(_747_),
    .Y(_749_)
);

OAI21X1 _4436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .B(_2342_),
    .C(_746_),
    .Y(_750_)
);

OAI21X1 _4437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_2266_),
    .C(_744_),
    .Y(_751_)
);

NAND3X1 _4438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_750_),
    .C(_751_),
    .Y(_752_)
);

NAND2X1 _4439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_11_bF$buf3),
    .Y(_753_)
);

OAI22X1 _4440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_753_),
    .C(_593_),
    .D(_589_),
    .Y(_754_)
);

NAND3X1 _4441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_749_),
    .C(_752_),
    .Y(_755_)
);

AOI21X1 _4442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_751_),
    .C(_742_),
    .Y(_757_)
);

AOI21X1 _4443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_748_),
    .B(_747_),
    .C(_743_),
    .Y(_758_)
);

INVX1 _4444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .Y(_759_)
);

OAI21X1 _4445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .B(_758_),
    .C(_759_),
    .Y(_760_)
);

NAND3X1 _4446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .B(_755_),
    .C(_760_),
    .Y(_761_)
);

INVX1 _4447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .Y(_762_)
);

NAND3X1 _4448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(_759_),
    .C(_752_),
    .Y(_763_)
);

OAI21X1 _4449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .B(_758_),
    .C(_754_),
    .Y(_764_)
);

NAND3X1 _4450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_763_),
    .B(_762_),
    .C(_764_),
    .Y(_765_)
);

AND2X2 _4451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_761_),
    .Y(_766_)
);

AOI21X1 _4452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_610_),
    .C(_596_),
    .Y(_768_)
);

OAI21X1 _4453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_595_),
    .C(_617_),
    .Y(_769_)
);

NAND2X1 _4454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf1),
    .B(breg_10_bF$buf2),
    .Y(_770_)
);

AND2X2 _4455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_11_bF$buf2),
    .Y(_771_)
);

AND2X2 _4456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_12_bF$buf0),
    .Y(_772_)
);

AOI22X1 _4457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_12_bF$buf3),
    .C(areg[6]),
    .D(breg_11_bF$buf1),
    .Y(_773_)
);

AOI21X1 _4458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_772_),
    .C(_773_),
    .Y(_774_)
);

XNOR2X1 _4459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_770_),
    .Y(_775_)
);

OAI21X1 _4460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(_600_),
    .C(_605_),
    .Y(_776_)
);

NAND2X1 _4461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_13_bF$buf0),
    .Y(_777_)
);

INVX2 _4462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .Y(_779_)
);

AND2X2 _4463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_15_bF$buf0),
    .Y(_780_)
);

NAND2X1 _4464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_604_),
    .Y(_781_)
);

AOI22X1 _4465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_15_bF$buf3),
    .C(areg_3_bF$buf0),
    .D(breg_14_bF$buf0),
    .Y(_782_)
);

INVX2 _4466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_782_),
    .Y(_783_)
);

NAND3X1 _4467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_783_),
    .C(_781_),
    .Y(_784_)
);

NOR2X1 _4468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_598_),
    .Y(_785_)
);

OAI21X1 _4469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_785_),
    .B(_782_),
    .C(_777_),
    .Y(_786_)
);

NAND3X1 _4470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .B(_786_),
    .C(_784_),
    .Y(_787_)
);

AOI21X1 _4471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_606_),
    .C(_599_),
    .Y(_788_)
);

NOR3X1 _4472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_782_),
    .C(_785_),
    .Y(_790_)
);

AOI21X1 _4473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_781_),
    .C(_779_),
    .Y(_791_)
);

OAI21X1 _4474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_790_),
    .C(_788_),
    .Y(_792_)
);

NAND3X1 _4475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_787_),
    .C(_792_),
    .Y(_793_)
);

INVX2 _4476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_770_),
    .Y(_794_)
);

XNOR2X1 _4477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_794_),
    .Y(_795_)
);

OAI21X1 _4478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_790_),
    .C(_776_),
    .Y(_796_)
);

NAND3X1 _4479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_788_),
    .C(_784_),
    .Y(_797_)
);

NAND3X1 _4480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_797_),
    .C(_796_),
    .Y(_798_)
);

NAND3X1 _4481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_793_),
    .C(_798_),
    .Y(_799_)
);

NOR3X1 _4482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_601_),
    .B(_609_),
    .C(_607_),
    .Y(_801_)
);

AOI21X1 _4483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_616_),
    .C(_801_),
    .Y(_802_)
);

AOI21X1 _4484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_797_),
    .B(_796_),
    .C(_795_),
    .Y(_803_)
);

AOI21X1 _4485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_787_),
    .B(_792_),
    .C(_775_),
    .Y(_804_)
);

OAI21X1 _4486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_804_),
    .C(_802_),
    .Y(_805_)
);

NAND3X1 _4487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_766_),
    .C(_805_),
    .Y(_806_)
);

NAND2X1 _4488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_761_),
    .B(_765_),
    .Y(_807_)
);

OAI21X1 _4489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_804_),
    .C(_769_),
    .Y(_808_)
);

NAND3X1 _4490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .B(_798_),
    .C(_802_),
    .Y(_809_)
);

NAND3X1 _4491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_807_),
    .B(_809_),
    .C(_808_),
    .Y(_810_)
);

NAND3X1 _4492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_810_),
    .C(_740_),
    .Y(_811_)
);

NOR3X1 _4493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_619_),
    .C(_622_),
    .Y(_812_)
);

AOI21X1 _4494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_630_),
    .C(_812_),
    .Y(_813_)
);

AOI21X1 _4495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_808_),
    .C(_807_),
    .Y(_814_)
);

AOI21X1 _4496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_805_),
    .C(_766_),
    .Y(_815_)
);

OAI21X1 _4497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_815_),
    .C(_813_),
    .Y(_816_)
);

NAND3X1 _4498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_816_),
    .C(_738_),
    .Y(_817_)
);

NAND3X1 _4499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_731_),
    .C(_726_),
    .Y(_818_)
);

NAND3X1 _4500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_735_),
    .C(_693_),
    .Y(_819_)
);

NAND2X1 _4501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_819_),
    .Y(_820_)
);

NOR3X1 _4502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_815_),
    .C(_813_),
    .Y(_822_)
);

AOI21X1 _4503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_810_),
    .C(_740_),
    .Y(_823_)
);

OAI21X1 _4504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_822_),
    .B(_823_),
    .C(_820_),
    .Y(_824_)
);

NAND3X1 _4505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .B(_692_),
    .C(_824_),
    .Y(_825_)
);

AOI21X1 _4506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_645_),
    .B(_643_),
    .C(_651_),
    .Y(_826_)
);

OAI21X1 _4507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_815_),
    .C(_740_),
    .Y(_827_)
);

NAND3X1 _4508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_810_),
    .C(_813_),
    .Y(_828_)
);

AOI21X1 _4509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_827_),
    .C(_820_),
    .Y(_829_)
);

AOI21X1 _4510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_816_),
    .C(_738_),
    .Y(_830_)
);

OAI21X1 _4511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(_830_),
    .C(_826_),
    .Y(_831_)
);

NAND3X1 _4512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_831_),
    .C(_825_),
    .Y(_833_)
);

INVX2 _4513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .Y(_834_)
);

NOR3X1 _4514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(_830_),
    .C(_826_),
    .Y(_835_)
);

AOI21X1 _4515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .B(_824_),
    .C(_692_),
    .Y(_836_)
);

OAI21X1 _4516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_836_),
    .C(_834_),
    .Y(_837_)
);

NAND3X1 _4517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_687_),
    .C(_837_),
    .Y(_838_)
);

AOI21X1 _4518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_657_),
    .C(_664_),
    .Y(_839_)
);

OAI21X1 _4519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(_830_),
    .C(_692_),
    .Y(_840_)
);

NAND3X1 _4520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_817_),
    .B(_826_),
    .C(_824_),
    .Y(_841_)
);

AOI21X1 _4521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_841_),
    .C(_834_),
    .Y(_842_)
);

AOI21X1 _4522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_825_),
    .C(_691_),
    .Y(_844_)
);

OAI21X1 _4523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_844_),
    .C(_839_),
    .Y(_845_)
);

NAND3X1 _4524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_845_),
    .C(_838_),
    .Y(_846_)
);

NOR3X1 _4525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_844_),
    .C(_839_),
    .Y(_847_)
);

AOI21X1 _4526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_837_),
    .C(_687_),
    .Y(_848_)
);

OAI21X1 _4527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_848_),
    .C(_685_),
    .Y(_849_)
);

NAND3X1 _4528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_684_),
    .C(_849_),
    .Y(_850_)
);

AOI21X1 _4529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_849_),
    .C(_684_),
    .Y(_851_)
);

INVX1 _4530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .Y(_852_)
);

NAND2X1 _4531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .B(_852_),
    .Y(_853_)
);

XNOR2X1 _4532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_853_),
    .Y(_1_[17])
);

AOI21X1 _4533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_850_),
    .C(_851_),
    .Y(_854_)
);

INVX1 _4534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_854_),
    .Y(_855_)
);

OAI21X1 _4535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_844_),
    .C(_687_),
    .Y(_856_)
);

NAND3X1 _4536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_833_),
    .C(_837_),
    .Y(_857_)
);

AOI21X1 _4537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_856_),
    .B(_857_),
    .C(_685_),
    .Y(_858_)
);

AOI21X1 _4538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_845_),
    .B(_838_),
    .C(_686_),
    .Y(_859_)
);

OAI21X1 _4539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_858_),
    .C(_684_),
    .Y(_860_)
);

NOR3X1 _4540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_659_),
    .B(_655_),
    .C(_662_),
    .Y(_861_)
);

AOI21X1 _4541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_671_),
    .C(_861_),
    .Y(_862_)
);

NAND3X1 _4542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_846_),
    .B(_862_),
    .C(_849_),
    .Y(_865_)
);

AOI22X1 _4543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_678_),
    .C(_860_),
    .D(_865_),
    .Y(_866_)
);

INVX1 _4544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .Y(_867_)
);

OAI21X1 _4545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_867_),
    .C(_855_),
    .Y(_868_)
);

OAI21X1 _4546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_848_),
    .B(_685_),
    .C(_838_),
    .Y(_869_)
);

NAND2X1 _4547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(_689_),
    .Y(_870_)
);

OAI21X1 _4548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .B(_836_),
    .C(_825_),
    .Y(_871_)
);

NAND2X1 _4549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_818_),
    .Y(_872_)
);

XOR2X1 _4550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_872_),
    .B(_697_),
    .Y(_873_)
);

INVX2 _4551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .Y(_874_)
);

OAI21X1 _4552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(_823_),
    .C(_811_),
    .Y(_876_)
);

NAND2X1 _4553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_713_),
    .B(_718_),
    .Y(_877_)
);

NOR2X1 _4554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_2608_),
    .Y(_878_)
);

INVX2 _4555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_878_),
    .Y(_879_)
);

OAI21X1 _4556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_700_),
    .C(_705_),
    .Y(_880_)
);

NAND2X1 _4557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_14_bF$buf3),
    .Y(_881_)
);

NOR2X1 _4558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_881_),
    .Y(_882_)
);

AOI22X1 _4559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_14_bF$buf2),
    .C(breg_7_bF$buf2),
    .D(areg_11_bF$buf1),
    .Y(_883_)
);

OAI21X1 _4560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .B(_883_),
    .C(_696_),
    .Y(_884_)
);

INVX1 _4561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .Y(_885_)
);

OR2X2 _4562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_339_),
    .B(_881_),
    .Y(_887_)
);

INVX1 _4563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .Y(_888_)
);

NAND3X1 _4564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .B(_888_),
    .C(_887_),
    .Y(_889_)
);

AOI21X1 _4565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_889_),
    .C(_880_),
    .Y(_890_)
);

AOI21X1 _4566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_706_),
    .C(_709_),
    .Y(_891_)
);

AOI21X1 _4567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_888_),
    .B(_887_),
    .C(_885_),
    .Y(_892_)
);

NOR3X1 _4568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_883_),
    .C(_882_),
    .Y(_893_)
);

NOR3X1 _4569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .B(_891_),
    .C(_892_),
    .Y(_894_)
);

OAI21X1 _4570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_894_),
    .B(_890_),
    .C(_879_),
    .Y(_895_)
);

OAI21X1 _4571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_893_),
    .C(_891_),
    .Y(_896_)
);

NAND3X1 _4572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_880_),
    .C(_889_),
    .Y(_898_)
);

NAND3X1 _4573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_878_),
    .B(_898_),
    .C(_896_),
    .Y(_899_)
);

AOI21X1 _4574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(_752_),
    .C(_754_),
    .Y(_900_)
);

OAI21X1 _4575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_900_),
    .B(_762_),
    .C(_755_),
    .Y(_901_)
);

NAND3X1 _4576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_899_),
    .B(_901_),
    .C(_895_),
    .Y(_902_)
);

AOI21X1 _4577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_898_),
    .B(_896_),
    .C(_878_),
    .Y(_903_)
);

NOR3X1 _4578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_879_),
    .C(_894_),
    .Y(_904_)
);

INVX1 _4579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_755_),
    .Y(_905_)
);

AOI21X1 _4580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_760_),
    .B(_741_),
    .C(_905_),
    .Y(_906_)
);

OAI21X1 _4581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_904_),
    .B(_903_),
    .C(_906_),
    .Y(_907_)
);

NAND3X1 _4582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_902_),
    .C(_907_),
    .Y(_909_)
);

AND2X2 _4583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_713_),
    .Y(_910_)
);

NAND3X1 _4584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_899_),
    .C(_906_),
    .Y(_911_)
);

OAI21X1 _4585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_904_),
    .B(_903_),
    .C(_901_),
    .Y(_912_)
);

NAND3X1 _4586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_910_),
    .B(_911_),
    .C(_912_),
    .Y(_913_)
);

NAND2X1 _4587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(_913_),
    .Y(_914_)
);

AOI21X1 _4588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .B(_798_),
    .C(_769_),
    .Y(_915_)
);

OAI21X1 _4589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_915_),
    .B(_807_),
    .C(_799_),
    .Y(_916_)
);

NAND2X1 _4590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_749_),
    .Y(_917_)
);

NAND2X1 _4591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_15_bF$buf1),
    .Y(_918_)
);

AOI22X1 _4592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf0),
    .B(areg_10_bF$buf0),
    .C(breg_9_bF$buf1),
    .D(areg[9]),
    .Y(_920_)
);

NOR2X1 _4593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_565_),
    .Y(_921_)
);

OAI21X1 _4594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_),
    .B(_920_),
    .C(_918_),
    .Y(_922_)
);

INVX1 _4595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .Y(_923_)
);

INVX1 _4596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .Y(_924_)
);

OR2X2 _4597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_565_),
    .Y(_925_)
);

NAND3X1 _4598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_924_),
    .C(_925_),
    .Y(_926_)
);

NAND2X1 _4599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_772_),
    .Y(_927_)
);

OAI21X1 _4600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_770_),
    .B(_773_),
    .C(_927_),
    .Y(_928_)
);

NAND3X1 _4601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_928_),
    .B(_922_),
    .C(_926_),
    .Y(_929_)
);

AOI21X1 _4602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_924_),
    .B(_925_),
    .C(_923_),
    .Y(_931_)
);

NOR3X1 _4603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(_920_),
    .C(_921_),
    .Y(_932_)
);

INVX1 _4604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .Y(_933_)
);

AOI22X1 _4605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_771_),
    .B(_772_),
    .C(_933_),
    .D(_794_),
    .Y(_934_)
);

OAI21X1 _4606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_932_),
    .C(_934_),
    .Y(_935_)
);

NAND3X1 _4607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_929_),
    .C(_935_),
    .Y(_936_)
);

AOI21X1 _4608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_746_),
    .C(_757_),
    .Y(_937_)
);

NAND3X1 _4609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_922_),
    .C(_926_),
    .Y(_938_)
);

OAI21X1 _4610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_932_),
    .C(_928_),
    .Y(_939_)
);

NAND3X1 _4611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_937_),
    .B(_938_),
    .C(_939_),
    .Y(_940_)
);

NAND2X1 _4612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(_940_),
    .Y(_942_)
);

AOI21X1 _4613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_784_),
    .C(_776_),
    .Y(_943_)
);

OAI21X1 _4614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_943_),
    .B(_795_),
    .C(_787_),
    .Y(_944_)
);

NAND2X1 _4615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_10_bF$buf1),
    .Y(_945_)
);

INVX2 _4616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .Y(_946_)
);

AND2X2 _4617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_12_bF$buf2),
    .Y(_947_)
);

AOI22X1 _4618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_12_bF$buf1),
    .C(areg_7_bF$buf3),
    .D(breg_11_bF$buf0),
    .Y(_948_)
);

AOI21X1 _4619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_947_),
    .C(_948_),
    .Y(_949_)
);

XNOR2X1 _4620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_946_),
    .Y(_950_)
);

OAI21X1 _4621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_782_),
    .C(_781_),
    .Y(_951_)
);

NAND2X1 _4622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_13_bF$buf3),
    .Y(_953_)
);

NAND2X1 _4623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_14_bF$buf3),
    .Y(_954_)
);

NAND3X1 _4624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_15_bF$buf2),
    .C(_954_),
    .Y(_955_)
);

NAND2X1 _4625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_15_bF$buf1),
    .Y(_956_)
);

NAND3X1 _4626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_14_bF$buf2),
    .C(_956_),
    .Y(_957_)
);

AOI21X1 _4627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_957_),
    .C(_953_),
    .Y(_958_)
);

INVX2 _4628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_953_),
    .Y(_959_)
);

AND2X2 _4629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_15_bF$buf0),
    .Y(_960_)
);

NAND2X1 _4630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .B(_960_),
    .Y(_961_)
);

AOI22X1 _4631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_15_bF$buf3),
    .C(areg_4_bF$buf1),
    .D(breg_14_bF$buf1),
    .Y(_962_)
);

INVX2 _4632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .Y(_964_)
);

AOI21X1 _4633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(_961_),
    .C(_959_),
    .Y(_965_)
);

OAI21X1 _4634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_958_),
    .C(_951_),
    .Y(_966_)
);

AOI21X1 _4635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_783_),
    .C(_785_),
    .Y(_967_)
);

NAND3X1 _4636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_959_),
    .B(_964_),
    .C(_961_),
    .Y(_968_)
);

NAND2X1 _4637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_15_bF$buf2),
    .Y(_969_)
);

NOR2X1 _4638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_969_),
    .Y(_970_)
);

OAI21X1 _4639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_970_),
    .B(_962_),
    .C(_953_),
    .Y(_971_)
);

NAND3X1 _4640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_967_),
    .C(_968_),
    .Y(_972_)
);

AOI21X1 _4641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_972_),
    .B(_966_),
    .C(_950_),
    .Y(_973_)
);

XNOR2X1 _4642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_945_),
    .Y(_975_)
);

NAND3X1 _4643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .B(_971_),
    .C(_968_),
    .Y(_976_)
);

OAI21X1 _4644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_958_),
    .C(_967_),
    .Y(_977_)
);

AOI21X1 _4645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(_977_),
    .C(_975_),
    .Y(_978_)
);

OAI21X1 _4646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_978_),
    .C(_944_),
    .Y(_979_)
);

NOR3X1 _4647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_788_),
    .C(_791_),
    .Y(_980_)
);

AOI21X1 _4648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_792_),
    .C(_980_),
    .Y(_981_)
);

NAND3X1 _4649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_976_),
    .C(_977_),
    .Y(_982_)
);

NAND3X1 _4650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(_972_),
    .C(_966_),
    .Y(_983_)
);

NAND3X1 _4651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .B(_983_),
    .C(_981_),
    .Y(_984_)
);

AOI21X1 _4652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(_984_),
    .C(_942_),
    .Y(_986_)
);

AND2X2 _4653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(_940_),
    .Y(_987_)
);

NAND3X1 _4654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_944_),
    .B(_982_),
    .C(_983_),
    .Y(_988_)
);

OAI21X1 _4655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_978_),
    .C(_981_),
    .Y(_989_)
);

AOI21X1 _4656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_989_),
    .C(_987_),
    .Y(_990_)
);

OAI21X1 _4657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_990_),
    .C(_916_),
    .Y(_991_)
);

NOR3X1 _4658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_804_),
    .C(_802_),
    .Y(_992_)
);

AOI21X1 _4659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_766_),
    .B(_805_),
    .C(_992_),
    .Y(_993_)
);

NAND3X1 _4660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_989_),
    .C(_987_),
    .Y(_994_)
);

NAND3X1 _4661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_979_),
    .C(_984_),
    .Y(_995_)
);

NAND3X1 _4662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_995_),
    .C(_993_),
    .Y(_997_)
);

AOI21X1 _4663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .B(_997_),
    .C(_914_),
    .Y(_998_)
);

NAND3X1 _4664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_910_),
    .B(_902_),
    .C(_907_),
    .Y(_999_)
);

NAND3X1 _4665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_911_),
    .C(_912_),
    .Y(_1000_)
);

NAND2X1 _4666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_999_),
    .B(_1000_),
    .Y(_1001_)
);

NAND3X1 _4667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_994_),
    .C(_995_),
    .Y(_1002_)
);

OAI21X1 _4668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_990_),
    .C(_993_),
    .Y(_1003_)
);

AOI21X1 _4669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_1003_),
    .C(_1001_),
    .Y(_1004_)
);

OAI21X1 _4670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_1004_),
    .C(_876_),
    .Y(_1005_)
);

AOI21X1 _4671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_738_),
    .C(_822_),
    .Y(_1006_)
);

NAND3X1 _4672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_1001_),
    .C(_1003_),
    .Y(_1008_)
);

NAND3X1 _4673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_991_),
    .C(_997_),
    .Y(_1009_)
);

NAND3X1 _4674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1009_),
    .C(_1006_),
    .Y(_1010_)
);

AOI21X1 _4675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1005_),
    .B(_1010_),
    .C(_874_),
    .Y(_1011_)
);

NAND3X1 _4676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1009_),
    .C(_876_),
    .Y(_1012_)
);

OAI21X1 _4677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_1004_),
    .C(_1006_),
    .Y(_1013_)
);

AOI21X1 _4678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1012_),
    .B(_1013_),
    .C(_873_),
    .Y(_1014_)
);

OAI21X1 _4679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(_1014_),
    .C(_871_),
    .Y(_1015_)
);

AOI21X1 _4680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_831_),
    .C(_835_),
    .Y(_1016_)
);

NAND3X1 _4681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_1012_),
    .C(_1013_),
    .Y(_1017_)
);

NOR3X1 _4682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_1004_),
    .C(_1006_),
    .Y(_1019_)
);

AOI21X1 _4683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1009_),
    .C(_876_),
    .Y(_1020_)
);

OAI21X1 _4684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(_1020_),
    .C(_874_),
    .Y(_1021_)
);

NAND3X1 _4685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(_1016_),
    .C(_1021_),
    .Y(_1022_)
);

AOI21X1 _4686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1015_),
    .B(_1022_),
    .C(_870_),
    .Y(_1023_)
);

INVX2 _4687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .Y(_1024_)
);

NAND3X1 _4688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(_1021_),
    .C(_871_),
    .Y(_1025_)
);

OAI21X1 _4689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(_1014_),
    .C(_1016_),
    .Y(_1026_)
);

AOI21X1 _4690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1026_),
    .B(_1025_),
    .C(_1024_),
    .Y(_1027_)
);

OAI21X1 _4691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1027_),
    .B(_1023_),
    .C(_869_),
    .Y(_1028_)
);

AOI21X1 _4692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_845_),
    .C(_847_),
    .Y(_1030_)
);

NAND3X1 _4693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1026_),
    .C(_1025_),
    .Y(_1031_)
);

NOR3X1 _4694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(_1014_),
    .C(_1016_),
    .Y(_1032_)
);

AOI21X1 _4695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(_1021_),
    .C(_871_),
    .Y(_1033_)
);

OAI21X1 _4696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1032_),
    .B(_1033_),
    .C(_870_),
    .Y(_1034_)
);

NAND3X1 _4697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(_1030_),
    .C(_1034_),
    .Y(_1035_)
);

NAND2X1 _4698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1028_),
    .B(_1035_),
    .Y(_1036_)
);

AND2X2 _4699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_1036_),
    .Y(_1037_)
);

NOR2X1 _4700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_868_),
    .Y(_1038_)
);

NOR2X1 _4701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1038_),
    .B(_1037_),
    .Y(_1_[18])
);

NAND3X1 _4702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(_869_),
    .C(_1034_),
    .Y(_1040_)
);

INVX1 _4703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .Y(_1041_)
);

NOR2X1 _4704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1041_),
    .B(_1037_),
    .Y(_1042_)
);

OAI21X1 _4705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(_870_),
    .C(_1025_),
    .Y(_1043_)
);

NAND2X1 _4706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(_872_),
    .Y(_1044_)
);

OAI21X1 _4707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_1020_),
    .C(_1012_),
    .Y(_1045_)
);

NAND2X1 _4708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_902_),
    .B(_909_),
    .Y(_1046_)
);

INVX1 _4709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .Y(_1047_)
);

AOI21X1 _4710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_995_),
    .C(_916_),
    .Y(_1048_)
);

OAI21X1 _4711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_1048_),
    .C(_1002_),
    .Y(_1049_)
);

OAI21X1 _4712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_879_),
    .C(_898_),
    .Y(_1051_)
);

OAI21X1 _4713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_883_),
    .C(_887_),
    .Y(_1052_)
);

NOR2X1 _4714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_2608_),
    .Y(_1053_)
);

NAND2X1 _4715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_13_bF$buf0),
    .Y(_1054_)
);

NAND2X1 _4716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg_14_bF$buf1),
    .Y(_1055_)
);

XOR2X1 _4717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(_1055_),
    .Y(_1056_)
);

NAND2X1 _4718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1056_),
    .Y(_1057_)
);

NAND2X1 _4719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_14_bF$buf0),
    .Y(_1058_)
);

INVX1 _4720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .Y(_1059_)
);

OAI21X1 _4721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_1059_),
    .C(_1054_),
    .Y(_1060_)
);

OAI21X1 _4722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_1058_),
    .C(_1060_),
    .Y(_1062_)
);

OAI21X1 _4723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_2608_),
    .C(_1062_),
    .Y(_1063_)
);

NAND3X1 _4724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .B(_1063_),
    .C(_1057_),
    .Y(_1064_)
);

INVX1 _4725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .Y(_1065_)
);

OAI21X1 _4726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_2608_),
    .C(_1056_),
    .Y(_1066_)
);

NAND2X1 _4727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1062_),
    .Y(_1067_)
);

NAND3X1 _4728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1067_),
    .B(_1065_),
    .C(_1066_),
    .Y(_1068_)
);

AND2X2 _4729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1068_),
    .B(_1064_),
    .Y(_1069_)
);

AOI21X1 _4730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .B(_926_),
    .C(_928_),
    .Y(_1070_)
);

OAI21X1 _4731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1070_),
    .B(_937_),
    .C(_929_),
    .Y(_1071_)
);

NAND2X1 _4732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1071_),
    .B(_1069_),
    .Y(_1073_)
);

NAND2X1 _4733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1068_),
    .Y(_1074_)
);

INVX1 _4734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_929_),
    .Y(_1075_)
);

AOI21X1 _4735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_935_),
    .C(_1075_),
    .Y(_1076_)
);

NAND2X1 _4736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1074_),
    .B(_1076_),
    .Y(_1077_)
);

NAND3X1 _4737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .B(_1077_),
    .C(_1073_),
    .Y(_1078_)
);

INVX1 _4738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .Y(_1079_)
);

NAND2X1 _4739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1076_),
    .B(_1069_),
    .Y(_1080_)
);

NAND2X1 _4740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1071_),
    .B(_1074_),
    .Y(_1081_)
);

NAND3X1 _4741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1081_),
    .B(_1079_),
    .C(_1080_),
    .Y(_1082_)
);

NAND2X1 _4742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(_1078_),
    .Y(_1084_)
);

AOI21X1 _4743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .B(_983_),
    .C(_944_),
    .Y(_1085_)
);

OAI21X1 _4744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_942_),
    .C(_988_),
    .Y(_1086_)
);

OAI21X1 _4745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_918_),
    .B(_920_),
    .C(_925_),
    .Y(_1087_)
);

INVX1 _4746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .Y(_1088_)
);

NAND2X1 _4747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf3),
    .B(areg_11_bF$buf0),
    .Y(_1089_)
);

NAND2X1 _4748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_15_bF$buf0),
    .Y(_1090_)
);

NOR2X1 _4749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_1090_),
    .Y(_1091_)
);

AOI22X1 _4750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_15_bF$buf3),
    .C(breg_9_bF$buf3),
    .D(areg_10_bF$buf3),
    .Y(_1092_)
);

OAI21X1 _4751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1091_),
    .B(_1092_),
    .C(_1089_),
    .Y(_1093_)
);

INVX2 _4752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .Y(_1095_)
);

OR2X2 _4753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_147_),
    .B(_1090_),
    .Y(_1096_)
);

INVX1 _4754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .Y(_1097_)
);

NAND3X1 _4755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1095_),
    .B(_1097_),
    .C(_1096_),
    .Y(_1098_)
);

NAND2X1 _4756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_947_),
    .Y(_1099_)
);

OAI21X1 _4757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_948_),
    .C(_1099_),
    .Y(_1100_)
);

NAND3X1 _4758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .B(_1093_),
    .C(_1098_),
    .Y(_1101_)
);

AOI21X1 _4759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1097_),
    .B(_1096_),
    .C(_1095_),
    .Y(_1102_)
);

NOR3X1 _4760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1092_),
    .C(_1091_),
    .Y(_1103_)
);

AOI22X1 _4761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_947_),
    .C(_949_),
    .D(_946_),
    .Y(_1104_)
);

OAI21X1 _4762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1103_),
    .C(_1104_),
    .Y(_1105_)
);

NAND3X1 _4763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_1101_),
    .C(_1105_),
    .Y(_1106_)
);

NAND3X1 _4764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1093_),
    .B(_1098_),
    .C(_1104_),
    .Y(_1107_)
);

OAI21X1 _4765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1103_),
    .C(_1100_),
    .Y(_1108_)
);

NAND3X1 _4766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .B(_1108_),
    .C(_1107_),
    .Y(_1109_)
);

AND2X2 _4767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .B(_1106_),
    .Y(_1110_)
);

AOI21X1 _4768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_968_),
    .C(_951_),
    .Y(_1111_)
);

OAI21X1 _4769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1111_),
    .B(_950_),
    .C(_976_),
    .Y(_1112_)
);

NAND2X1 _4770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_10_bF$buf0),
    .Y(_1113_)
);

INVX1 _4771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1113_),
    .Y(_1114_)
);

AND2X2 _4772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_11_bF$buf3),
    .Y(_1116_)
);

AND2X2 _4773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_12_bF$buf0),
    .Y(_1117_)
);

AOI22X1 _4774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf1),
    .B(breg_12_bF$buf3),
    .C(areg_8_bF$buf2),
    .D(breg_11_bF$buf2),
    .Y(_1118_)
);

AOI21X1 _4775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .B(_1117_),
    .C(_1118_),
    .Y(_1119_)
);

XNOR2X1 _4776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(_1114_),
    .Y(_1120_)
);

OAI21X1 _4777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_953_),
    .B(_962_),
    .C(_961_),
    .Y(_1121_)
);

NAND2X1 _4778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_13_bF$buf2),
    .Y(_1122_)
);

NAND2X1 _4779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_14_bF$buf0),
    .Y(_1123_)
);

NAND3X1 _4780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_15_bF$buf1),
    .C(_1123_),
    .Y(_1124_)
);

NAND3X1 _4781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_14_bF$buf3),
    .C(_969_),
    .Y(_1125_)
);

AOI21X1 _4782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1125_),
    .C(_1122_),
    .Y(_1128_)
);

INVX2 _4783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1122_),
    .Y(_1129_)
);

AND2X2 _4784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_14_bF$buf2),
    .Y(_1130_)
);

NAND2X1 _4785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(_1130_),
    .Y(_1131_)
);

OAI21X1 _4786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_220_),
    .C(_969_),
    .Y(_1132_)
);

AOI21X1 _4787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1132_),
    .B(_1131_),
    .C(_1129_),
    .Y(_1133_)
);

OAI21X1 _4788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(_1128_),
    .C(_1121_),
    .Y(_1134_)
);

AOI21X1 _4789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_959_),
    .B(_964_),
    .C(_970_),
    .Y(_1135_)
);

NAND3X1 _4790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .B(_1132_),
    .C(_1131_),
    .Y(_1136_)
);

NAND3X1 _4791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1122_),
    .B(_1124_),
    .C(_1125_),
    .Y(_1137_)
);

NAND3X1 _4792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1135_),
    .C(_1136_),
    .Y(_1139_)
);

AOI21X1 _4793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1134_),
    .C(_1120_),
    .Y(_1140_)
);

XNOR2X1 _4794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(_1113_),
    .Y(_1141_)
);

NAND3X1 _4795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1121_),
    .B(_1137_),
    .C(_1136_),
    .Y(_1142_)
);

OAI21X1 _4796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .B(_1128_),
    .C(_1135_),
    .Y(_1143_)
);

AOI21X1 _4797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1143_),
    .C(_1141_),
    .Y(_1144_)
);

OAI21X1 _4798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1140_),
    .B(_1144_),
    .C(_1112_),
    .Y(_1145_)
);

NOR3X1 _4799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_967_),
    .B(_958_),
    .C(_965_),
    .Y(_1146_)
);

AOI21X1 _4800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_975_),
    .B(_977_),
    .C(_1146_),
    .Y(_1147_)
);

NAND3X1 _4801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1142_),
    .C(_1143_),
    .Y(_1148_)
);

NAND3X1 _4802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1120_),
    .B(_1139_),
    .C(_1134_),
    .Y(_1150_)
);

NAND3X1 _4803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .B(_1150_),
    .C(_1147_),
    .Y(_1151_)
);

AOI21X1 _4804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1151_),
    .B(_1145_),
    .C(_1110_),
    .Y(_1152_)
);

NAND2X1 _4805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1106_),
    .B(_1109_),
    .Y(_1153_)
);

NAND3X1 _4806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_1148_),
    .C(_1150_),
    .Y(_1154_)
);

OAI21X1 _4807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1140_),
    .B(_1144_),
    .C(_1147_),
    .Y(_1155_)
);

AOI21X1 _4808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1155_),
    .C(_1153_),
    .Y(_1156_)
);

OAI21X1 _4809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1156_),
    .C(_1086_),
    .Y(_1157_)
);

NOR3X1 _4810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_978_),
    .C(_981_),
    .Y(_1158_)
);

AOI21X1 _4811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_987_),
    .B(_989_),
    .C(_1158_),
    .Y(_1159_)
);

NAND3X1 _4812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1153_),
    .C(_1155_),
    .Y(_1161_)
);

NAND3X1 _4813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1151_),
    .B(_1145_),
    .C(_1110_),
    .Y(_1162_)
);

NAND3X1 _4814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1161_),
    .B(_1162_),
    .C(_1159_),
    .Y(_1163_)
);

AOI21X1 _4815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1163_),
    .B(_1157_),
    .C(_1084_),
    .Y(_1164_)
);

NAND3X1 _4816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1079_),
    .B(_1077_),
    .C(_1073_),
    .Y(_1165_)
);

NAND3X1 _4817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .B(_1081_),
    .C(_1080_),
    .Y(_1166_)
);

NAND2X1 _4818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1165_),
    .Y(_1167_)
);

NAND3X1 _4819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1086_),
    .B(_1161_),
    .C(_1162_),
    .Y(_1168_)
);

OAI21X1 _4820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1156_),
    .C(_1159_),
    .Y(_1169_)
);

AOI21X1 _4821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1169_),
    .C(_1167_),
    .Y(_1170_)
);

OAI21X1 _4822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1170_),
    .C(_1049_),
    .Y(_1172_)
);

NOR3X1 _4823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_990_),
    .C(_993_),
    .Y(_1173_)
);

AOI21X1 _4824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1001_),
    .B(_1003_),
    .C(_1173_),
    .Y(_1174_)
);

NAND3X1 _4825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(_1168_),
    .C(_1169_),
    .Y(_1175_)
);

NAND3X1 _4826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1084_),
    .B(_1163_),
    .C(_1157_),
    .Y(_1176_)
);

NAND3X1 _4827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1176_),
    .C(_1174_),
    .Y(_1177_)
);

AOI21X1 _4828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1177_),
    .B(_1172_),
    .C(_1047_),
    .Y(_1178_)
);

NAND3X1 _4829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1176_),
    .C(_1049_),
    .Y(_1179_)
);

OAI21X1 _4830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1170_),
    .C(_1174_),
    .Y(_1180_)
);

AOI21X1 _4831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .B(_1180_),
    .C(_1046_),
    .Y(_1181_)
);

OAI21X1 _4832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1181_),
    .C(_1045_),
    .Y(_1183_)
);

AOI21X1 _4833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_1013_),
    .C(_1019_),
    .Y(_1184_)
);

NAND3X1 _4834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .B(_1179_),
    .C(_1180_),
    .Y(_1185_)
);

NAND3X1 _4835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1177_),
    .C(_1172_),
    .Y(_1186_)
);

NAND3X1 _4836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1186_),
    .C(_1184_),
    .Y(_1187_)
);

AOI21X1 _4837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1187_),
    .B(_1183_),
    .C(_1044_),
    .Y(_1188_)
);

INVX2 _4838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1044_),
    .Y(_1189_)
);

NAND3X1 _4839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1186_),
    .C(_1045_),
    .Y(_1190_)
);

OAI21X1 _4840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1181_),
    .C(_1184_),
    .Y(_1191_)
);

AOI21X1 _4841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1190_),
    .B(_1191_),
    .C(_1189_),
    .Y(_1192_)
);

OAI21X1 _4842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1188_),
    .B(_1192_),
    .C(_1043_),
    .Y(_1194_)
);

AOI21X1 _4843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1026_),
    .C(_1032_),
    .Y(_1195_)
);

NAND3X1 _4844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1189_),
    .B(_1190_),
    .C(_1191_),
    .Y(_1196_)
);

NOR3X1 _4845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1181_),
    .C(_1184_),
    .Y(_1197_)
);

AOI21X1 _4846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1186_),
    .C(_1045_),
    .Y(_1198_)
);

OAI21X1 _4847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1198_),
    .C(_1044_),
    .Y(_1199_)
);

NAND3X1 _4848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1195_),
    .C(_1199_),
    .Y(_1200_)
);

NAND2X1 _4849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(_1200_),
    .Y(_1201_)
);

XNOR2X1 _4850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_1201_),
    .Y(_1_[19])
);

AOI22X1 _4851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(_1200_),
    .C(_1035_),
    .D(_1028_),
    .Y(_1202_)
);

NAND3X1 _4852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1043_),
    .C(_1199_),
    .Y(_1204_)
);

AOI21X1 _4853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1199_),
    .C(_1043_),
    .Y(_1205_)
);

AOI21X1 _4854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1204_),
    .B(_1040_),
    .C(_1205_),
    .Y(_1206_)
);

AOI21X1 _4855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_854_),
    .C(_1206_),
    .Y(_1207_)
);

NAND2X1 _4856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_866_),
    .Y(_1208_)
);

OAI21X1 _4857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_1208_),
    .C(_1207_),
    .Y(_1209_)
);

OAI21X1 _4858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1198_),
    .B(_1044_),
    .C(_1190_),
    .Y(_1210_)
);

INVX1 _4859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .Y(_1211_)
);

AOI21X1 _4860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .B(_1180_),
    .C(_1211_),
    .Y(_1212_)
);

OAI21X1 _4861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1074_),
    .B(_1076_),
    .C(_1078_),
    .Y(_1213_)
);

INVX2 _4862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .Y(_1215_)
);

NAND2X1 _4863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1175_),
    .Y(_1216_)
);

INVX1 _4864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .Y(_1217_)
);

OAI21X1 _4865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_1058_),
    .C(_1057_),
    .Y(_1218_)
);

NAND2X1 _4866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf2),
    .B(areg_13_bF$buf3),
    .Y(_1219_)
);

INVX2 _4867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1220_)
);

NAND2X1 _4868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1053_),
    .Y(_1221_)
);

INVX1 _4869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .Y(_1222_)
);

AOI22X1 _4870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf1),
    .B(areg_13_bF$buf2),
    .C(breg_8_bF$buf1),
    .D(areg[12]),
    .Y(_1223_)
);

NOR2X1 _4871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1223_),
    .B(_1222_),
    .Y(_1224_)
);

XOR2X1 _4872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(_1224_),
    .Y(_1226_)
);

NAND2X1 _4873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .B(_1105_),
    .Y(_1227_)
);

OAI21X1 _4874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1227_),
    .B(_1088_),
    .C(_1101_),
    .Y(_1228_)
);

NAND2X1 _4875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1228_),
    .Y(_1229_)
);

XNOR2X1 _4876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(_1224_),
    .Y(_1230_)
);

INVX1 _4877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .Y(_1231_)
);

AOI21X1 _4878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .B(_1105_),
    .C(_1231_),
    .Y(_1232_)
);

NAND2X1 _4879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(_1230_),
    .Y(_1233_)
);

NAND3X1 _4880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1217_),
    .B(_1233_),
    .C(_1229_),
    .Y(_1234_)
);

NAND2X1 _4881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(_1226_),
    .Y(_1235_)
);

NAND2X1 _4882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1228_),
    .Y(_1237_)
);

NAND3X1 _4883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1235_),
    .C(_1237_),
    .Y(_1238_)
);

NAND2X1 _4884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1234_),
    .B(_1238_),
    .Y(_1239_)
);

AOI21X1 _4885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .B(_1150_),
    .C(_1112_),
    .Y(_1240_)
);

OAI21X1 _4886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1110_),
    .B(_1240_),
    .C(_1154_),
    .Y(_1241_)
);

OAI21X1 _4887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1092_),
    .C(_1096_),
    .Y(_1242_)
);

NOR2X1 _4888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_1090_),
    .Y(_1243_)
);

AOI22X1 _4889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf0),
    .B(areg_15_bF$buf2),
    .C(breg_9_bF$buf2),
    .D(areg_11_bF$buf3),
    .Y(_1244_)
);

OAI21X1 _4890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(_1244_),
    .C(_1058_),
    .Y(_1245_)
);

INVX1 _4891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .Y(_1246_)
);

OR2X2 _4892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_1090_),
    .Y(_1248_)
);

OAI21X1 _4893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2266_),
    .B(_2458_),
    .C(_335_),
    .Y(_1249_)
);

NAND3X1 _4894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1246_),
    .B(_1249_),
    .C(_1248_),
    .Y(_1250_)
);

NAND2X1 _4895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .B(_1117_),
    .Y(_1251_)
);

OAI21X1 _4896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1113_),
    .B(_1118_),
    .C(_1251_),
    .Y(_1252_)
);

NAND3X1 _4897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1252_),
    .B(_1245_),
    .C(_1250_),
    .Y(_1253_)
);

INVX1 _4898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1245_),
    .Y(_1254_)
);

OAI21X1 _4899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_1090_),
    .C(_1249_),
    .Y(_1255_)
);

NOR2X1 _4900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(_1255_),
    .Y(_1256_)
);

INVX1 _4901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1252_),
    .Y(_1257_)
);

OAI21X1 _4902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1256_),
    .B(_1254_),
    .C(_1257_),
    .Y(_1259_)
);

NAND3X1 _4903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .B(_1253_),
    .C(_1259_),
    .Y(_1260_)
);

INVX1 _4904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .Y(_1261_)
);

NAND3X1 _4905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1245_),
    .B(_1250_),
    .C(_1257_),
    .Y(_1262_)
);

OAI21X1 _4906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1256_),
    .B(_1254_),
    .C(_1252_),
    .Y(_1263_)
);

NAND3X1 _4907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1261_),
    .B(_1262_),
    .C(_1263_),
    .Y(_1264_)
);

NAND2X1 _4908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1260_),
    .B(_1264_),
    .Y(_1265_)
);

AOI21X1 _4909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1136_),
    .C(_1121_),
    .Y(_1266_)
);

OAI21X1 _4910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1120_),
    .C(_1142_),
    .Y(_1267_)
);

NAND2X1 _4911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf3),
    .B(areg_10_bF$buf2),
    .Y(_1268_)
);

INVX2 _4912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1268_),
    .Y(_1270_)
);

NAND2X1 _4913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf1),
    .B(breg_11_bF$buf1),
    .Y(_1271_)
);

NAND2X1 _4914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_12_bF$buf2),
    .Y(_1272_)
);

NAND2X1 _4915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_11_bF$buf0),
    .Y(_1273_)
);

OAI21X1 _4916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_2698_),
    .C(_1273_),
    .Y(_1274_)
);

OAI21X1 _4917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1271_),
    .B(_1272_),
    .C(_1274_),
    .Y(_1275_)
);

XNOR2X1 _4918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(_1270_),
    .Y(_1276_)
);

NOR2X1 _4919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(_1130_),
    .Y(_1277_)
);

OAI21X1 _4920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(_1122_),
    .C(_1131_),
    .Y(_1278_)
);

NAND2X1 _4921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_13_bF$buf1),
    .Y(_1279_)
);

INVX2 _4922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1279_),
    .Y(_1281_)
);

AND2X2 _4923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_15_bF$buf0),
    .Y(_1282_)
);

NAND2X1 _4924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1130_),
    .B(_1282_),
    .Y(_1283_)
);

AOI22X1 _4925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_15_bF$buf3),
    .C(areg[6]),
    .D(breg_14_bF$buf1),
    .Y(_1284_)
);

INVX2 _4926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1284_),
    .Y(_1285_)
);

NAND3X1 _4927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1285_),
    .C(_1283_),
    .Y(_1286_)
);

NAND2X1 _4928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .B(breg_15_bF$buf2),
    .Y(_1287_)
);

NOR2X1 _4929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(_1287_),
    .Y(_1288_)
);

OAI21X1 _4930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1288_),
    .B(_1284_),
    .C(_1279_),
    .Y(_1289_)
);

NAND3X1 _4931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1286_),
    .B(_1289_),
    .C(_1278_),
    .Y(_1290_)
);

NOR2X1 _4932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_1123_),
    .Y(_1292_)
);

AOI21X1 _4933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .B(_1132_),
    .C(_1292_),
    .Y(_1293_)
);

NOR3X1 _4934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1279_),
    .B(_1284_),
    .C(_1288_),
    .Y(_1294_)
);

AOI21X1 _4935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1285_),
    .B(_1283_),
    .C(_1281_),
    .Y(_1295_)
);

OAI21X1 _4936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1294_),
    .C(_1293_),
    .Y(_1296_)
);

NAND3X1 _4937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1296_),
    .C(_1276_),
    .Y(_1297_)
);

XNOR2X1 _4938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(_1268_),
    .Y(_1298_)
);

NOR3X1 _4939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1294_),
    .B(_1293_),
    .C(_1295_),
    .Y(_1299_)
);

AOI21X1 _4940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1286_),
    .B(_1289_),
    .C(_1278_),
    .Y(_1300_)
);

OAI21X1 _4941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(_1300_),
    .C(_1298_),
    .Y(_1301_)
);

AOI21X1 _4942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1297_),
    .B(_1301_),
    .C(_1267_),
    .Y(_1303_)
);

NOR3X1 _4943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .B(_1128_),
    .C(_1133_),
    .Y(_1304_)
);

AOI21X1 _4944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1143_),
    .C(_1304_),
    .Y(_1305_)
);

OAI21X1 _4945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1294_),
    .C(_1278_),
    .Y(_1306_)
);

NAND3X1 _4946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1289_),
    .C(_1286_),
    .Y(_1307_)
);

AOI21X1 _4947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1307_),
    .B(_1306_),
    .C(_1298_),
    .Y(_1308_)
);

AOI21X1 _4948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1290_),
    .C(_1276_),
    .Y(_1309_)
);

NOR3X1 _4949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1308_),
    .B(_1305_),
    .C(_1309_),
    .Y(_1310_)
);

OAI21X1 _4950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1310_),
    .B(_1303_),
    .C(_1265_),
    .Y(_1311_)
);

AOI21X1 _4951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1262_),
    .B(_1263_),
    .C(_1261_),
    .Y(_1312_)
);

AOI21X1 _4952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .B(_1259_),
    .C(_1242_),
    .Y(_1314_)
);

NOR2X1 _4953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(_1314_),
    .Y(_1315_)
);

OAI21X1 _4954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1309_),
    .B(_1308_),
    .C(_1305_),
    .Y(_1316_)
);

NAND3X1 _4955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1297_),
    .C(_1301_),
    .Y(_1317_)
);

NAND3X1 _4956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1317_),
    .C(_1315_),
    .Y(_1318_)
);

AOI21X1 _4957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1318_),
    .C(_1241_),
    .Y(_1319_)
);

NOR3X1 _4958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1140_),
    .B(_1144_),
    .C(_1147_),
    .Y(_1320_)
);

AOI21X1 _4959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1153_),
    .B(_1155_),
    .C(_1320_),
    .Y(_1321_)
);

AOI21X1 _4960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1317_),
    .C(_1315_),
    .Y(_1322_)
);

NOR3X1 _4961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(_1303_),
    .C(_1310_),
    .Y(_1323_)
);

NOR3X1 _4962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .B(_1322_),
    .C(_1323_),
    .Y(_1325_)
);

NOR3X1 _4963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .B(_1319_),
    .C(_1325_),
    .Y(_1326_)
);

AND2X2 _4964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .B(_1234_),
    .Y(_1327_)
);

OAI21X1 _4965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1323_),
    .B(_1322_),
    .C(_1321_),
    .Y(_1328_)
);

NAND3X1 _4966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1311_),
    .C(_1318_),
    .Y(_1329_)
);

AOI21X1 _4967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1329_),
    .B(_1328_),
    .C(_1327_),
    .Y(_1330_)
);

OAI21X1 _4968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(_1330_),
    .C(_1216_),
    .Y(_1331_)
);

INVX1 _4969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .Y(_1332_)
);

AOI21X1 _4970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(_1169_),
    .C(_1332_),
    .Y(_1333_)
);

NAND3X1 _4971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1328_),
    .B(_1329_),
    .C(_1327_),
    .Y(_1334_)
);

OAI21X1 _4972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1325_),
    .B(_1319_),
    .C(_1239_),
    .Y(_1336_)
);

NAND3X1 _4973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1333_),
    .C(_1336_),
    .Y(_1337_)
);

AOI21X1 _4974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(_1331_),
    .C(_1215_),
    .Y(_1338_)
);

NAND3X1 _4975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1336_),
    .C(_1216_),
    .Y(_1339_)
);

OAI21X1 _4976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(_1330_),
    .C(_1333_),
    .Y(_1340_)
);

AOI21X1 _4977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1339_),
    .B(_1340_),
    .C(_1213_),
    .Y(_1341_)
);

OAI21X1 _4978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1341_),
    .B(_1338_),
    .C(_1212_),
    .Y(_1342_)
);

NAND2X1 _4979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .B(_1185_),
    .Y(_1343_)
);

NAND3X1 _4980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_1339_),
    .C(_1340_),
    .Y(_1344_)
);

NOR3X1 _4981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1333_),
    .B(_1330_),
    .C(_1326_),
    .Y(_1345_)
);

AOI21X1 _4982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1336_),
    .C(_1216_),
    .Y(_1347_)
);

OAI21X1 _4983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1345_),
    .B(_1347_),
    .C(_1215_),
    .Y(_1348_)
);

NAND3X1 _4984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1344_),
    .B(_1343_),
    .C(_1348_),
    .Y(_1349_)
);

NAND3X1 _4985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1349_),
    .C(_1210_),
    .Y(_1350_)
);

AOI21X1 _4986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1189_),
    .B(_1191_),
    .C(_1197_),
    .Y(_1351_)
);

AOI21X1 _4987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1344_),
    .B(_1348_),
    .C(_1343_),
    .Y(_1352_)
);

NOR3X1 _4988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(_1212_),
    .C(_1341_),
    .Y(_1353_)
);

OAI21X1 _4989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1353_),
    .C(_1351_),
    .Y(_1354_)
);

NAND2X1 _4990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1354_),
    .Y(_1355_)
);

XNOR2X1 _4991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1209_),
    .B(_1355_),
    .Y(_1_[20])
);

INVX1 _4992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .Y(_1357_)
);

AOI21X1 _4993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(_1209_),
    .C(_1357_),
    .Y(_1358_)
);

OAI21X1 _4994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1347_),
    .B(_1215_),
    .C(_1339_),
    .Y(_1359_)
);

OAI21X1 _4995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1232_),
    .C(_1234_),
    .Y(_1360_)
);

OAI21X1 _4996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1239_),
    .C(_1329_),
    .Y(_1361_)
);

NAND2X1 _4997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1224_),
    .B(_1218_),
    .Y(_1362_)
);

INVX2 _4998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .Y(_1363_)
);

OAI21X1 _4999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2266_),
    .B(_2608_),
    .C(_1221_),
    .Y(_1364_)
);

OAI21X1 _5000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2266_),
    .B(_1221_),
    .C(_1364_),
    .Y(_1365_)
);

INVX1 _5001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .Y(_1366_)
);

OAI21X1 _5002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(_1363_),
    .C(_1366_),
    .Y(_1368_)
);

AOI21X1 _5003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .B(_1259_),
    .C(_1363_),
    .Y(_1369_)
);

NAND2X1 _5004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1369_),
    .Y(_1370_)
);

NAND3X1 _5005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1370_),
    .C(_1368_),
    .Y(_1371_)
);

INVX1 _5006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .Y(_1372_)
);

NAND2X1 _5007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1366_),
    .B(_1369_),
    .Y(_1373_)
);

OAI21X1 _5008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(_1363_),
    .C(_1365_),
    .Y(_1374_)
);

NAND3X1 _5009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1372_),
    .B(_1373_),
    .C(_1374_),
    .Y(_1375_)
);

NAND2X1 _5010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(_1375_),
    .Y(_1376_)
);

OAI21X1 _5011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(_1303_),
    .C(_1317_),
    .Y(_1377_)
);

OAI21X1 _5012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(_1244_),
    .C(_1248_),
    .Y(_1379_)
);

NAND2X1 _5013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_11_bF$buf2),
    .Y(_1380_)
);

NAND2X1 _5014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_14_bF$buf2),
    .Y(_1381_)
);

OAI21X1 _5015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2454_),
    .B(_2458_),
    .C(_881_),
    .Y(_1382_)
);

OAI21X1 _5016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1380_),
    .B(_1381_),
    .C(_1382_),
    .Y(_1383_)
);

OAI21X1 _5017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .B(_2781_),
    .C(_1383_),
    .Y(_1384_)
);

NAND2X1 _5018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_11_bF$buf1),
    .Y(_1385_)
);

OR2X2 _5019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_1385_),
    .Y(_1386_)
);

NAND3X1 _5020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1382_),
    .C(_1386_),
    .Y(_1387_)
);

NOR2X1 _5021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1271_),
    .B(_1272_),
    .Y(_1388_)
);

AOI21X1 _5022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1270_),
    .B(_1274_),
    .C(_1388_),
    .Y(_1389_)
);

INVX1 _5023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .Y(_1390_)
);

NAND3X1 _5024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .B(_1384_),
    .C(_1390_),
    .Y(_1391_)
);

AOI21X1 _5025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1382_),
    .B(_1386_),
    .C(_1220_),
    .Y(_1392_)
);

NOR2X1 _5026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .B(_1383_),
    .Y(_1393_)
);

OAI21X1 _5027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1393_),
    .B(_1392_),
    .C(_1389_),
    .Y(_1394_)
);

NAND3X1 _5028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1379_),
    .B(_1391_),
    .C(_1394_),
    .Y(_1395_)
);

INVX1 _5029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1379_),
    .Y(_1396_)
);

NAND3X1 _5030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .B(_1389_),
    .C(_1384_),
    .Y(_1397_)
);

OAI21X1 _5031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1393_),
    .B(_1392_),
    .C(_1390_),
    .Y(_1398_)
);

NAND3X1 _5032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1396_),
    .B(_1397_),
    .C(_1398_),
    .Y(_1401_)
);

AND2X2 _5033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .B(_1401_),
    .Y(_1402_)
);

AOI21X1 _5034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1276_),
    .C(_1299_),
    .Y(_1403_)
);

NAND2X1 _5035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_12_bF$buf1),
    .Y(_1404_)
);

OAI21X1 _5036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2614_),
    .B(_2527_),
    .C(_1272_),
    .Y(_1405_)
);

OAI21X1 _5037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(_1404_),
    .C(_1405_),
    .Y(_1406_)
);

XNOR2X1 _5038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1406_),
    .B(_708_),
    .Y(_1407_)
);

OAI21X1 _5039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1279_),
    .B(_1284_),
    .C(_1283_),
    .Y(_1408_)
);

NAND2X1 _5040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_13_bF$buf0),
    .Y(_1409_)
);

OAI21X1 _5041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_220_),
    .C(_1282_),
    .Y(_1410_)
);

INVX4 _5042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf1),
    .Y(_1412_)
);

AND2X2 _5043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_14_bF$buf0),
    .Y(_1413_)
);

OAI21X1 _5044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_1412_),
    .C(_1413_),
    .Y(_1414_)
);

AOI21X1 _5045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1410_),
    .B(_1414_),
    .C(_1409_),
    .Y(_1415_)
);

INVX2 _5046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1409_),
    .Y(_1416_)
);

NAND2X1 _5047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1282_),
    .B(_1413_),
    .Y(_1417_)
);

OAI21X1 _5048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_220_),
    .C(_1287_),
    .Y(_1418_)
);

AOI21X1 _5049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1418_),
    .B(_1417_),
    .C(_1416_),
    .Y(_1419_)
);

OAI21X1 _5050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1419_),
    .C(_1408_),
    .Y(_1420_)
);

AOI21X1 _5051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1285_),
    .C(_1288_),
    .Y(_1421_)
);

NAND3X1 _5052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1418_),
    .C(_1417_),
    .Y(_1423_)
);

NAND2X1 _5053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_14_bF$buf3),
    .Y(_1424_)
);

NOR2X1 _5054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1287_),
    .B(_1424_),
    .Y(_1425_)
);

NOR2X1 _5055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1282_),
    .B(_1413_),
    .Y(_1426_)
);

OAI21X1 _5056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1425_),
    .C(_1409_),
    .Y(_1427_)
);

NAND3X1 _5057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1421_),
    .B(_1423_),
    .C(_1427_),
    .Y(_1428_)
);

AOI21X1 _5058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1428_),
    .C(_1407_),
    .Y(_1429_)
);

INVX2 _5059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .Y(_1430_)
);

XNOR2X1 _5060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1406_),
    .B(_1430_),
    .Y(_1431_)
);

NAND3X1 _5061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1423_),
    .C(_1427_),
    .Y(_1432_)
);

OAI21X1 _5062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1419_),
    .C(_1421_),
    .Y(_1434_)
);

AOI21X1 _5063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1434_),
    .B(_1432_),
    .C(_1431_),
    .Y(_1435_)
);

OAI21X1 _5064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1429_),
    .B(_1435_),
    .C(_1403_),
    .Y(_1436_)
);

OAI21X1 _5065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1298_),
    .B(_1300_),
    .C(_1290_),
    .Y(_1437_)
);

NAND3X1 _5066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1432_),
    .B(_1434_),
    .C(_1431_),
    .Y(_1438_)
);

NAND3X1 _5067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1428_),
    .C(_1407_),
    .Y(_1439_)
);

NAND3X1 _5068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .B(_1438_),
    .C(_1437_),
    .Y(_1440_)
);

NAND3X1 _5069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(_1440_),
    .C(_1402_),
    .Y(_1441_)
);

NAND2X1 _5070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .B(_1401_),
    .Y(_1442_)
);

AOI21X1 _5071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .B(_1438_),
    .C(_1437_),
    .Y(_1443_)
);

NOR3X1 _5072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1429_),
    .B(_1435_),
    .C(_1403_),
    .Y(_1445_)
);

OAI21X1 _5073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1445_),
    .B(_1443_),
    .C(_1442_),
    .Y(_1446_)
);

NAND3X1 _5074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1377_),
    .B(_1446_),
    .C(_1441_),
    .Y(_1447_)
);

AOI21X1 _5075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1315_),
    .C(_1310_),
    .Y(_1448_)
);

NOR3X1 _5076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(_1443_),
    .C(_1445_),
    .Y(_1449_)
);

AOI21X1 _5077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(_1440_),
    .C(_1402_),
    .Y(_1450_)
);

OAI21X1 _5078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1450_),
    .C(_1448_),
    .Y(_1451_)
);

NAND3X1 _5079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1376_),
    .B(_1447_),
    .C(_1451_),
    .Y(_1452_)
);

AND2X2 _5080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(_1375_),
    .Y(_1453_)
);

OAI21X1 _5081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1450_),
    .C(_1377_),
    .Y(_1454_)
);

NAND3X1 _5082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1446_),
    .B(_1441_),
    .C(_1448_),
    .Y(_1456_)
);

NAND3X1 _5083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .B(_1454_),
    .C(_1453_),
    .Y(_1457_)
);

NAND3X1 _5084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1452_),
    .C(_1457_),
    .Y(_1458_)
);

AOI21X1 _5085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1328_),
    .B(_1327_),
    .C(_1325_),
    .Y(_1459_)
);

AOI21X1 _5086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .B(_1454_),
    .C(_1453_),
    .Y(_1460_)
);

AOI21X1 _5087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1447_),
    .B(_1451_),
    .C(_1376_),
    .Y(_1461_)
);

OAI21X1 _5088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1461_),
    .C(_1459_),
    .Y(_1462_)
);

NAND3X1 _5089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .B(_1458_),
    .C(_1462_),
    .Y(_1463_)
);

INVX2 _5090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .Y(_1464_)
);

NOR3X1 _5091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1461_),
    .C(_1459_),
    .Y(_1465_)
);

AOI21X1 _5092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(_1457_),
    .C(_1361_),
    .Y(_1467_)
);

OAI21X1 _5093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1465_),
    .B(_1467_),
    .C(_1464_),
    .Y(_1468_)
);

NAND3X1 _5094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1463_),
    .B(_1359_),
    .C(_1468_),
    .Y(_1469_)
);

AOI21X1 _5095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_1340_),
    .C(_1345_),
    .Y(_1470_)
);

OAI21X1 _5096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1461_),
    .C(_1361_),
    .Y(_1471_)
);

NAND3X1 _5097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(_1457_),
    .C(_1459_),
    .Y(_1472_)
);

AOI21X1 _5098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1471_),
    .B(_1472_),
    .C(_1464_),
    .Y(_1473_)
);

AOI21X1 _5099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1458_),
    .B(_1462_),
    .C(_1360_),
    .Y(_1474_)
);

OAI21X1 _5100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1474_),
    .C(_1470_),
    .Y(_1475_)
);

NAND3X1 _5101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1475_),
    .C(_1353_),
    .Y(_1476_)
);

OAI21X1 _5102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1474_),
    .C(_1359_),
    .Y(_1478_)
);

NAND3X1 _5103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1463_),
    .B(_1468_),
    .C(_1470_),
    .Y(_1479_)
);

NAND3X1 _5104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(_1479_),
    .C(_1349_),
    .Y(_1480_)
);

NAND2X1 _5105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(_1476_),
    .Y(_1481_)
);

INVX2 _5106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .Y(_1482_)
);

XNOR2X1 _5107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1482_),
    .Y(_1_[21])
);

OAI21X1 _5108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1350_),
    .C(_1476_),
    .Y(_1483_)
);

NOR2X1 _5109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1355_),
    .Y(_1484_)
);

AOI21X1 _5110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1484_),
    .B(_1209_),
    .C(_1483_),
    .Y(_1485_)
);

NOR2X1 _5111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(_1473_),
    .Y(_1486_)
);

OAI21X1 _5112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .B(_1464_),
    .C(_1458_),
    .Y(_1488_)
);

NAND3X1 _5113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1372_),
    .B(_1370_),
    .C(_1368_),
    .Y(_1489_)
);

OAI21X1 _5114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1369_),
    .C(_1489_),
    .Y(_1490_)
);

INVX2 _5115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .Y(_1491_)
);

AOI21X1 _5116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1446_),
    .B(_1441_),
    .C(_1377_),
    .Y(_1492_)
);

OAI21X1 _5117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .B(_1492_),
    .C(_1447_),
    .Y(_1493_)
);

NAND2X1 _5118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(_1222_),
    .Y(_1494_)
);

INVX2 _5119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1494_),
    .Y(_1495_)
);

NAND2X1 _5120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1391_),
    .B(_1395_),
    .Y(_1496_)
);

XNOR2X1 _5121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1495_),
    .Y(_1497_)
);

OAI21X1 _5122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1442_),
    .B(_1443_),
    .C(_1440_),
    .Y(_1499_)
);

OAI21X1 _5123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_1219_),
    .C(_1386_),
    .Y(_1500_)
);

NAND2X1 _5124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg[12]),
    .Y(_1501_)
);

NAND2X1 _5125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_14_bF$buf1),
    .Y(_1502_)
);

NOR2X1 _5126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .B(_1502_),
    .Y(_1503_)
);

AOI22X1 _5127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf0),
    .B(areg_14_bF$buf0),
    .C(breg_9_bF$buf3),
    .D(areg_13_bF$buf1),
    .Y(_1504_)
);

OAI21X1 _5128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .B(_1504_),
    .C(_1501_),
    .Y(_1505_)
);

INVX1 _5129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .Y(_1506_)
);

NOR2X1 _5130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1504_),
    .B(_1503_),
    .Y(_1507_)
);

NAND2X1 _5131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1506_),
    .B(_1507_),
    .Y(_1508_)
);

NOR2X1 _5132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(_1404_),
    .Y(_1510_)
);

AOI21X1 _5133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1430_),
    .B(_1405_),
    .C(_1510_),
    .Y(_1511_)
);

INVX1 _5134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .Y(_1512_)
);

NAND3X1 _5135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1505_),
    .B(_1512_),
    .C(_1508_),
    .Y(_1513_)
);

INVX1 _5136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1505_),
    .Y(_1514_)
);

AND2X2 _5137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1507_),
    .B(_1506_),
    .Y(_1515_)
);

OAI21X1 _5138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1514_),
    .C(_1511_),
    .Y(_1516_)
);

NAND3X1 _5139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .B(_1513_),
    .C(_1516_),
    .Y(_1517_)
);

INVX1 _5140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .Y(_1518_)
);

NAND3X1 _5141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(_1505_),
    .C(_1508_),
    .Y(_1519_)
);

OAI21X1 _5142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1514_),
    .C(_1512_),
    .Y(_1520_)
);

NAND3X1 _5143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1519_),
    .C(_1520_),
    .Y(_1521_)
);

NAND2X1 _5144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(_1521_),
    .Y(_1522_)
);

AOI21X1 _5145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1423_),
    .B(_1427_),
    .C(_1408_),
    .Y(_1523_)
);

OAI21X1 _5146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .B(_1523_),
    .C(_1432_),
    .Y(_1524_)
);

NAND2X1 _5147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf3),
    .B(areg_11_bF$buf0),
    .Y(_1525_)
);

NAND2X1 _5148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_15_bF$buf1),
    .Y(_1526_)
);

XOR2X1 _5149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1404_),
    .B(_1526_),
    .Y(_1527_)
);

XOR2X1 _5150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1525_),
    .Y(_1528_)
);

OAI21X1 _5151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1409_),
    .C(_1417_),
    .Y(_1529_)
);

NAND2X1 _5152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_13_bF$buf3),
    .Y(_1531_)
);

AND2X2 _5153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf1),
    .B(breg_15_bF$buf0),
    .Y(_1532_)
);

OAI21X1 _5154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_220_),
    .C(_1532_),
    .Y(_1533_)
);

AND2X2 _5155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_14_bF$buf2),
    .Y(_1534_)
);

OAI21X1 _5156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_1412_),
    .C(_1534_),
    .Y(_1535_)
);

AOI21X1 _5157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .B(_1535_),
    .C(_1531_),
    .Y(_1536_)
);

INVX2 _5158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1531_),
    .Y(_1537_)
);

NAND2X1 _5159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1532_),
    .B(_1534_),
    .Y(_1538_)
);

OAI22X1 _5160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_1412_),
    .C(_2116_),
    .D(_220_),
    .Y(_1539_)
);

AOI21X1 _5161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .B(_1538_),
    .C(_1537_),
    .Y(_1540_)
);

OAI21X1 _5162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1540_),
    .C(_1529_),
    .Y(_1542_)
);

AOI21X1 _5163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1418_),
    .C(_1425_),
    .Y(_1543_)
);

NAND3X1 _5164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(_1539_),
    .C(_1538_),
    .Y(_1544_)
);

AND2X2 _5165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1532_),
    .B(_1534_),
    .Y(_1545_)
);

NOR2X1 _5166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1532_),
    .B(_1534_),
    .Y(_1546_)
);

OAI21X1 _5167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1545_),
    .B(_1546_),
    .C(_1531_),
    .Y(_1547_)
);

NAND3X1 _5168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1543_),
    .B(_1544_),
    .C(_1547_),
    .Y(_1548_)
);

AOI21X1 _5169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1542_),
    .B(_1548_),
    .C(_1528_),
    .Y(_1549_)
);

XNOR2X1 _5170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1525_),
    .Y(_1550_)
);

NAND3X1 _5171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_1544_),
    .C(_1547_),
    .Y(_1551_)
);

OAI21X1 _5172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1540_),
    .C(_1543_),
    .Y(_1553_)
);

AOI21X1 _5173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(_1551_),
    .C(_1550_),
    .Y(_1554_)
);

OAI21X1 _5174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1554_),
    .C(_1524_),
    .Y(_1555_)
);

NOR3X1 _5175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(_1421_),
    .C(_1415_),
    .Y(_1556_)
);

AOI21X1 _5176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1434_),
    .B(_1431_),
    .C(_1556_),
    .Y(_1557_)
);

NAND3X1 _5177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1551_),
    .B(_1553_),
    .C(_1550_),
    .Y(_1558_)
);

NOR3X1 _5178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1540_),
    .B(_1543_),
    .C(_1536_),
    .Y(_1559_)
);

AOI21X1 _5179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1544_),
    .B(_1547_),
    .C(_1529_),
    .Y(_1560_)
);

OAI21X1 _5180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .B(_1559_),
    .C(_1528_),
    .Y(_1561_)
);

NAND3X1 _5181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1558_),
    .C(_1561_),
    .Y(_1562_)
);

AOI21X1 _5182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .B(_1555_),
    .C(_1522_),
    .Y(_1564_)
);

NAND3X1 _5183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1513_),
    .C(_1516_),
    .Y(_1565_)
);

NAND3X1 _5184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .B(_1519_),
    .C(_1520_),
    .Y(_1566_)
);

NAND2X1 _5185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1565_),
    .B(_1566_),
    .Y(_1567_)
);

NAND3X1 _5186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1524_),
    .B(_1558_),
    .C(_1561_),
    .Y(_1568_)
);

OAI21X1 _5187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1554_),
    .C(_1557_),
    .Y(_1569_)
);

AOI21X1 _5188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(_1569_),
    .C(_1567_),
    .Y(_1570_)
);

OAI21X1 _5189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1570_),
    .C(_1499_),
    .Y(_1571_)
);

AOI21X1 _5190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(_1402_),
    .C(_1445_),
    .Y(_1572_)
);

NAND3X1 _5191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1568_),
    .B(_1569_),
    .C(_1567_),
    .Y(_1573_)
);

NOR3X1 _5192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1557_),
    .C(_1549_),
    .Y(_1575_)
);

AOI21X1 _5193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1558_),
    .B(_1561_),
    .C(_1524_),
    .Y(_1576_)
);

OAI21X1 _5194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1575_),
    .B(_1576_),
    .C(_1522_),
    .Y(_1577_)
);

NAND3X1 _5195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1577_),
    .C(_1572_),
    .Y(_1578_)
);

AOI21X1 _5196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1571_),
    .B(_1578_),
    .C(_1497_),
    .Y(_1579_)
);

INVX2 _5197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .Y(_1580_)
);

NAND3X1 _5198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1499_),
    .B(_1573_),
    .C(_1577_),
    .Y(_1581_)
);

OAI21X1 _5199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1570_),
    .C(_1572_),
    .Y(_1582_)
);

AOI21X1 _5200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1581_),
    .B(_1582_),
    .C(_1580_),
    .Y(_1583_)
);

OAI21X1 _5201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1579_),
    .B(_1583_),
    .C(_1493_),
    .Y(_1584_)
);

NOR3X1 _5202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1450_),
    .C(_1449_),
    .Y(_1586_)
);

AOI21X1 _5203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1376_),
    .B(_1451_),
    .C(_1586_),
    .Y(_1587_)
);

NAND3X1 _5204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(_1581_),
    .C(_1582_),
    .Y(_1588_)
);

NAND3X1 _5205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .B(_1571_),
    .C(_1578_),
    .Y(_1589_)
);

NAND3X1 _5206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1589_),
    .C(_1587_),
    .Y(_1590_)
);

AOI21X1 _5207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .B(_1590_),
    .C(_1491_),
    .Y(_1591_)
);

NAND3X1 _5208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1589_),
    .C(_1493_),
    .Y(_1592_)
);

OAI21X1 _5209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1579_),
    .B(_1583_),
    .C(_1587_),
    .Y(_1593_)
);

AOI21X1 _5210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1593_),
    .C(_1490_),
    .Y(_1594_)
);

OAI21X1 _5211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .C(_1488_),
    .Y(_1595_)
);

AOI21X1 _5212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .B(_1462_),
    .C(_1465_),
    .Y(_1597_)
);

NAND3X1 _5213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1592_),
    .C(_1593_),
    .Y(_1598_)
);

NAND3X1 _5214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1491_),
    .B(_1584_),
    .C(_1590_),
    .Y(_1599_)
);

NAND3X1 _5215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1600_)
);

AOI22X1 _5216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1486_),
    .C(_1600_),
    .D(_1595_),
    .Y(_1601_)
);

INVX1 _5217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1601_),
    .Y(_1602_)
);

NAND3X1 _5218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_1488_),
    .C(_1599_),
    .Y(_1603_)
);

OAI21X1 _5219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .C(_1597_),
    .Y(_1604_)
);

AOI21X1 _5220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1604_),
    .C(_1469_),
    .Y(_1605_)
);

INVX1 _5221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1605_),
    .Y(_1606_)
);

NAND2X1 _5222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(_1602_),
    .Y(_1608_)
);

XNOR2X1 _5223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1608_),
    .Y(_1_[22])
);

AOI21X1 _5224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1595_),
    .B(_1600_),
    .C(_1469_),
    .Y(_1609_)
);

INVX1 _5225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1609_),
    .Y(_1610_)
);

NOR2X1 _5226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1605_),
    .B(_1601_),
    .Y(_1611_)
);

OAI21X1 _5227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1611_),
    .C(_1610_),
    .Y(_1612_)
);

NOR3X1 _5228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .C(_1597_),
    .Y(_1613_)
);

AOI21X1 _5229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1589_),
    .C(_1493_),
    .Y(_1614_)
);

OAI21X1 _5230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1614_),
    .B(_1491_),
    .C(_1592_),
    .Y(_1615_)
);

NAND2X1 _5231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1495_),
    .B(_1496_),
    .Y(_1616_)
);

AOI21X1 _5232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1577_),
    .C(_1499_),
    .Y(_1618_)
);

OAI21X1 _5233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1497_),
    .C(_1581_),
    .Y(_1619_)
);

NAND2X1 _5234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1517_),
    .Y(_1620_)
);

INVX1 _5235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .Y(_1621_)
);

OAI21X1 _5236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1522_),
    .B(_1576_),
    .C(_1568_),
    .Y(_1622_)
);

OAI21X1 _5237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .B(_1502_),
    .C(_1508_),
    .Y(_1623_)
);

AOI22X1 _5238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf3),
    .B(areg_13_bF$buf0),
    .C(breg_11_bF$buf2),
    .D(areg[12]),
    .Y(_1624_)
);

NAND2X1 _5239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf1),
    .B(areg_13_bF$buf3),
    .Y(_1625_)
);

NOR2X1 _5240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1625_),
    .Y(_1626_)
);

NOR2X1 _5241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .B(_1626_),
    .Y(_1627_)
);

NAND2X1 _5242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_15_bF$buf0),
    .Y(_1629_)
);

AND2X2 _5243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1404_),
    .B(_1526_),
    .Y(_1630_)
);

OAI22X1 _5244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_1629_),
    .C(_1630_),
    .D(_1525_),
    .Y(_1631_)
);

NAND2X1 _5245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1631_),
    .Y(_1632_)
);

NOR2X1 _5246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1631_),
    .Y(_1633_)
);

INVX1 _5247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1633_),
    .Y(_1634_)
);

NAND3X1 _5248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1623_),
    .B(_1632_),
    .C(_1634_),
    .Y(_1635_)
);

NOR2X1 _5249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .B(_1515_),
    .Y(_1636_)
);

INVX1 _5250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1632_),
    .Y(_1637_)
);

OAI21X1 _5251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(_1633_),
    .C(_1636_),
    .Y(_1638_)
);

AND2X2 _5252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1635_),
    .B(_1638_),
    .Y(_1640_)
);

AOI21X1 _5253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1553_),
    .B(_1550_),
    .C(_1559_),
    .Y(_1641_)
);

INVX1 _5254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1629_),
    .Y(_1642_)
);

AOI22X1 _5255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_8_bF$buf3),
    .B(areg_15_bF$buf3),
    .C(areg_11_bF$buf3),
    .D(breg_12_bF$buf3),
    .Y(_1643_)
);

AOI21X1 _5256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1095_),
    .B(_1642_),
    .C(_1643_),
    .Y(_1644_)
);

XOR2X1 _5257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1644_),
    .B(_1502_),
    .Y(_1645_)
);

OAI21X1 _5258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1546_),
    .B(_1531_),
    .C(_1538_),
    .Y(_1646_)
);

NAND2X1 _5259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf0),
    .B(breg_13_bF$buf2),
    .Y(_1647_)
);

AND2X2 _5260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_15_bF$buf3),
    .Y(_1648_)
);

OAI21X1 _5261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2342_),
    .B(_220_),
    .C(_1648_),
    .Y(_1649_)
);

AND2X2 _5262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_14_bF$buf1),
    .Y(_1651_)
);

OAI21X1 _5263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_1412_),
    .C(_1651_),
    .Y(_1652_)
);

AOI21X1 _5264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .B(_1652_),
    .C(_1647_),
    .Y(_1653_)
);

INVX1 _5265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .Y(_1654_)
);

NAND2X1 _5266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1648_),
    .B(_1651_),
    .Y(_1655_)
);

NAND2X1 _5267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_14_bF$buf0),
    .Y(_1656_)
);

OAI21X1 _5268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2116_),
    .B(_1412_),
    .C(_1656_),
    .Y(_1657_)
);

AOI21X1 _5269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1655_),
    .C(_1654_),
    .Y(_1658_)
);

OAI21X1 _5270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(_1658_),
    .C(_1646_),
    .Y(_1659_)
);

AOI21X1 _5271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(_1539_),
    .C(_1545_),
    .Y(_1660_)
);

NAND3X1 _5272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1654_),
    .B(_1657_),
    .C(_1655_),
    .Y(_1662_)
);

NAND3X1 _5273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(_1649_),
    .C(_1652_),
    .Y(_1663_)
);

NAND3X1 _5274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1662_),
    .B(_1663_),
    .C(_1660_),
    .Y(_1664_)
);

AOI21X1 _5275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1664_),
    .C(_1645_),
    .Y(_1665_)
);

XNOR2X1 _5276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1644_),
    .B(_1502_),
    .Y(_1666_)
);

NAND3X1 _5277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1662_),
    .B(_1663_),
    .C(_1646_),
    .Y(_1667_)
);

OAI21X1 _5278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(_1658_),
    .C(_1660_),
    .Y(_1668_)
);

AOI21X1 _5279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1668_),
    .B(_1667_),
    .C(_1666_),
    .Y(_1669_)
);

OAI21X1 _5280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .B(_1669_),
    .C(_1641_),
    .Y(_1670_)
);

OAI21X1 _5281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1560_),
    .C(_1551_),
    .Y(_1671_)
);

NAND3X1 _5282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1668_),
    .B(_1667_),
    .C(_1666_),
    .Y(_1673_)
);

NAND3X1 _5283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1664_),
    .C(_1645_),
    .Y(_1674_)
);

NAND3X1 _5284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1674_),
    .C(_1671_),
    .Y(_1675_)
);

AOI21X1 _5285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1670_),
    .B(_1675_),
    .C(_1640_),
    .Y(_1676_)
);

NAND2X1 _5286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1638_),
    .B(_1635_),
    .Y(_1677_)
);

AOI21X1 _5287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1674_),
    .C(_1671_),
    .Y(_1678_)
);

NOR3X1 _5288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .B(_1669_),
    .C(_1641_),
    .Y(_1679_)
);

NOR3X1 _5289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(_1678_),
    .C(_1679_),
    .Y(_1680_)
);

OAI21X1 _5290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1680_),
    .B(_1676_),
    .C(_1622_),
    .Y(_1681_)
);

AOI21X1 _5291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1569_),
    .B(_1567_),
    .C(_1575_),
    .Y(_1682_)
);

OAI21X1 _5292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1679_),
    .B(_1678_),
    .C(_1677_),
    .Y(_1684_)
);

NAND3X1 _5293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1670_),
    .B(_1675_),
    .C(_1640_),
    .Y(_1685_)
);

NAND3X1 _5294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1684_),
    .B(_1685_),
    .C(_1682_),
    .Y(_1686_)
);

AOI21X1 _5295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_),
    .B(_1681_),
    .C(_1621_),
    .Y(_1687_)
);

NAND3X1 _5296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1684_),
    .B(_1685_),
    .C(_1622_),
    .Y(_1688_)
);

OAI21X1 _5297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1680_),
    .B(_1676_),
    .C(_1682_),
    .Y(_1689_)
);

AOI21X1 _5298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1688_),
    .B(_1689_),
    .C(_1620_),
    .Y(_1690_)
);

OAI21X1 _5299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .B(_1690_),
    .C(_1619_),
    .Y(_1691_)
);

NOR3X1 _5300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1570_),
    .C(_1572_),
    .Y(_1692_)
);

AOI21X1 _5301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(_1582_),
    .C(_1692_),
    .Y(_1693_)
);

NAND3X1 _5302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(_1688_),
    .C(_1689_),
    .Y(_1695_)
);

NAND3X1 _5303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1621_),
    .B(_1686_),
    .C(_1681_),
    .Y(_1696_)
);

NAND3X1 _5304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(_1696_),
    .C(_1693_),
    .Y(_1697_)
);

AOI21X1 _5305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1697_),
    .B(_1691_),
    .C(_1616_),
    .Y(_1698_)
);

INVX1 _5306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .Y(_1699_)
);

NAND3X1 _5307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1619_),
    .B(_1695_),
    .C(_1696_),
    .Y(_1700_)
);

OAI21X1 _5308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .B(_1690_),
    .C(_1693_),
    .Y(_1701_)
);

AOI21X1 _5309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1700_),
    .B(_1701_),
    .C(_1699_),
    .Y(_1702_)
);

OAI21X1 _5310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .B(_1702_),
    .C(_1615_),
    .Y(_1703_)
);

NOR3X1 _5311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1579_),
    .B(_1583_),
    .C(_1587_),
    .Y(_1704_)
);

AOI21X1 _5312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1593_),
    .C(_1704_),
    .Y(_1706_)
);

NAND3X1 _5313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1699_),
    .B(_1700_),
    .C(_1701_),
    .Y(_1707_)
);

NAND3X1 _5314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(_1697_),
    .C(_1691_),
    .Y(_1708_)
);

NAND3X1 _5315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1707_),
    .B(_1708_),
    .C(_1706_),
    .Y(_1709_)
);

AOI21X1 _5316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1703_),
    .B(_1709_),
    .C(_1613_),
    .Y(_1710_)
);

NAND3X1 _5317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1615_),
    .B(_1707_),
    .C(_1708_),
    .Y(_1711_)
);

OAI21X1 _5318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .B(_1702_),
    .C(_1706_),
    .Y(_1712_)
);

AOI21X1 _5319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1711_),
    .B(_1712_),
    .C(_1603_),
    .Y(_1713_)
);

NOR2X1 _5320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1713_),
    .B(_1710_),
    .Y(_1714_)
);

XNOR2X1 _5321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1714_),
    .Y(_1_[23])
);

INVX1 _5322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1711_),
    .Y(_1715_)
);

NAND2X1 _5323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1700_),
    .B(_1707_),
    .Y(_1716_)
);

NAND2X1 _5324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1688_),
    .B(_1695_),
    .Y(_1717_)
);

INVX1 _5325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1717_),
    .Y(_1718_)
);

OAI21X1 _5326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1636_),
    .B(_1633_),
    .C(_1632_),
    .Y(_1719_)
);

OAI21X1 _5327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(_1678_),
    .C(_1675_),
    .Y(_1720_)
);

INVX1 _5328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1720_),
    .Y(_1721_)
);

INVX2 _5329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1626_),
    .Y(_1722_)
);

OAI22X1 _5330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1629_),
    .C(_1643_),
    .D(_1502_),
    .Y(_1723_)
);

NOR2X1 _5331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2773_),
    .B(_1723_),
    .Y(_1724_)
);

NAND2X1 _5332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2773_),
    .B(_1723_),
    .Y(_1726_)
);

INVX1 _5333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .Y(_1727_)
);

NOR2X1 _5334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1727_),
    .Y(_1728_)
);

XNOR2X1 _5335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1728_),
    .B(_1722_),
    .Y(_1729_)
);

AND2X2 _5336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1667_),
    .Y(_1730_)
);

NAND2X1 _5337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_14_bF$buf3),
    .Y(_1731_)
);

NOR2X1 _5338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1731_),
    .Y(_1732_)
);

AOI22X1 _5339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_14_bF$buf2),
    .C(areg_11_bF$buf2),
    .D(breg_13_bF$buf0),
    .Y(_1733_)
);

OAI21X1 _5340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1732_),
    .B(_1733_),
    .C(_1625_),
    .Y(_1734_)
);

NOR2X1 _5341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1733_),
    .B(_1732_),
    .Y(_1735_)
);

NAND3X1 _5342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_13_bF$buf2),
    .C(_1735_),
    .Y(_1738_)
);

AND2X2 _5343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1734_),
    .Y(_1739_)
);

INVX1 _5344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1648_),
    .Y(_1740_)
);

OAI21X1 _5345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1740_),
    .B(_1656_),
    .C(_1662_),
    .Y(_1741_)
);

NAND2X1 _5346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_15_bF$buf2),
    .Y(_1742_)
);

NAND2X1 _5347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .B(breg_15_bF$buf1),
    .Y(_1743_)
);

OAI21X1 _5348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2614_),
    .B(_220_),
    .C(_1743_),
    .Y(_1744_)
);

OAI21X1 _5349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1656_),
    .B(_1742_),
    .C(_1744_),
    .Y(_1745_)
);

XNOR2X1 _5350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1745_),
    .B(_1090_),
    .Y(_1746_)
);

XNOR2X1 _5351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1746_),
    .B(_1741_),
    .Y(_1747_)
);

XNOR2X1 _5352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1747_),
    .B(_1739_),
    .Y(_1749_)
);

XOR2X1 _5353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1749_),
    .B(_1730_),
    .Y(_1750_)
);

XNOR2X1 _5354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1750_),
    .B(_1729_),
    .Y(_1751_)
);

NAND2X1 _5355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1721_),
    .B(_1751_),
    .Y(_1752_)
);

OR2X2 _5356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1751_),
    .B(_1721_),
    .Y(_1753_)
);

AOI21X1 _5357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1752_),
    .B(_1753_),
    .C(_1719_),
    .Y(_1754_)
);

INVX2 _5358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1719_),
    .Y(_1755_)
);

OR2X2 _5359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1750_),
    .B(_1729_),
    .Y(_1756_)
);

NAND2X1 _5360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1729_),
    .B(_1750_),
    .Y(_1757_)
);

AOI21X1 _5361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1757_),
    .B(_1756_),
    .C(_1720_),
    .Y(_1758_)
);

NOR2X1 _5362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1721_),
    .B(_1751_),
    .Y(_1760_)
);

NOR3X1 _5363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1758_),
    .B(_1755_),
    .C(_1760_),
    .Y(_1761_)
);

OAI21X1 _5364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(_1761_),
    .C(_1718_),
    .Y(_1762_)
);

OAI21X1 _5365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1760_),
    .B(_1758_),
    .C(_1755_),
    .Y(_1763_)
);

NAND3X1 _5366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1719_),
    .B(_1752_),
    .C(_1753_),
    .Y(_1764_)
);

NAND3X1 _5367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1763_),
    .B(_1717_),
    .C(_1764_),
    .Y(_1765_)
);

NAND3X1 _5368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1716_),
    .B(_1765_),
    .C(_1762_),
    .Y(_1766_)
);

AOI21X1 _5369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .B(_1762_),
    .C(_1716_),
    .Y(_1767_)
);

INVX1 _5370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .Y(_1768_)
);

NAND3X1 _5371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1715_),
    .B(_1766_),
    .C(_1768_),
    .Y(_1769_)
);

INVX1 _5372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1766_),
    .Y(_1771_)
);

OAI21X1 _5373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1771_),
    .B(_1767_),
    .C(_1711_),
    .Y(_1772_)
);

AND2X2 _5374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1769_),
    .B(_1772_),
    .Y(_1773_)
);

OAI22X1 _5375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1601_),
    .B(_1605_),
    .C(_1710_),
    .D(_1713_),
    .Y(_1774_)
);

INVX1 _5376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1774_),
    .Y(_1775_)
);

NAND2X1 _5377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1711_),
    .B(_1712_),
    .Y(_1776_)
);

OAI21X1 _5378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1710_),
    .B(_1713_),
    .C(_1609_),
    .Y(_1777_)
);

OAI21X1 _5379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1776_),
    .C(_1777_),
    .Y(_1778_)
);

AOI21X1 _5380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1775_),
    .B(_1483_),
    .C(_1778_),
    .Y(_1779_)
);

AND2X2 _5381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(_1350_),
    .Y(_1780_)
);

NAND3X1 _5382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1780_),
    .B(_1482_),
    .C(_1775_),
    .Y(_1782_)
);

OAI21X1 _5383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1207_),
    .B(_1782_),
    .C(_1779_),
    .Y(_1783_)
);

NOR3X1 _5384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_298_),
    .C(_485_),
    .Y(_1784_)
);

OAI21X1 _5385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_296_),
    .C(_487_),
    .Y(_1785_)
);

AOI21X1 _5386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1784_),
    .B(_124_),
    .C(_1785_),
    .Y(_1786_)
);

NAND3X1 _5387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_125_),
    .B(_1784_),
    .C(_2596_),
    .Y(_1787_)
);

NOR3X1 _5388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1481_),
    .B(_1774_),
    .C(_1355_),
    .Y(_1788_)
);

NAND3X1 _5389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .B(_1202_),
    .C(_1788_),
    .Y(_1789_)
);

AOI21X1 _5390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .B(_1787_),
    .C(_1789_),
    .Y(_1790_)
);

NOR2X1 _5391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1783_),
    .B(_1790_),
    .Y(_1791_)
);

XNOR2X1 _5392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1791_),
    .B(_1773_),
    .Y(_1_[24])
);

NAND2X1 _5393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1772_),
    .B(_1769_),
    .Y(_1793_)
);

OAI21X1 _5394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1791_),
    .B(_1793_),
    .C(_1769_),
    .Y(_1794_)
);

OAI21X1 _5395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1758_),
    .B(_1755_),
    .C(_1753_),
    .Y(_1795_)
);

OAI21X1 _5396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1722_),
    .C(_1726_),
    .Y(_1796_)
);

INVX1 _5397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1796_),
    .Y(_1797_)
);

OAI21X1 _5398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1730_),
    .B(_1749_),
    .C(_1757_),
    .Y(_1798_)
);

OAI21X1 _5399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1731_),
    .C(_1738_),
    .Y(_1799_)
);

INVX1 _5400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .Y(_1800_)
);

INVX1 _5401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1741_),
    .Y(_1801_)
);

NOR2X1 _5402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1746_),
    .B(_1801_),
    .Y(_1803_)
);

AOI21X1 _5403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1739_),
    .B(_1747_),
    .C(_1803_),
    .Y(_1804_)
);

INVX1 _5404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1804_),
    .Y(_1805_)
);

NAND2X1 _5405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .B(breg_13_bF$buf3),
    .Y(_1806_)
);

NAND2X1 _5406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_14_bF$buf1),
    .Y(_1807_)
);

NOR2X1 _5407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1625_),
    .B(_1807_),
    .Y(_1808_)
);

AOI22X1 _5408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf3),
    .B(areg_14_bF$buf0),
    .C(breg_12_bF$buf1),
    .D(areg_13_bF$buf1),
    .Y(_1809_)
);

OAI21X1 _5409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1808_),
    .B(_1809_),
    .C(_1806_),
    .Y(_1810_)
);

NOR2X1 _5410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1808_),
    .Y(_1811_)
);

NAND3X1 _5411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .B(breg_13_bF$buf2),
    .C(_1811_),
    .Y(_1812_)
);

AND2X2 _5412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1812_),
    .B(_1810_),
    .Y(_1814_)
);

OAI22X1 _5413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1656_),
    .B(_1742_),
    .C(_1745_),
    .D(_1090_),
    .Y(_1815_)
);

NOR2X1 _5414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2458_),
    .B(_220_),
    .Y(_1816_)
);

NAND2X1 _5415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_15_bF$buf2),
    .Y(_1817_)
);

OAI21X1 _5416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2454_),
    .B(_528_),
    .C(_1742_),
    .Y(_1818_)
);

OAI21X1 _5417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1268_),
    .B(_1817_),
    .C(_1818_),
    .Y(_1819_)
);

XNOR2X1 _5418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1819_),
    .B(_1816_),
    .Y(_1820_)
);

XOR2X1 _5419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1820_),
    .B(_1815_),
    .Y(_1821_)
);

XOR2X1 _5420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1821_),
    .B(_1814_),
    .Y(_1822_)
);

NOR2X1 _5421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .B(_1805_),
    .Y(_1823_)
);

XNOR2X1 _5422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1821_),
    .B(_1814_),
    .Y(_1825_)
);

NOR2X1 _5423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1804_),
    .B(_1825_),
    .Y(_1826_)
);

OAI21X1 _5424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_1826_),
    .C(_1800_),
    .Y(_1827_)
);

XOR2X1 _5425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1804_),
    .Y(_1828_)
);

NAND2X1 _5426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(_1828_),
    .Y(_1829_)
);

AOI21X1 _5427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1829_),
    .C(_1798_),
    .Y(_1830_)
);

NOR2X1 _5428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1730_),
    .B(_1749_),
    .Y(_1831_)
);

AOI21X1 _5429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1729_),
    .B(_1750_),
    .C(_1831_),
    .Y(_1832_)
);

NAND2X1 _5430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1829_),
    .Y(_1833_)
);

NOR2X1 _5431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(_1833_),
    .Y(_1834_)
);

OAI21X1 _5432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1830_),
    .B(_1834_),
    .C(_1797_),
    .Y(_1836_)
);

NAND2X1 _5433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(_1833_),
    .Y(_1837_)
);

NAND3X1 _5434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1829_),
    .C(_1798_),
    .Y(_1838_)
);

NAND3X1 _5435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1796_),
    .B(_1837_),
    .C(_1838_),
    .Y(_1839_)
);

AOI21X1 _5436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1839_),
    .B(_1836_),
    .C(_1795_),
    .Y(_1840_)
);

NAND3X1 _5437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1839_),
    .B(_1795_),
    .C(_1836_),
    .Y(_1841_)
);

INVX2 _5438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .Y(_1842_)
);

OAI21X1 _5439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(_1840_),
    .C(_1765_),
    .Y(_1843_)
);

INVX1 _5440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .Y(_1844_)
);

INVX1 _5441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .Y(_1845_)
);

NAND3X1 _5442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1845_),
    .C(_1844_),
    .Y(_1847_)
);

NAND3X1 _5443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1843_),
    .B(_1847_),
    .C(_1771_),
    .Y(_1848_)
);

AOI21X1 _5444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1845_),
    .C(_1844_),
    .Y(_1849_)
);

NOR3X1 _5445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .B(_1840_),
    .C(_1842_),
    .Y(_1850_)
);

OAI21X1 _5446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1850_),
    .B(_1849_),
    .C(_1766_),
    .Y(_1851_)
);

NAND2X1 _5447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(_1851_),
    .Y(_1852_)
);

XNOR2X1 _5448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1794_),
    .B(_1852_),
    .Y(_1_[25])
);

NAND2X1 _5449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(_1769_),
    .Y(_1853_)
);

NAND2X1 _5450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1851_),
    .B(_1853_),
    .Y(_1854_)
);

NOR2X1 _5451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_1793_),
    .Y(_1855_)
);

OAI21X1 _5452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1790_),
    .B(_1783_),
    .C(_1855_),
    .Y(_1857_)
);

INVX1 _5453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1795_),
    .Y(_1858_)
);

NAND2X1 _5454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1839_),
    .B(_1836_),
    .Y(_1859_)
);

OAI21X1 _5455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1830_),
    .B(_1797_),
    .C(_1838_),
    .Y(_1860_)
);

AOI21X1 _5456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(_1828_),
    .C(_1826_),
    .Y(_1861_)
);

OAI21X1 _5457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1625_),
    .B(_1807_),
    .C(_1812_),
    .Y(_1862_)
);

NAND2X1 _5458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_1820_),
    .Y(_1863_)
);

NAND2X1 _5459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1814_),
    .B(_1821_),
    .Y(_1864_)
);

NAND2X1 _5460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1863_),
    .B(_1864_),
    .Y(_1865_)
);

NAND2X1 _5461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf0),
    .B(breg_14_bF$buf3),
    .Y(_1866_)
);

NOR2X1 _5462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1866_),
    .Y(_1868_)
);

AOI22X1 _5463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .B(breg_14_bF$buf2),
    .C(breg_13_bF$buf1),
    .D(areg_13_bF$buf3),
    .Y(_1869_)
);

NOR2X1 _5464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1869_),
    .B(_1868_),
    .Y(_1870_)
);

INVX2 _5465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .Y(_1871_)
);

AOI22X1 _5466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1270_),
    .B(_1871_),
    .C(_1818_),
    .D(_1816_),
    .Y(_1872_)
);

OAI22X1 _5467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .B(_528_),
    .C(_2458_),
    .D(_1412_),
    .Y(_1873_)
);

OAI21X1 _5468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(_1817_),
    .C(_1873_),
    .Y(_1874_)
);

XNOR2X1 _5469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1874_),
    .B(_1807_),
    .Y(_1875_)
);

XNOR2X1 _5470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1875_),
    .B(_1872_),
    .Y(_1876_)
);

XNOR2X1 _5471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(_1870_),
    .Y(_1877_)
);

XOR2X1 _5472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1877_),
    .B(_1865_),
    .Y(_1879_)
);

NOR2X1 _5473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .B(_1879_),
    .Y(_1880_)
);

AND2X2 _5474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1879_),
    .B(_1862_),
    .Y(_1881_)
);

OAI21X1 _5475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1881_),
    .B(_1880_),
    .C(_1861_),
    .Y(_1882_)
);

INVX1 _5476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .Y(_1883_)
);

OAI21X1 _5477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1823_),
    .B(_1800_),
    .C(_1883_),
    .Y(_1884_)
);

INVX1 _5478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .Y(_1885_)
);

NOR2X1 _5479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1865_),
    .B(_1877_),
    .Y(_1886_)
);

NAND2X1 _5480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1865_),
    .B(_1877_),
    .Y(_1887_)
);

INVX1 _5481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1887_),
    .Y(_1888_)
);

OAI21X1 _5482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1888_),
    .B(_1886_),
    .C(_1885_),
    .Y(_1890_)
);

NAND2X1 _5483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .B(_1879_),
    .Y(_1891_)
);

NAND3X1 _5484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1890_),
    .C(_1891_),
    .Y(_1892_)
);

NAND2X1 _5485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1892_),
    .B(_1882_),
    .Y(_1893_)
);

NAND2X1 _5486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1860_),
    .Y(_1894_)
);

AOI21X1 _5487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1796_),
    .B(_1837_),
    .C(_1834_),
    .Y(_1895_)
);

AND2X2 _5488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1882_),
    .B(_1892_),
    .Y(_1896_)
);

NAND2X1 _5489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .B(_1895_),
    .Y(_1897_)
);

NAND2X1 _5490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1897_),
    .B(_1894_),
    .Y(_1898_)
);

OAI21X1 _5491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(_1859_),
    .C(_1898_),
    .Y(_1899_)
);

NAND2X1 _5492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .B(_1860_),
    .Y(_1901_)
);

NAND2X1 _5493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1895_),
    .Y(_1902_)
);

NAND2X1 _5494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1902_),
    .B(_1901_),
    .Y(_1903_)
);

NAND2X1 _5495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1903_),
    .B(_1842_),
    .Y(_1904_)
);

AOI21X1 _5496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1904_),
    .B(_1899_),
    .C(_1850_),
    .Y(_1905_)
);

NAND2X1 _5497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1898_),
    .B(_1842_),
    .Y(_1906_)
);

OAI21X1 _5498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(_1859_),
    .C(_1903_),
    .Y(_1907_)
);

AOI21X1 _5499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(_1906_),
    .C(_1847_),
    .Y(_1908_)
);

NOR2X1 _5500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1908_),
    .B(_1905_),
    .Y(_1909_)
);

AOI21X1 _5501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1854_),
    .B(_1857_),
    .C(_1909_),
    .Y(_1910_)
);

AND2X2 _5502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1851_),
    .B(_1848_),
    .Y(_1912_)
);

NAND2X1 _5503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1912_),
    .B(_1773_),
    .Y(_1913_)
);

OAI21X1 _5504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1791_),
    .B(_1913_),
    .C(_1854_),
    .Y(_1914_)
);

INVX1 _5505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1909_),
    .Y(_1915_)
);

NOR2X1 _5506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1915_),
    .B(_1914_),
    .Y(_1916_)
);

NOR2X1 _5507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(_1916_),
    .Y(_1_[26])
);

NAND2X1 _5508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(_1906_),
    .Y(_1917_)
);

NOR2X1 _5509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1847_),
    .B(_1917_),
    .Y(_1918_)
);

NOR2X1 _5510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1895_),
    .Y(_1919_)
);

OAI21X1 _5511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1886_),
    .B(_1885_),
    .C(_1887_),
    .Y(_1920_)
);

NOR2X1 _5512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_1875_),
    .Y(_1922_)
);

INVX1 _5513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .Y(_1923_)
);

NOR2X1 _5514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .B(_1876_),
    .Y(_1924_)
);

NOR2X1 _5515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1922_),
    .B(_1924_),
    .Y(_1925_)
);

NOR2X1 _5516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2608_),
    .B(_1412_),
    .Y(_1926_)
);

OAI22X1 _5517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(_1817_),
    .C(_1874_),
    .D(_1807_),
    .Y(_1927_)
);

NAND2X1 _5518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf0),
    .B(areg_15_bF$buf1),
    .Y(_1928_)
);

OAI21X1 _5519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .B(_528_),
    .C(_1731_),
    .Y(_1929_)
);

OAI21X1 _5520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(_1928_),
    .C(_1929_),
    .Y(_1930_)
);

XNOR2X1 _5521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1866_),
    .Y(_1931_)
);

XNOR2X1 _5522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1931_),
    .B(_1927_),
    .Y(_1933_)
);

XNOR2X1 _5523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1933_),
    .B(_1926_),
    .Y(_1934_)
);

XOR2X1 _5524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(_1934_),
    .Y(_1935_)
);

NAND2X1 _5525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(_1935_),
    .Y(_1936_)
);

XNOR2X1 _5526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(_1934_),
    .Y(_1937_)
);

OAI21X1 _5527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1866_),
    .C(_1937_),
    .Y(_1938_)
);

NAND3X1 _5528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1920_),
    .B(_1936_),
    .C(_1938_),
    .Y(_1939_)
);

INVX1 _5529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1920_),
    .Y(_1940_)
);

OAI21X1 _5530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1866_),
    .C(_1935_),
    .Y(_1941_)
);

NAND2X1 _5531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(_1937_),
    .Y(_1942_)
);

NAND3X1 _5532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1940_),
    .B(_1942_),
    .C(_1941_),
    .Y(_1944_)
);

NAND2X1 _5533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1944_),
    .Y(_1945_)
);

NAND2X1 _5534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1892_),
    .B(_1945_),
    .Y(_1946_)
);

INVX1 _5535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1892_),
    .Y(_1947_)
);

NAND3X1 _5536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1944_),
    .C(_1947_),
    .Y(_1948_)
);

AOI21X1 _5537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1946_),
    .B(_1948_),
    .C(_1919_),
    .Y(_1949_)
);

NAND2X1 _5538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_1946_),
    .Y(_1950_)
);

NOR2X1 _5539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1950_),
    .Y(_1951_)
);

OAI22X1 _5540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1903_),
    .C(_1951_),
    .D(_1949_),
    .Y(_1952_)
);

AOI21X1 _5541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1894_),
    .B(_1897_),
    .C(_1841_),
    .Y(_1953_)
);

OAI21X1 _5542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1895_),
    .B(_1893_),
    .C(_1950_),
    .Y(_1955_)
);

NAND3X1 _5543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1946_),
    .B(_1948_),
    .C(_1919_),
    .Y(_1956_)
);

NAND3X1 _5544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1955_),
    .B(_1956_),
    .C(_1953_),
    .Y(_1957_)
);

NAND2X1 _5545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1957_),
    .B(_1952_),
    .Y(_1958_)
);

OAI21X1 _5546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(_1918_),
    .C(_1958_),
    .Y(_1959_)
);

INVX1 _5547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1918_),
    .Y(_1960_)
);

OAI21X1 _5548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_1769_),
    .C(_1848_),
    .Y(_1961_)
);

NAND2X1 _5549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_854_),
    .Y(_1962_)
);

AND2X2 _5550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_1204_),
    .Y(_1963_)
);

OAI21X1 _5551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1963_),
    .C(_1962_),
    .Y(_1964_)
);

NAND2X1 _5552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_1350_),
    .Y(_1966_)
);

NAND2X1 _5553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(_1966_),
    .Y(_1967_)
);

INVX1 _5554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1778_),
    .Y(_1968_)
);

OAI21X1 _5555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1967_),
    .B(_1774_),
    .C(_1968_),
    .Y(_1969_)
);

AOI21X1 _5556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1788_),
    .B(_1964_),
    .C(_1969_),
    .Y(_1970_)
);

NAND3X1 _5557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_295_),
    .B(_125_),
    .C(_486_),
    .Y(_1971_)
);

NOR2X1 _5558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2765_),
    .B(_1971_),
    .Y(_1972_)
);

NOR2X1 _5559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1782_),
    .Y(_1973_)
);

OAI21X1 _5560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1972_),
    .B(_492_),
    .C(_1973_),
    .Y(_1974_)
);

AOI21X1 _5561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .B(_1974_),
    .C(_1913_),
    .Y(_1975_)
);

OAI21X1 _5562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .B(_1961_),
    .C(_1915_),
    .Y(_1977_)
);

AND2X2 _5563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1952_),
    .B(_1957_),
    .Y(_1978_)
);

NAND3X1 _5564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1960_),
    .B(_1978_),
    .C(_1977_),
    .Y(_1979_)
);

NAND2X1 _5565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1959_),
    .B(_1979_),
    .Y(_1_[27])
);

OAI21X1 _5566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .B(_1908_),
    .C(_1978_),
    .Y(_1980_)
);

NOR3X1 _5567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1793_),
    .B(_1852_),
    .C(_1980_),
    .Y(_1981_)
);

OAI21X1 _5568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1790_),
    .B(_1783_),
    .C(_1981_),
    .Y(_1982_)
);

NAND3X1 _5569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1906_),
    .B(_1907_),
    .C(_1847_),
    .Y(_1983_)
);

NAND2X1 _5570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1850_),
    .B(_1917_),
    .Y(_1984_)
);

AOI21X1 _5571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1983_),
    .B(_1984_),
    .C(_1958_),
    .Y(_1985_)
);

NOR2X1 _5572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .B(_1951_),
    .Y(_1987_)
);

OAI21X1 _5573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1918_),
    .B(_1953_),
    .C(_1987_),
    .Y(_1988_)
);

INVX1 _5574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .Y(_1989_)
);

AOI21X1 _5575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .B(_1961_),
    .C(_1989_),
    .Y(_1990_)
);

AOI21X1 _5576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1942_),
    .B(_1941_),
    .C(_1940_),
    .Y(_1991_)
);

OAI21X1 _5577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(_1934_),
    .C(_1936_),
    .Y(_1992_)
);

INVX1 _5578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1927_),
    .Y(_1993_)
);

NAND2X1 _5579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1926_),
    .B(_1933_),
    .Y(_1994_)
);

OAI21X1 _5580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1993_),
    .B(_1931_),
    .C(_1994_),
    .Y(_1995_)
);

OAI22X1 _5581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(_1928_),
    .C(_1930_),
    .D(_1866_),
    .Y(_1996_)
);

NAND2X1 _5582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf2),
    .B(breg_15_bF$buf3),
    .Y(_1998_)
);

NOR2X1 _5583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_1059_),
    .Y(_1999_)
);

INVX1 _5584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1999_),
    .Y(_2000_)
);

NOR2X1 _5585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1928_),
    .B(_2000_),
    .Y(_2001_)
);

AOI21X1 _5586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf3),
    .B(areg_15_bF$buf0),
    .C(_1999_),
    .Y(_2002_)
);

NOR2X1 _5587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2002_),
    .B(_2001_),
    .Y(_2003_)
);

XNOR2X1 _5588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_1998_),
    .Y(_2004_)
);

XOR2X1 _5589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(_1996_),
    .Y(_2005_)
);

NAND2X1 _5590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2005_),
    .B(_1995_),
    .Y(_2006_)
);

INVX1 _5591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2006_),
    .Y(_2007_)
);

NOR2X1 _5592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2005_),
    .B(_1995_),
    .Y(_2009_)
);

NOR2X1 _5593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2009_),
    .B(_2007_),
    .Y(_2010_)
);

XOR2X1 _5594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1992_),
    .B(_2010_),
    .Y(_2011_)
);

OR2X2 _5595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2011_),
    .B(_1991_),
    .Y(_2012_)
);

NAND2X1 _5596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1991_),
    .B(_2011_),
    .Y(_2013_)
);

AND2X2 _5597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2012_),
    .B(_2013_),
    .Y(_2014_)
);

OAI21X1 _5598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1950_),
    .B(_1901_),
    .C(_1948_),
    .Y(_2015_)
);

XOR2X1 _5599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .B(_2015_),
    .Y(_2016_)
);

INVX1 _5600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .Y(_2017_)
);

AOI21X1 _5601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(_1982_),
    .C(_2017_),
    .Y(_2018_)
);

NAND3X1 _5602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1912_),
    .B(_1773_),
    .C(_1985_),
    .Y(_2020_)
);

OAI21X1 _5603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1791_),
    .B(_2020_),
    .C(_1990_),
    .Y(_2021_)
);

NOR2X1 _5604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(_2021_),
    .Y(_2022_)
);

NOR2X1 _5605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2018_),
    .B(_2022_),
    .Y(_1_[28])
);

INVX1 _5606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .Y(_2023_)
);

NOR2X1 _5607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1956_),
    .B(_2023_),
    .Y(_2024_)
);

INVX1 _5608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .Y(_2025_)
);

AOI21X1 _5609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .B(_1974_),
    .C(_2020_),
    .Y(_2026_)
);

OAI21X1 _5610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1854_),
    .B(_1980_),
    .C(_1988_),
    .Y(_2027_)
);

OAI21X1 _5611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .B(_2027_),
    .C(_2016_),
    .Y(_2028_)
);

NOR2X1 _5612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_2023_),
    .Y(_2030_)
);

NAND2X1 _5613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2010_),
    .B(_1992_),
    .Y(_2031_)
);

NAND2X1 _5614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_2004_),
    .Y(_2032_)
);

INVX1 _5615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2001_),
    .Y(_2033_)
);

OAI21X1 _5616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2002_),
    .B(_1998_),
    .C(_2033_),
    .Y(_2034_)
);

AOI22X1 _5617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_15_bF$buf3),
    .C(areg_14_bF$buf3),
    .D(breg_15_bF$buf2),
    .Y(_2035_)
);

AOI21X1 _5618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1871_),
    .B(_1999_),
    .C(_2035_),
    .Y(_2036_)
);

NAND2X1 _5619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2036_),
    .B(_2034_),
    .Y(_2037_)
);

INVX1 _5620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .Y(_2038_)
);

NOR2X1 _5621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2036_),
    .B(_2034_),
    .Y(_2039_)
);

NOR2X1 _5622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2039_),
    .B(_2038_),
    .Y(_2041_)
);

XNOR2X1 _5623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2041_),
    .B(_2032_),
    .Y(_2042_)
);

XOR2X1 _5624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2042_),
    .B(_2006_),
    .Y(_2043_)
);

NAND2X1 _5625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2043_),
    .B(_2031_),
    .Y(_2044_)
);

OR2X2 _5626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2031_),
    .B(_2043_),
    .Y(_2045_)
);

NAND2X1 _5627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2044_),
    .B(_2045_),
    .Y(_2046_)
);

XOR2X1 _5628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_2013_),
    .Y(_2047_)
);

XOR2X1 _5629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2030_),
    .B(_2047_),
    .Y(_2048_)
);

NAND3X1 _5630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2025_),
    .B(_2048_),
    .C(_2028_),
    .Y(_2049_)
);

INVX1 _5631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2048_),
    .Y(_2050_)
);

OAI21X1 _5632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2018_),
    .B(_2024_),
    .C(_2050_),
    .Y(_2052_)
);

NAND2X1 _5633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2052_),
    .B(_2049_),
    .Y(_1_[29])
);

NAND2X1 _5634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(_2048_),
    .Y(_2053_)
);

INVX1 _5635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .Y(_2054_)
);

OAI21X1 _5636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .B(_2027_),
    .C(_2054_),
    .Y(_2055_)
);

OAI21X1 _5637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2030_),
    .B(_2024_),
    .C(_2047_),
    .Y(_2056_)
);

NOR2X1 _5638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2013_),
    .B(_2046_),
    .Y(_2057_)
);

INVX1 _5639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2041_),
    .Y(_2058_)
);

NOR2X1 _5640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2032_),
    .B(_2058_),
    .Y(_2059_)
);

NOR2X1 _5641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .B(_1999_),
    .Y(_2060_)
);

XNOR2X1 _5642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .B(_2060_),
    .Y(_2062_)
);

XNOR2X1 _5643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2059_),
    .B(_2062_),
    .Y(_2063_)
);

NAND2X1 _5644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2042_),
    .B(_2007_),
    .Y(_2064_)
);

OAI21X1 _5645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2031_),
    .B(_2043_),
    .C(_2064_),
    .Y(_2065_)
);

XNOR2X1 _5646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2063_),
    .Y(_2066_)
);

XOR2X1 _5647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2057_),
    .B(_2066_),
    .Y(_2067_)
);

NAND3X1 _5648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2056_),
    .B(_2067_),
    .C(_2055_),
    .Y(_2068_)
);

AOI21X1 _5649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(_1982_),
    .C(_2053_),
    .Y(_2069_)
);

INVX1 _5650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2056_),
    .Y(_2070_)
);

INVX1 _5651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2067_),
    .Y(_2071_)
);

OAI21X1 _5652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2069_),
    .B(_2070_),
    .C(_2071_),
    .Y(_2073_)
);

NAND2X1 _5653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2068_),
    .Y(_1_[30])
);

NAND2X1 _5654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2066_),
    .B(_2057_),
    .Y(_2074_)
);

OAI21X1 _5655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2069_),
    .B(_2070_),
    .C(_2067_),
    .Y(_2075_)
);

AOI21X1 _5656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2045_),
    .C(_2063_),
    .Y(_2076_)
);

NAND2X1 _5657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2062_),
    .B(_2059_),
    .Y(_2077_)
);

OAI21X1 _5658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .B(_1999_),
    .C(_1871_),
    .Y(_2078_)
);

NAND2X1 _5659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2078_),
    .B(_2077_),
    .Y(_2079_)
);

NOR2X1 _5660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2079_),
    .B(_2076_),
    .Y(_2080_)
);

NAND3X1 _5661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .B(_2080_),
    .C(_2075_),
    .Y(_1_[31])
);

XOR2X1 _5662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_2620_),
    .Y(_1_[1])
);

BUFX2 _5663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[0]),
    .Y(y[0])
);

BUFX2 _5664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[1]),
    .Y(y[1])
);

BUFX2 _5665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[2]),
    .Y(y[2])
);

BUFX2 _5666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[3]),
    .Y(y[3])
);

BUFX2 _5667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[4]),
    .Y(y[4])
);

BUFX2 _5668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[5]),
    .Y(y[5])
);

BUFX2 _5669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[6]),
    .Y(y[6])
);

BUFX2 _5670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[7]),
    .Y(y[7])
);

BUFX2 _5671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[8]),
    .Y(y[8])
);

BUFX2 _5672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[9]),
    .Y(y[9])
);

BUFX2 _5673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[10]),
    .Y(y[10])
);

BUFX2 _5674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[11]),
    .Y(y[11])
);

BUFX2 _5675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[12]),
    .Y(y[12])
);

BUFX2 _5676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[13]),
    .Y(y[13])
);

BUFX2 _5677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[14]),
    .Y(y[14])
);

BUFX2 _5678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[15]),
    .Y(y[15])
);

BUFX2 _5679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[16]),
    .Y(y[16])
);

BUFX2 _5680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[17]),
    .Y(y[17])
);

BUFX2 _5681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[18]),
    .Y(y[18])
);

BUFX2 _5682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[19]),
    .Y(y[19])
);

BUFX2 _5683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[20]),
    .Y(y[20])
);

BUFX2 _5684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[21]),
    .Y(y[21])
);

BUFX2 _5685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[22]),
    .Y(y[22])
);

BUFX2 _5686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[23]),
    .Y(y[23])
);

BUFX2 _5687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[24]),
    .Y(y[24])
);

BUFX2 _5688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[25]),
    .Y(y[25])
);

BUFX2 _5689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[26]),
    .Y(y[26])
);

BUFX2 _5690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[27]),
    .Y(y[27])
);

BUFX2 _5691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[28]),
    .Y(y[28])
);

BUFX2 _5692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[29]),
    .Y(y[29])
);

BUFX2 _5693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[30]),
    .Y(y[30])
);

BUFX2 _5694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_[31]),
    .Y(y[31])
);

DFFPOSX1 _5695_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_0_[0]),
    .Q(_2816_[0])
);

DFFPOSX1 _5696_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1_[1]),
    .Q(_2816_[1])
);

DFFPOSX1 _5697_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1_[2]),
    .Q(_2816_[2])
);

DFFPOSX1 _5698_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1_[3]),
    .Q(_2816_[3])
);

DFFPOSX1 _5699_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1_[4]),
    .Q(_2816_[4])
);

DFFPOSX1 _5700_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1_[5]),
    .Q(_2816_[5])
);

DFFPOSX1 _5701_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1_[6]),
    .Q(_2816_[6])
);

DFFPOSX1 _5702_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1_[7]),
    .Q(_2816_[7])
);

DFFPOSX1 _5703_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1_[8]),
    .Q(_2816_[8])
);

DFFPOSX1 _5704_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1_[9]),
    .Q(_2816_[9])
);

DFFPOSX1 _5705_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1_[10]),
    .Q(_2816_[10])
);

DFFPOSX1 _5706_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1_[11]),
    .Q(_2816_[11])
);

DFFPOSX1 _5707_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1_[12]),
    .Q(_2816_[12])
);

DFFPOSX1 _5708_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1_[13]),
    .Q(_2816_[13])
);

DFFPOSX1 _5709_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1_[14]),
    .Q(_2816_[14])
);

DFFPOSX1 _5710_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1_[15]),
    .Q(_2816_[15])
);

DFFPOSX1 _5711_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1_[16]),
    .Q(_2816_[16])
);

DFFPOSX1 _5712_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1_[17]),
    .Q(_2816_[17])
);

DFFPOSX1 _5713_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1_[18]),
    .Q(_2816_[18])
);

DFFPOSX1 _5714_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1_[19]),
    .Q(_2816_[19])
);

DFFPOSX1 _5715_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1_[20]),
    .Q(_2816_[20])
);

DFFPOSX1 _5716_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1_[21]),
    .Q(_2816_[21])
);

DFFPOSX1 _5717_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1_[22]),
    .Q(_2816_[22])
);

DFFPOSX1 _5718_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1_[23]),
    .Q(_2816_[23])
);

DFFPOSX1 _5719_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(_1_[24]),
    .Q(_2816_[24])
);

DFFPOSX1 _5720_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(_1_[25]),
    .Q(_2816_[25])
);

DFFPOSX1 _5721_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(_1_[26]),
    .Q(_2816_[26])
);

DFFPOSX1 _5722_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(_1_[27]),
    .Q(_2816_[27])
);

DFFPOSX1 _5723_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(_1_[28]),
    .Q(_2816_[28])
);

DFFPOSX1 _5724_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(_1_[29]),
    .Q(_2816_[29])
);

DFFPOSX1 _5725_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(_1_[30]),
    .Q(_2816_[30])
);

DFFPOSX1 _5726_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(_1_[31]),
    .Q(_2816_[31])
);

DFFPOSX1 _5727_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(a[0]),
    .Q(areg[0])
);

DFFPOSX1 _5728_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(a[1]),
    .Q(areg[1])
);

DFFPOSX1 _5729_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(a[2]),
    .Q(areg[2])
);

DFFPOSX1 _5730_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(a[3]),
    .Q(areg[3])
);

DFFPOSX1 _5731_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(a[4]),
    .Q(areg[4])
);

DFFPOSX1 _5732_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(a[5]),
    .Q(areg[5])
);

DFFPOSX1 _5733_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(a[6]),
    .Q(areg[6])
);

DFFPOSX1 _5734_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(a[7]),
    .Q(areg[7])
);

DFFPOSX1 _5735_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(a[8]),
    .Q(areg[8])
);

DFFPOSX1 _5736_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(a[9]),
    .Q(areg[9])
);

DFFPOSX1 _5737_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(a[10]),
    .Q(areg[10])
);

DFFPOSX1 _5738_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(a[11]),
    .Q(areg[11])
);

DFFPOSX1 _5739_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(a[12]),
    .Q(areg[12])
);

DFFPOSX1 _5740_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(a[13]),
    .Q(areg[13])
);

DFFPOSX1 _5741_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(a[14]),
    .Q(areg[14])
);

DFFPOSX1 _5742_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(a[15]),
    .Q(areg[15])
);

DFFPOSX1 _5743_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(b[0]),
    .Q(breg[0])
);

DFFPOSX1 _5744_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(b[1]),
    .Q(breg[1])
);

DFFPOSX1 _5745_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(b[2]),
    .Q(breg[2])
);

DFFPOSX1 _5746_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(b[3]),
    .Q(breg[3])
);

DFFPOSX1 _5747_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(b[4]),
    .Q(breg[4])
);

DFFPOSX1 _5748_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(b[5]),
    .Q(breg[5])
);

DFFPOSX1 _5749_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(b[6]),
    .Q(breg[6])
);

DFFPOSX1 _5750_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(b[7]),
    .Q(breg[7])
);

DFFPOSX1 _5751_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(b[8]),
    .Q(breg[8])
);

DFFPOSX1 _5752_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(b[9]),
    .Q(breg[9])
);

DFFPOSX1 _5753_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(b[10]),
    .Q(breg[10])
);

DFFPOSX1 _5754_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(b[11]),
    .Q(breg[11])
);

DFFPOSX1 _5755_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(b[12]),
    .Q(breg[12])
);

DFFPOSX1 _5756_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(b[13]),
    .Q(breg[13])
);

DFFPOSX1 _5757_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(b[14]),
    .Q(breg[14])
);

DFFPOSX1 _5758_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(b[15]),
    .Q(breg[15])
);

endmodule
