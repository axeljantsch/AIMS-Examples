/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module multiplierBeh(
    inout vdd,
    inout gnd,
    input [31:0] a,
    input [31:0] b,
    input clk,
    output [63:0] y
);

wire _11689_ ;
wire _11269_ ;
wire _9837_ ;
wire _9417_ ;
wire _4972_ ;
wire _4552_ ;
wire _4132_ ;
wire _5757_ ;
wire _5337_ ;
wire _9590_ ;
wire _9170_ ;
wire [31:0] a ;
wire [31:0] b ;
wire _1677_ ;
wire _1257_ ;
wire _7903_ ;
wire [63:0] y ;
wire _5090_ ;
wire _588_ ;
wire _168_ ;
wire _11901_ ;
wire _3823_ ;
wire _3403_ ;
wire _6295_ ;
wire _10293_ ;
wire _4608_ ;
wire _8861_ ;
wire _8441_ ;
wire _8021_ ;
wire _11498_ ;
wire _11078_ ;
wire _9646_ ;
wire _9226_ ;
wire _4781_ ;
wire _4361_ ;
wire _800_ ;
wire _5986_ ;
wire _5566_ ;
wire _5146_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _7712_ ;
wire _10769_ ;
wire _10349_ ;
wire _397_ ;
wire _11710_ ;
wire _8917_ ;
wire _3632_ ;
wire _3212_ ;
wire _4837_ ;
wire _4417_ ;
wire _8670_ ;
wire _8250_ ;
wire _9875_ ;
wire _9455_ ;
wire _9035_ ;
wire _4590_ ;
wire _4170_ ;
wire _2903_ ;
wire _5795_ ;
wire _5375_ ;
wire _1295_ ;
wire _7941_ ;
wire _7521_ ;
wire _7101_ ;
wire _10998_ ;
wire _10578_ ;
wire _10158_ ;
wire _8726_ ;
wire _8306_ ;
wire _3861_ ;
wire _3441_ ;
wire _3021_ ;
wire _4646_ ;
wire _4226_ ;
wire _9684_ ;
wire _9264_ ;
wire _2712_ ;
wire _5184_ ;
wire _3917_ ;
wire _6389_ ;
wire _7750_ ;
wire _7330_ ;
wire _10387_ ;
wire _8955_ ;
wire _8535_ ;
wire _8115_ ;
wire _3670_ ;
wire _3250_ ;
wire _4875_ ;
wire _4455_ ;
wire _4035_ ;
wire _6601_ ;
wire _9493_ ;
wire _9073_ ;
wire _7806_ ;
wire _2941_ ;
wire _2521_ ;
wire _2101_ ;
wire _11804_ ;
wire _3726_ ;
wire _3306_ ;
wire _6198_ ;
wire _10196_ ;
wire _8764_ ;
wire _8344_ ;
wire _9969_ ;
wire _9549_ ;
wire _9129_ ;
wire _4684_ ;
wire _4264_ ;
wire _703_ ;
wire _5889_ ;
wire _5469_ ;
wire _5049_ ;
wire _6830_ ;
wire _6410_ ;
wire _1389_ ;
wire _7615_ ;
wire _2750_ ;
wire _2330_ ;
wire _11613_ ;
wire _3955_ ;
wire _3535_ ;
wire _3115_ ;
wire _8993_ ;
wire _8573_ ;
wire _8153_ ;
wire _19_ ;
wire _1601_ ;
wire _9778_ ;
wire _9358_ ;
wire _4493_ ;
wire _4073_ ;
wire _932_ ;
wire _512_ ;
wire _2806_ ;
wire _5698_ ;
wire _5278_ ;
wire _1198_ ;
wire _7844_ ;
wire _7424_ ;
wire _7004_ ;
wire _11842_ ;
wire _11422_ ;
wire _11002_ ;
wire _8629_ ;
wire _8209_ ;
wire _3764_ ;
wire _3344_ ;
wire _4969_ ;
wire _4549_ ;
wire _4129_ ;
wire _5910_ ;
wire _8382_ ;
wire _1830_ ;
wire _1410_ ;
wire _9587_ ;
wire _9167_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _5087_ ;
wire _7653_ ;
wire _7233_ ;
wire _11651_ ;
wire _11231_ ;
wire _8858_ ;
wire _8438_ ;
wire _8018_ ;
wire _3993_ ;
wire _3573_ ;
wire _3153_ ;
wire _4778_ ;
wire _4358_ ;
wire _8191_ ;
wire _57_ ;
wire _6924_ ;
wire _6504_ ;
wire _9396_ ;
wire _10922_ ;
wire _10502_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _7709_ ;
wire _2844_ ;
wire _2424_ ;
wire _2004_ ;
wire _11707_ ;
wire _3629_ ;
wire _3209_ ;
wire _7882_ ;
wire _7462_ ;
wire _7042_ ;
wire _10099_ ;
wire _11880_ ;
wire _11460_ ;
wire _11040_ ;
wire _8667_ ;
wire _8247_ ;
wire _3382_ ;
wire _4587_ ;
wire _4167_ ;
wire _606_ ;
wire _6733_ ;
wire _6313_ ;
wire _10731_ ;
wire _10311_ ;
wire _7938_ ;
wire _7518_ ;
wire _2653_ ;
wire _2233_ ;
wire _11516_ ;
wire _3858_ ;
wire _3438_ ;
wire _3018_ ;
wire _7691_ ;
wire _7271_ ;
wire _8896_ ;
wire _8476_ ;
wire _8056_ ;
wire _3191_ ;
wire _1924_ ;
wire _1504_ ;
wire _4396_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _6962_ ;
wire _6542_ ;
wire _6122_ ;
wire _10960_ ;
wire _10540_ ;
wire _10120_ ;
wire _7747_ ;
wire _7327_ ;
wire _2882_ ;
wire _2462_ ;
wire _2042_ ;
wire _11745_ ;
wire _11325_ ;
wire _3667_ ;
wire _3247_ ;
wire _7080_ ;
wire _5813_ ;
wire _8285_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2938_ ;
wire _2518_ ;
wire _6771_ ;
wire _6351_ ;
wire _7976_ ;
wire _7556_ ;
wire _7136_ ;
wire _2691_ ;
wire _2271_ ;
wire _11554_ ;
wire _11134_ ;
wire _3896_ ;
wire _3476_ ;
wire _3056_ ;
wire _9702_ ;
wire _5622_ ;
wire _5202_ ;
wire _8094_ ;
wire _6827_ ;
wire _6407_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _9299_ ;
wire _10825_ ;
wire _10405_ ;
wire _873_ ;
wire _453_ ;
wire _2747_ ;
wire _2327_ ;
wire _6580_ ;
wire _6160_ ;
wire _7785_ ;
wire _7365_ ;
wire _2080_ ;
wire _11783_ ;
wire _11363_ ;
wire _3285_ ;
wire _9931_ ;
wire _9511_ ;
wire _5851_ ;
wire _5431_ ;
wire _5011_ ;
wire _929_ ;
wire _509_ ;
wire _6636_ ;
wire _6216_ ;
wire _1771_ ;
wire _1351_ ;
wire _10634_ ;
wire _10214_ ;
wire _682_ ;
wire _262_ ;
wire _2976_ ;
wire _2556_ ;
wire _2136_ ;
wire _11839_ ;
wire _11419_ ;
wire _4702_ ;
wire _7594_ ;
wire _7174_ ;
wire _11592_ ;
wire _11172_ ;
wire _5907_ ;
wire _8799_ ;
wire _8379_ ;
wire _3094_ ;
wire _9740_ ;
wire _9320_ ;
wire _1827_ ;
wire _1407_ ;
wire _4299_ ;
wire _5660_ ;
wire _5240_ ;
wire _738_ ;
wire _318_ ;
wire _6865_ ;
wire _6445_ ;
wire _6025_ ;
wire _1580_ ;
wire _1160_ ;
wire _10863_ ;
wire _10443_ ;
wire _10023_ ;
wire _491_ ;
wire _2785_ ;
wire _2365_ ;
wire _11648_ ;
wire _11228_ ;
wire _4931_ ;
wire _4511_ ;
wire _5716_ ;
wire _8188_ ;
wire _1636_ ;
wire _1216_ ;
wire _10919_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _6674_ ;
wire _6254_ ;
wire _10672_ ;
wire _10252_ ;
wire _7879_ ;
wire _7459_ ;
wire _7039_ ;
wire _2594_ ;
wire _2174_ ;
wire _8820_ ;
wire _8400_ ;
wire _11877_ ;
wire _11457_ ;
wire _11037_ ;
wire _3799_ ;
wire _3379_ ;
wire _9605_ ;
wire _4740_ ;
wire _4320_ ;
wire _5945_ ;
wire _5525_ ;
wire _5105_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _10728_ ;
wire _10308_ ;
wire _776_ ;
wire _356_ ;
wire _6483_ ;
wire _6063_ ;
wire _10481_ ;
wire _10061_ ;
wire _7688_ ;
wire _7268_ ;
wire _11686_ ;
wire _11266_ ;
wire _3188_ ;
wire _9834_ ;
wire _9414_ ;
wire _5754_ ;
wire _5334_ ;
wire _6959_ ;
wire _6539_ ;
wire _6119_ ;
wire _1674_ ;
wire _1254_ ;
wire _7900_ ;
wire _10957_ ;
wire _10537_ ;
wire _10117_ ;
wire _585_ ;
wire _165_ ;
wire _2879_ ;
wire _2459_ ;
wire _2039_ ;
wire _3820_ ;
wire _3400_ ;
wire _6292_ ;
wire _10290_ ;
wire _4605_ ;
wire _7497_ ;
wire _7077_ ;
wire _11495_ ;
wire _11075_ ;
wire _9643_ ;
wire _9223_ ;
wire _5983_ ;
wire _5563_ ;
wire _5143_ ;
wire areg_25_bF$buf0 ;
wire areg_25_bF$buf1 ;
wire areg_25_bF$buf2 ;
wire areg_25_bF$buf3 ;
wire areg_25_bF$buf4 ;
wire _6768_ ;
wire _6348_ ;
wire _1483_ ;
wire _1063_ ;
wire _10766_ ;
wire _10346_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _8914_ ;
wire _4834_ ;
wire _4414_ ;
wire _5619_ ;
wire _9872_ ;
wire _9452_ ;
wire _9032_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _2900_ ;
wire _5792_ ;
wire _5372_ ;
wire _6997_ ;
wire _6577_ ;
wire _6157_ ;
wire _1292_ ;
wire _10995_ ;
wire _10575_ ;
wire _10155_ ;
wire _2497_ ;
wire _2077_ ;
wire _8723_ ;
wire _8303_ ;
wire _9928_ ;
wire _9508_ ;
wire _4643_ ;
wire _4223_ ;
wire _5848_ ;
wire _5428_ ;
wire _5008_ ;
wire _9681_ ;
wire _9261_ ;
wire _1768_ ;
wire _1348_ ;
wire _5181_ ;
wire _679_ ;
wire _259_ ;
wire _3914_ ;
wire _6386_ ;
wire _10384_ ;
wire _8952_ ;
wire _8532_ ;
wire _8112_ ;
wire _11589_ ;
wire _11169_ ;
wire _9737_ ;
wire _9317_ ;
wire _4872_ ;
wire _4452_ ;
wire _4032_ ;
wire _5657_ ;
wire _5237_ ;
wire _9490_ ;
wire _9070_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _7803_ ;
wire _488_ ;
wire _11801_ ;
wire _3723_ ;
wire _3303_ ;
wire _6195_ ;
wire _10193_ ;
wire _4928_ ;
wire _4508_ ;
wire _8761_ ;
wire _8341_ ;
wire _11398_ ;
wire _9966_ ;
wire _9546_ ;
wire _9126_ ;
wire _4681_ ;
wire _4261_ ;
wire _700_ ;
wire _5886_ ;
wire _5466_ ;
wire _5046_ ;
wire _1386_ ;
wire _7612_ ;
wire _10669_ ;
wire _10249_ ;
wire _297_ ;
wire _11610_ ;
wire _8817_ ;
wire _3952_ ;
wire _3532_ ;
wire _3112_ ;
wire areg_7_bF$buf0 ;
wire areg_7_bF$buf1 ;
wire areg_7_bF$buf2 ;
wire areg_7_bF$buf3 ;
wire areg_7_bF$buf4 ;
wire _4737_ ;
wire _4317_ ;
wire _8990_ ;
wire _8570_ ;
wire _8150_ ;
wire _16_ ;
wire _9775_ ;
wire _9355_ ;
wire _4490_ ;
wire _4070_ ;
wire _2803_ ;
wire _5695_ ;
wire _5275_ ;
wire _1195_ ;
wire _7841_ ;
wire _7421_ ;
wire _7001_ ;
wire _10898_ ;
wire _10478_ ;
wire _10058_ ;
wire _8626_ ;
wire _8206_ ;
wire _3761_ ;
wire _3341_ ;
wire _4966_ ;
wire _4546_ ;
wire _4126_ ;
wire _9584_ ;
wire _9164_ ;
wire _2612_ ;
wire _5084_ ;
wire _3817_ ;
wire _6289_ ;
wire _7650_ ;
wire _7230_ ;
wire _10287_ ;
wire _8855_ ;
wire _8435_ ;
wire _8015_ ;
wire _3990_ ;
wire _3570_ ;
wire _3150_ ;
wire _4775_ ;
wire _4355_ ;
wire _54_ ;
wire _6921_ ;
wire _6501_ ;
wire _9393_ ;
wire _7706_ ;
wire _2841_ ;
wire _2421_ ;
wire _2001_ ;
wire _11704_ ;
wire _3626_ ;
wire _3206_ ;
wire _6098_ ;
wire _10096_ ;
wire _8664_ ;
wire _8244_ ;
wire _9869_ ;
wire _9449_ ;
wire _9029_ ;
wire _4584_ ;
wire _4164_ ;
wire _603_ ;
wire _5789_ ;
wire _5369_ ;
wire _6730_ ;
wire _6310_ ;
wire _1289_ ;
wire _7935_ ;
wire _7515_ ;
wire _2650_ ;
wire _2230_ ;
wire _11513_ ;
wire _3855_ ;
wire _3435_ ;
wire _3015_ ;
wire _8893_ ;
wire _8473_ ;
wire _8053_ ;
wire _1921_ ;
wire _1501_ ;
wire _9678_ ;
wire _9258_ ;
wire _4393_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _5598_ ;
wire _5178_ ;
wire _92_ ;
wire _1098_ ;
wire _7744_ ;
wire _7324_ ;
wire _11742_ ;
wire _11322_ ;
wire _8949_ ;
wire _8529_ ;
wire _8109_ ;
wire _3664_ ;
wire _3244_ ;
wire _4869_ ;
wire _4449_ ;
wire _4029_ ;
wire _5810_ ;
wire _8282_ ;
wire _1730_ ;
wire _1310_ ;
wire _9487_ ;
wire _9067_ ;
wire _641_ ;
wire _221_ ;
wire _2935_ ;
wire _2515_ ;
wire _7973_ ;
wire _7553_ ;
wire _7133_ ;
wire _11551_ ;
wire _11131_ ;
wire _8758_ ;
wire _8338_ ;
wire _3893_ ;
wire _3473_ ;
wire _3053_ ;
wire _4678_ ;
wire _4258_ ;
wire _8091_ ;
wire _6824_ ;
wire _6404_ ;
wire _9296_ ;
wire _10822_ ;
wire _10402_ ;
wire _870_ ;
wire _450_ ;
wire _7609_ ;
wire _2744_ ;
wire _2324_ ;
wire _11607_ ;
wire _3949_ ;
wire _3529_ ;
wire _3109_ ;
wire _7782_ ;
wire _7362_ ;
wire _11780_ ;
wire _11360_ ;
wire _8987_ ;
wire _8567_ ;
wire _8147_ ;
wire _3282_ ;
wire _4487_ ;
wire _4067_ ;
wire _926_ ;
wire _506_ ;
wire _6633_ ;
wire _6213_ ;
wire _10631_ ;
wire _10211_ ;
wire _7838_ ;
wire _7418_ ;
wire _2973_ ;
wire _2553_ ;
wire _2133_ ;
wire _11836_ ;
wire _11416_ ;
wire _3758_ ;
wire _3338_ ;
wire _7591_ ;
wire _7171_ ;
wire _5904_ ;
wire _8796_ ;
wire _8376_ ;
wire _3091_ ;
wire _1824_ ;
wire _1404_ ;
wire _4296_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _6862_ ;
wire _6442_ ;
wire _6022_ ;
wire _10860_ ;
wire _10440_ ;
wire _10020_ ;
wire _7647_ ;
wire _7227_ ;
wire _2782_ ;
wire _2362_ ;
wire _11645_ ;
wire _11225_ ;
wire _3987_ ;
wire _3567_ ;
wire _3147_ ;
wire _5713_ ;
wire _8185_ ;
wire _6918_ ;
wire _1633_ ;
wire _1213_ ;
wire _10916_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2838_ ;
wire _2418_ ;
wire _6671_ ;
wire _6251_ ;
wire _7876_ ;
wire _7456_ ;
wire _7036_ ;
wire _2591_ ;
wire _2171_ ;
wire _11874_ ;
wire _11454_ ;
wire _11034_ ;
wire _3796_ ;
wire _3376_ ;
wire _9602_ ;
wire _5942_ ;
wire _5522_ ;
wire _5102_ ;
wire _6727_ ;
wire _6307_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _9199_ ;
wire _10725_ ;
wire _10305_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _6480_ ;
wire _6060_ ;
wire _7685_ ;
wire _7265_ ;
wire _11683_ ;
wire _11263_ ;
wire _3185_ ;
wire _9831_ ;
wire _9411_ ;
wire _1918_ ;
wire _5751_ ;
wire _5331_ ;
wire _829_ ;
wire _409_ ;
wire breg_27_bF$buf0 ;
wire breg_27_bF$buf1 ;
wire _89_ ;
wire breg_27_bF$buf2 ;
wire breg_27_bF$buf3 ;
wire _6956_ ;
wire breg_27_bF$buf4 ;
wire _6536_ ;
wire breg_27_bF$buf5 ;
wire _6116_ ;
wire _1671_ ;
wire _1251_ ;
wire _10954_ ;
wire _10534_ ;
wire _10114_ ;
wire _582_ ;
wire _162_ ;
wire _2876_ ;
wire _2456_ ;
wire _2036_ ;
wire _11739_ ;
wire _11319_ ;
wire _4602_ ;
wire _7494_ ;
wire _7074_ ;
wire _11492_ ;
wire _11072_ ;
wire _5807_ ;
wire _8699_ ;
wire _8279_ ;
wire breg_5_bF$buf0 ;
wire breg_5_bF$buf1 ;
wire breg_5_bF$buf2 ;
wire breg_5_bF$buf3 ;
wire _9640_ ;
wire _9220_ ;
wire _1727_ ;
wire _1307_ ;
wire _4199_ ;
wire _5980_ ;
wire _5560_ ;
wire _5140_ ;
wire _638_ ;
wire _218_ ;
wire _6765_ ;
wire _6345_ ;
wire _1480_ ;
wire _1060_ ;
wire _10763_ ;
wire _10343_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _8911_ ;
wire _11548_ ;
wire _11128_ ;
wire _3146__bF$buf0 ;
wire _3146__bF$buf1 ;
wire _3146__bF$buf2 ;
wire _3146__bF$buf3 ;
wire _4831_ ;
wire _4411_ ;
wire _5616_ ;
wire _8088_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _10819_ ;
wire _867_ ;
wire _447_ ;
wire _6994_ ;
wire _6574_ ;
wire _6154_ ;
wire _10992_ ;
wire _10572_ ;
wire _10152_ ;
wire _7779_ ;
wire _7359_ ;
wire _2494_ ;
wire _2074_ ;
wire _8720_ ;
wire _8300_ ;
wire _11777_ ;
wire _11357_ ;
wire _3699_ ;
wire _3279_ ;
wire _9925_ ;
wire _9505_ ;
wire _4640_ ;
wire _4220_ ;
wire _5845_ ;
wire _5425_ ;
wire _5005_ ;
wire _1765_ ;
wire _1345_ ;
wire _10628_ ;
wire _10208_ ;
wire _676_ ;
wire _256_ ;
wire _3911_ ;
wire _6383_ ;
wire _10381_ ;
wire _7588_ ;
wire _7168_ ;
wire _11586_ ;
wire _11166_ ;
wire _3088_ ;
wire _9734_ ;
wire _9314_ ;
wire _5654_ ;
wire _5234_ ;
wire _6859_ ;
wire _6439_ ;
wire _6019_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _7800_ ;
wire _10857_ ;
wire _10437_ ;
wire _10017_ ;
wire _485_ ;
wire _2779_ ;
wire _2359_ ;
wire _3720_ ;
wire _3300_ ;
wire _6192_ ;
wire _10190_ ;
wire _4925_ ;
wire _4505_ ;
wire _7397_ ;
wire _11395_ ;
wire _9963_ ;
wire _9543_ ;
wire _9123_ ;
wire _5883_ ;
wire _5463_ ;
wire _5043_ ;
wire _6668_ ;
wire _6248_ ;
wire _1383_ ;
wire _10666_ ;
wire _10246_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _8814_ ;
wire _4734_ ;
wire _4314_ ;
wire _5939_ ;
wire _5519_ ;
wire _13_ ;
wire _9772_ ;
wire _9352_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _2800_ ;
wire _5692_ ;
wire _5272_ ;
wire _6897_ ;
wire _6477_ ;
wire _6057_ ;
wire _1192_ ;
wire _10895_ ;
wire _10475_ ;
wire _10055_ ;
wire _2397_ ;
wire _8623_ ;
wire _8203_ ;
wire _9828_ ;
wire _9408_ ;
wire _4963_ ;
wire _4543_ ;
wire _4123_ ;
wire _5748_ ;
wire _5328_ ;
wire _9581_ ;
wire _9161_ ;
wire _1668_ ;
wire _1248_ ;
wire _5081_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _3814_ ;
wire _6286_ ;
wire _10284_ ;
wire _8852_ ;
wire _8432_ ;
wire _8012_ ;
wire _11489_ ;
wire _11069_ ;
wire _9637_ ;
wire _9217_ ;
wire _4772_ ;
wire _4352_ ;
wire _5977_ ;
wire _5557_ ;
wire _5137_ ;
wire _51_ ;
wire _9390_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _7703_ ;
wire _388_ ;
wire _11701_ ;
wire _8908_ ;
wire _3623_ ;
wire _3203_ ;
wire _6095_ ;
wire _10093_ ;
wire _4828_ ;
wire _4408_ ;
wire _8661_ ;
wire _8241_ ;
wire _11298_ ;
wire _9866_ ;
wire _9446_ ;
wire _9026_ ;
wire _4581_ ;
wire _4161_ ;
wire _600_ ;
wire _5786_ ;
wire _5366_ ;
wire _1286_ ;
wire _7932_ ;
wire _7512_ ;
wire _10989_ ;
wire _10569_ ;
wire _10149_ ;
wire _197_ ;
wire _11510_ ;
wire _8717_ ;
wire _3852_ ;
wire _3432_ ;
wire _3012_ ;
wire _4637_ ;
wire _4217_ ;
wire _8890_ ;
wire _8470_ ;
wire _8050_ ;
wire _9675_ ;
wire _9255_ ;
wire _4390_ ;
wire _2703_ ;
wire _5595_ ;
wire _5175_ ;
wire _3908_ ;
wire _1095_ ;
wire _7741_ ;
wire _7321_ ;
wire _10798_ ;
wire _10378_ ;
wire _8946_ ;
wire _8526_ ;
wire _8106_ ;
wire _3661_ ;
wire _3241_ ;
wire _4866_ ;
wire _4446_ ;
wire _4026_ ;
wire _9484_ ;
wire _9064_ ;
wire _2932_ ;
wire _2512_ ;
wire _3717_ ;
wire _6189_ ;
wire _7970_ ;
wire _7550_ ;
wire _7130_ ;
wire _10187_ ;
wire _8755_ ;
wire _8335_ ;
wire _3890_ ;
wire _3470_ ;
wire _3050_ ;
wire areg_20_bF$buf0 ;
wire areg_20_bF$buf1 ;
wire areg_20_bF$buf2 ;
wire areg_20_bF$buf3 ;
wire areg_20_bF$buf4 ;
wire _4675_ ;
wire _4255_ ;
wire _6821_ ;
wire _6401_ ;
wire _9293_ ;
wire _7606_ ;
wire _2741_ ;
wire _2321_ ;
wire _11604_ ;
wire _3946_ ;
wire _3526_ ;
wire _3106_ ;
wire _7_ ;
wire _8984_ ;
wire _8564_ ;
wire _8144_ ;
wire _9769_ ;
wire _9349_ ;
wire _4484_ ;
wire _4064_ ;
wire _923_ ;
wire _503_ ;
wire _5689_ ;
wire _5269_ ;
wire _6630_ ;
wire _6210_ ;
wire _1189_ ;
wire _7835_ ;
wire _7415_ ;
wire _2970_ ;
wire _2550_ ;
wire _2130_ ;
wire _11833_ ;
wire _11413_ ;
wire _3755_ ;
wire _3335_ ;
wire _5901_ ;
wire _8793_ ;
wire _8373_ ;
wire _1821_ ;
wire _1401_ ;
wire _9998_ ;
wire _9578_ ;
wire _9158_ ;
wire _4293_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _5498_ ;
wire _5078_ ;
wire _7644_ ;
wire _7224_ ;
wire _11642_ ;
wire _11222_ ;
wire _8849_ ;
wire _8429_ ;
wire _8009_ ;
wire _3984_ ;
wire _3564_ ;
wire _3144_ ;
wire _4769_ ;
wire _4349_ ;
wire _5710_ ;
wire _8182_ ;
wire _48_ ;
wire _6915_ ;
wire _1630_ ;
wire _1210_ ;
wire _9387_ ;
wire _10913_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2835_ ;
wire _2415_ ;
wire _7873_ ;
wire _7453_ ;
wire _7033_ ;
wire _11871_ ;
wire _11451_ ;
wire _11031_ ;
wire _8658_ ;
wire _8238_ ;
wire _3793_ ;
wire _3373_ ;
wire _4998_ ;
wire _4578_ ;
wire _4158_ ;
wire areg_2_bF$buf0 ;
wire areg_2_bF$buf1 ;
wire areg_2_bF$buf2 ;
wire areg_2_bF$buf3 ;
wire _6724_ ;
wire areg_2_bF$buf4 ;
wire _6304_ ;
wire _9196_ ;
wire _10722_ ;
wire _10302_ ;
wire _770_ ;
wire _350_ ;
wire _7929_ ;
wire _7509_ ;
wire _2644_ ;
wire _2224_ ;
wire _11507_ ;
wire _3849_ ;
wire _3429_ ;
wire _3009_ ;
wire _7682_ ;
wire _7262_ ;
wire _11680_ ;
wire _11260_ ;
wire _8887_ ;
wire _8467_ ;
wire _8047_ ;
wire _3182_ ;
wire _1915_ ;
wire _4387_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _6953_ ;
wire _6533_ ;
wire _6113_ ;
wire _10951_ ;
wire _10531_ ;
wire _10111_ ;
wire _7738_ ;
wire _7318_ ;
wire _2873_ ;
wire _2453_ ;
wire _2033_ ;
wire _11736_ ;
wire _11316_ ;
wire _3658_ ;
wire _3238_ ;
wire _7491_ ;
wire _7071_ ;
wire _5804_ ;
wire _8696_ ;
wire _8276_ ;
wire _1724_ ;
wire _1304_ ;
wire _4196_ ;
wire _635_ ;
wire _215_ ;
wire _2929_ ;
wire _2509_ ;
wire _6762_ ;
wire _6342_ ;
wire _10760_ ;
wire _10340_ ;
wire _7967_ ;
wire _7547_ ;
wire _7127_ ;
wire _2682_ ;
wire _2262_ ;
wire _11545_ ;
wire _11125_ ;
wire _3887_ ;
wire _3467_ ;
wire _3047_ ;
wire _5613_ ;
wire _8085_ ;
wire _6818_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _10816_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _6991_ ;
wire _6571_ ;
wire _6151_ ;
wire _7776_ ;
wire _7356_ ;
wire _2491_ ;
wire _2071_ ;
wire _11774_ ;
wire _11354_ ;
wire _3696_ ;
wire _3276_ ;
wire _9922_ ;
wire _9502_ ;
wire _5842_ ;
wire _5422_ ;
wire _5002_ ;
wire _6627_ ;
wire breg_19_bF$buf0 ;
wire _6207_ ;
wire breg_19_bF$buf1 ;
wire breg_19_bF$buf2 ;
wire breg_19_bF$buf3 ;
wire _1762_ ;
wire breg_19_bF$buf4 ;
wire _1342_ ;
wire breg_19_bF$buf5 ;
wire _9099_ ;
wire _10625_ ;
wire _10205_ ;
wire _673_ ;
wire _253_ ;
wire _2967_ ;
wire _2547_ ;
wire _2127_ ;
wire _6380_ ;
wire _7585_ ;
wire _7165_ ;
wire _11583_ ;
wire _11163_ ;
wire _3085_ ;
wire _9731_ ;
wire _9311_ ;
wire _1818_ ;
wire _5651_ ;
wire _5231_ ;
wire _729_ ;
wire _309_ ;
wire _6856_ ;
wire _6436_ ;
wire _6016_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _10854_ ;
wire _10434_ ;
wire _10014_ ;
wire _482_ ;
wire _2776_ ;
wire _2356_ ;
wire _11639_ ;
wire _11219_ ;
wire _4922_ ;
wire _4502_ ;
wire _7394_ ;
wire _11392_ ;
wire _5707_ ;
wire _8599_ ;
wire _8179_ ;
wire _9960_ ;
wire _9540_ ;
wire _9120_ ;
wire _1627_ ;
wire _1207_ ;
wire _4099_ ;
wire _5880_ ;
wire _5460_ ;
wire _5040_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _6665_ ;
wire _6245_ ;
wire _1380_ ;
wire _10663_ ;
wire _10243_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _8811_ ;
wire _11868_ ;
wire _11448_ ;
wire _11028_ ;
wire _4731_ ;
wire _4311_ ;
wire _5936_ ;
wire _5516_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _10719_ ;
wire _767_ ;
wire _347_ ;
wire _6894_ ;
wire _6474_ ;
wire _6054_ ;
wire _10892_ ;
wire _10472_ ;
wire _10052_ ;
wire _7679_ ;
wire _7259_ ;
wire _2394_ ;
wire _8620_ ;
wire _8200_ ;
wire _11677_ ;
wire _11257_ ;
wire _3599_ ;
wire _3179_ ;
wire _9825_ ;
wire _9405_ ;
wire _4960_ ;
wire _4540_ ;
wire _4120_ ;
wire _5745_ ;
wire _5325_ ;
wire _1665_ ;
wire _1245_ ;
wire _10948_ ;
wire _10528_ ;
wire _10108_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _3811_ ;
wire _6283_ ;
wire _10281_ ;
wire _7488_ ;
wire _7068_ ;
wire _11486_ ;
wire _11066_ ;
wire _9634_ ;
wire _9214_ ;
wire _5974_ ;
wire _5554_ ;
wire _5134_ ;
wire _6759_ ;
wire _6339_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _7700_ ;
wire _10757_ ;
wire _10337_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _8905_ ;
wire _3620_ ;
wire _3200_ ;
wire _6092_ ;
wire _4116__bF$buf0 ;
wire _4116__bF$buf1 ;
wire _4116__bF$buf2 ;
wire _4116__bF$buf3 ;
wire _4116__bF$buf4 ;
wire _10090_ ;
wire _4825_ ;
wire _4405_ ;
wire _7297_ ;
wire _11295_ ;
wire _9863_ ;
wire _9443_ ;
wire _9023_ ;
wire _5783_ ;
wire _5363_ ;
wire _6988_ ;
wire _6568_ ;
wire _6148_ ;
wire _1283_ ;
wire _10986_ ;
wire _10566_ ;
wire _10146_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _8714_ ;
wire _9919_ ;
wire _4634_ ;
wire _4214_ ;
wire _5839_ ;
wire _5419_ ;
wire _9672_ ;
wire _9252_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _5592_ ;
wire _5172_ ;
wire _3905_ ;
wire _6797_ ;
wire _6377_ ;
wire _1092_ ;
wire _10795_ ;
wire _10375_ ;
wire _2297_ ;
wire _8943_ ;
wire _8523_ ;
wire _8103_ ;
wire breg_22_bF$buf0 ;
wire breg_22_bF$buf1 ;
wire breg_22_bF$buf2 ;
wire breg_22_bF$buf3 ;
wire breg_22_bF$buf4 ;
wire _9728_ ;
wire _9308_ ;
wire _4863_ ;
wire _4443_ ;
wire _4023_ ;
wire _5648_ ;
wire _5228_ ;
wire _9481_ ;
wire _9061_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire breg_0_bF$buf0 ;
wire breg_0_bF$buf1 ;
wire breg_0_bF$buf2 ;
wire breg_0_bF$buf3 ;
wire _3714_ ;
wire breg_0_bF$buf4 ;
wire breg_0_bF$buf5 ;
wire breg_0_bF$buf6 ;
wire _6186_ ;
wire _10184_ ;
wire _4919_ ;
wire _8752_ ;
wire _8332_ ;
wire _11389_ ;
wire _9957_ ;
wire _9537_ ;
wire _9117_ ;
wire _4672_ ;
wire _4252_ ;
wire _5877_ ;
wire _5457_ ;
wire _5037_ ;
wire _9290_ ;
wire _1797_ ;
wire _1377_ ;
wire _7603_ ;
wire _288_ ;
wire _11601_ ;
wire _8808_ ;
wire _3943_ ;
wire _3523_ ;
wire _3103_ ;
wire _4_ ;
wire _4728_ ;
wire _4308_ ;
wire _8981_ ;
wire _8561_ ;
wire _8141_ ;
wire _11198_ ;
wire _9766_ ;
wire _9346_ ;
wire _4481_ ;
wire _4061_ ;
wire _920_ ;
wire _500_ ;
wire _5686_ ;
wire _5266_ ;
wire _1186_ ;
wire _7832_ ;
wire _7412_ ;
wire _10889_ ;
wire _10469_ ;
wire _10049_ ;
wire _11830_ ;
wire _11410_ ;
wire _8617_ ;
wire _3752_ ;
wire _3332_ ;
wire _4957_ ;
wire _4537_ ;
wire _4117_ ;
wire _8790_ ;
wire _8370_ ;
wire _9995_ ;
wire _9575_ ;
wire _9155_ ;
wire _4290_ ;
wire _2603_ ;
wire _5495_ ;
wire _5075_ ;
wire _3808_ ;
wire _7641_ ;
wire _7221_ ;
wire _10698_ ;
wire _10278_ ;
wire _8846_ ;
wire _8426_ ;
wire _8006_ ;
wire _3981_ ;
wire _3561_ ;
wire _3141_ ;
wire _4766_ ;
wire _4346_ ;
wire areg_31_bF$buf0 ;
wire areg_31_bF$buf1 ;
wire areg_31_bF$buf2 ;
wire areg_31_bF$buf3 ;
wire areg_31_bF$buf4 ;
wire _45_ ;
wire _6912_ ;
wire _9384_ ;
wire _10910_ ;
wire _2832_ ;
wire _2412_ ;
wire _3617_ ;
wire _6089_ ;
wire _7870_ ;
wire _7450_ ;
wire _7030_ ;
wire _10087_ ;
wire _8655_ ;
wire _8235_ ;
wire _3790_ ;
wire _3370_ ;
wire _4995_ ;
wire _4575_ ;
wire _4155_ ;
wire _6721_ ;
wire _6301_ ;
wire _9193_ ;
wire _7926_ ;
wire _7506_ ;
wire _2641_ ;
wire _2221_ ;
wire _11504_ ;
wire _3846_ ;
wire _3426_ ;
wire _3006_ ;
wire _8884_ ;
wire _8464_ ;
wire _8044_ ;
wire _1912_ ;
wire _9669_ ;
wire _9249_ ;
wire _4384_ ;
wire _823_ ;
wire _403_ ;
wire _5589_ ;
wire _5315__bF$buf0 ;
wire _5169_ ;
wire _5315__bF$buf1 ;
wire _5315__bF$buf2 ;
wire _5315__bF$buf3 ;
wire _5315__bF$buf4 ;
wire _83_ ;
wire _6950_ ;
wire _6530_ ;
wire _6110_ ;
wire _1089_ ;
wire _7735_ ;
wire _7315_ ;
wire _2870_ ;
wire _2450_ ;
wire _2030_ ;
wire _11733_ ;
wire _11313_ ;
wire _3655_ ;
wire _3235_ ;
wire _5801_ ;
wire _8693_ ;
wire _8273_ ;
wire _1721_ ;
wire _1301_ ;
wire _9898_ ;
wire _9478_ ;
wire _9058_ ;
wire _4193_ ;
wire _632_ ;
wire _212_ ;
wire _2926_ ;
wire _2506_ ;
wire _5398_ ;
wire _7964_ ;
wire _7544_ ;
wire _7124_ ;
wire _11542_ ;
wire _11122_ ;
wire _8749_ ;
wire _8329_ ;
wire _3884_ ;
wire _3464_ ;
wire _3044_ ;
wire _4669_ ;
wire _4249_ ;
wire _5610_ ;
wire _8082_ ;
wire _6815_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _9287_ ;
wire _10813_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _7773_ ;
wire _7353_ ;
wire _11771_ ;
wire _11351_ ;
wire _8978_ ;
wire _8558_ ;
wire _8138_ ;
wire _3693_ ;
wire _3273_ ;
wire _4898_ ;
wire _4478_ ;
wire _4058_ ;
wire _917_ ;
wire _6624_ ;
wire _6204_ ;
wire _9096_ ;
wire _10622_ ;
wire _10202_ ;
wire _670_ ;
wire _250_ ;
wire _7829_ ;
wire _7409_ ;
wire _2964_ ;
wire _2544_ ;
wire _2124_ ;
wire _11827_ ;
wire _11407_ ;
wire _3749_ ;
wire _3329_ ;
wire _7582_ ;
wire _7162_ ;
wire _11580_ ;
wire _11160_ ;
wire _8787_ ;
wire _8367_ ;
wire _3082_ ;
wire _1815_ ;
wire _4287_ ;
wire _726_ ;
wire _306_ ;
wire _6853_ ;
wire _6433_ ;
wire _6013_ ;
wire _10851_ ;
wire _10431_ ;
wire _10011_ ;
wire _7638_ ;
wire _7218_ ;
wire _2773_ ;
wire _2353_ ;
wire _11636_ ;
wire _11216_ ;
wire _3978_ ;
wire _3558_ ;
wire _3138_ ;
wire _7391_ ;
wire _5704_ ;
wire _8596_ ;
wire _8176_ ;
wire _5453__bF$buf0 ;
wire _5453__bF$buf1 ;
wire _5453__bF$buf2 ;
wire _5453__bF$buf3 ;
wire _5453__bF$buf4 ;
wire _5453__bF$buf5 ;
wire _6909_ ;
wire _1624_ ;
wire _1204_ ;
wire _4096_ ;
wire _10907_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2829_ ;
wire _2409_ ;
wire _6662_ ;
wire _6242_ ;
wire _10660_ ;
wire _10240_ ;
wire _7867_ ;
wire _7447_ ;
wire _7027_ ;
wire _2582_ ;
wire _2162_ ;
wire _11865_ ;
wire _11445_ ;
wire _11025_ ;
wire _3787_ ;
wire _3367_ ;
wire _5933_ ;
wire _5513_ ;
wire _6718_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _10716_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _6891_ ;
wire _6471_ ;
wire _6051_ ;
wire _7676_ ;
wire _7256_ ;
wire _2391_ ;
wire _11674_ ;
wire _11254_ ;
wire _3596_ ;
wire _3176_ ;
wire _9822_ ;
wire _9402_ ;
wire _2287__bF$buf0 ;
wire _2287__bF$buf1 ;
wire _2287__bF$buf2 ;
wire _1909_ ;
wire _2287__bF$buf3 ;
wire _5742_ ;
wire _5322_ ;
wire _6947_ ;
wire _6527_ ;
wire _6107_ ;
wire _1662_ ;
wire _1242_ ;
wire _10945_ ;
wire _10525_ ;
wire _10105_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2867_ ;
wire _2447_ ;
wire _2027_ ;
wire _6280_ ;
wire _7485_ ;
wire _7065_ ;
wire _11483_ ;
wire _11063_ ;
wire _9631_ ;
wire _9211_ ;
wire _1718_ ;
wire _5971_ ;
wire _5551_ ;
wire _5131_ ;
wire _629_ ;
wire _209_ ;
wire _6756_ ;
wire _6336_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _10754_ ;
wire _10334_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _8902_ ;
wire _11539_ ;
wire _11119_ ;
wire _4822_ ;
wire _4402_ ;
wire _7294_ ;
wire _11292_ ;
wire _5607_ ;
wire _8499_ ;
wire _8079_ ;
wire _9860_ ;
wire _9440_ ;
wire _9020_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _5780_ ;
wire _5360_ ;
wire _858_ ;
wire _438_ ;
wire _6985_ ;
wire _6565_ ;
wire _6145_ ;
wire _1280_ ;
wire _10983_ ;
wire _10563_ ;
wire _10143_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _8711_ ;
wire _11768_ ;
wire _11348_ ;
wire _9916_ ;
wire _4631_ ;
wire _4211_ ;
wire _5836_ ;
wire _5416_ ;
wire _1756_ ;
wire _1336_ ;
wire _10619_ ;
wire _667_ ;
wire _247_ ;
wire _3902_ ;
wire _6794_ ;
wire _6374_ ;
wire _10792_ ;
wire _10372_ ;
wire _7999_ ;
wire _7579_ ;
wire _7159_ ;
wire _2294_ ;
wire _8940_ ;
wire _8520_ ;
wire _8100_ ;
wire _11577_ ;
wire _11157_ ;
wire _3499_ ;
wire _3079_ ;
wire _9725_ ;
wire _9305_ ;
wire _4860_ ;
wire _4440_ ;
wire _4020_ ;
wire _5645_ ;
wire _5225_ ;
wire _4434__bF$buf0 ;
wire _4434__bF$buf1 ;
wire _4434__bF$buf2 ;
wire _4434__bF$buf3 ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _10848_ ;
wire _10428_ ;
wire _10008_ ;
wire _896_ ;
wire _476_ ;
wire _3711_ ;
wire _6183_ ;
wire _10181_ ;
wire _4916_ ;
wire _7388_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _11386_ ;
wire _9954_ ;
wire _9534_ ;
wire _9114_ ;
wire _5874_ ;
wire _5454_ ;
wire _5034_ ;
wire _6659_ ;
wire _6239_ ;
wire _1794_ ;
wire _1374_ ;
wire _7600_ ;
wire _10657_ ;
wire _10237_ ;
wire _285_ ;
wire _2999_ ;
wire _2579_ ;
wire _2159_ ;
wire _8805_ ;
wire _3940_ ;
wire _3520_ ;
wire _3100_ ;
wire _1_ ;
wire _4725_ ;
wire _4305_ ;
wire _7197_ ;
wire _11195_ ;
wire _9763_ ;
wire _9343_ ;
wire _5683_ ;
wire _5263_ ;
wire _6888_ ;
wire _6468_ ;
wire _6048_ ;
wire _1183_ ;
wire _10886_ ;
wire _10466_ ;
wire _10046_ ;
wire _2388_ ;
wire _8614_ ;
wire breg_14_bF$buf0 ;
wire breg_14_bF$buf1 ;
wire breg_14_bF$buf2 ;
wire breg_14_bF$buf3 ;
wire _9819_ ;
wire _4954_ ;
wire _4534_ ;
wire _4114_ ;
wire _5739_ ;
wire _5319_ ;
wire _9992_ ;
wire _9572_ ;
wire _9152_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _5492_ ;
wire _5072_ ;
wire _3805_ ;
wire _6697_ ;
wire _6277_ ;
wire _10695_ ;
wire _10275_ ;
wire _2197_ ;
wire _8843_ ;
wire _8423_ ;
wire _8003_ ;
wire _9628_ ;
wire _9208_ ;
wire _4763_ ;
wire _4343_ ;
wire _5968_ ;
wire _5548_ ;
wire _5128_ ;
wire _42_ ;
wire _9381_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _3614_ ;
wire _6086_ ;
wire _10084_ ;
wire _4819_ ;
wire _8652_ ;
wire _8232_ ;
wire _11289_ ;
wire _9857_ ;
wire _9437_ ;
wire _9017_ ;
wire _4992_ ;
wire _4572_ ;
wire _4152_ ;
wire _5777_ ;
wire _5357_ ;
wire _9190_ ;
wire _1697_ ;
wire _1277_ ;
wire _7923_ ;
wire _7503_ ;
wire _188_ ;
wire _11501_ ;
wire _8708_ ;
wire _3843_ ;
wire _3423_ ;
wire _3003_ ;
wire _4628_ ;
wire _4208_ ;
wire _8881_ ;
wire _8461_ ;
wire _8041_ ;
wire _11098_ ;
wire _9666_ ;
wire _9246_ ;
wire _4381_ ;
wire _820_ ;
wire _400_ ;
wire _5586_ ;
wire _5166_ ;
wire _80_ ;
wire _1086_ ;
wire _7732_ ;
wire _7312_ ;
wire _10789_ ;
wire _10369_ ;
wire _11730_ ;
wire _11310_ ;
wire _8937_ ;
wire _8517_ ;
wire _3652_ ;
wire _3232_ ;
wire _4857_ ;
wire _4437_ ;
wire _4017_ ;
wire _8690_ ;
wire _8270_ ;
wire _9895_ ;
wire _9475_ ;
wire _9055_ ;
wire _4190_ ;
wire _2923_ ;
wire _2503_ ;
wire _5395_ ;
wire _3708_ ;
wire _7961_ ;
wire _7541_ ;
wire _7121_ ;
wire _10598_ ;
wire _10178_ ;
wire _2586__bF$buf0 ;
wire _2586__bF$buf1 ;
wire _2586__bF$buf2 ;
wire _2586__bF$buf3 ;
wire _2586__bF$buf4 ;
wire _8746_ ;
wire _8326_ ;
wire _3881_ ;
wire _3461_ ;
wire _3041_ ;
wire _4666_ ;
wire _4246_ ;
wire _6812_ ;
wire _9284_ ;
wire _10810_ ;
wire _2732_ ;
wire _2312_ ;
wire _3937_ ;
wire _3517_ ;
wire _7770_ ;
wire _7350_ ;
wire _8975_ ;
wire _8555_ ;
wire _8135_ ;
wire _3690_ ;
wire _3270_ ;
wire _4895_ ;
wire _4475_ ;
wire _4055_ ;
wire _914_ ;
wire _6621_ ;
wire _6201_ ;
wire _9093_ ;
wire _7826_ ;
wire _7406_ ;
wire _2961_ ;
wire _2541_ ;
wire _2121_ ;
wire _11824_ ;
wire _11404_ ;
wire _3746_ ;
wire _3326_ ;
wire _8784_ ;
wire _8364_ ;
wire _1812_ ;
wire _9989_ ;
wire _9569_ ;
wire _9149_ ;
wire _4284_ ;
wire _723_ ;
wire _303_ ;
wire _5489_ ;
wire _5069_ ;
wire _6850_ ;
wire _6430_ ;
wire _6010_ ;
wire _7635_ ;
wire _7215_ ;
wire _2770_ ;
wire _2350_ ;
wire _11633_ ;
wire _11213_ ;
wire _3975_ ;
wire _3555_ ;
wire _3135_ ;
wire _5701_ ;
wire _8593_ ;
wire _8173_ ;
wire _39_ ;
wire _6906_ ;
wire _1621_ ;
wire _1201_ ;
wire _9798_ ;
wire _9378_ ;
wire _4093_ ;
wire _10904_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2826_ ;
wire _2406_ ;
wire _5298_ ;
wire _7864_ ;
wire _7444_ ;
wire _7024_ ;
wire _11862_ ;
wire _11442_ ;
wire _11022_ ;
wire _8649_ ;
wire _8229_ ;
wire _3784_ ;
wire _3364_ ;
wire _4989_ ;
wire _4569_ ;
wire _4149_ ;
wire _5930_ ;
wire _5510_ ;
wire _6715_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _9187_ ;
wire _10713_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire _7673_ ;
wire _7253_ ;
wire clk ;
wire _11671_ ;
wire _11251_ ;
wire _8878_ ;
wire _8458_ ;
wire _8038_ ;
wire _3593_ ;
wire _3173_ ;
wire _1906_ ;
wire _4798_ ;
wire _4378_ ;
wire _817_ ;
wire _77_ ;
wire _6944_ ;
wire _6524_ ;
wire _6104_ ;
wire _10942_ ;
wire _10522_ ;
wire _10102_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _7729_ ;
wire _7309_ ;
wire _2864_ ;
wire _2444_ ;
wire _2024_ ;
wire _11727_ ;
wire _11307_ ;
wire _3649_ ;
wire _3229_ ;
wire _7225__bF$buf0 ;
wire _7225__bF$buf1 ;
wire _7225__bF$buf2 ;
wire _7225__bF$buf3 ;
wire _7225__bF$buf4 ;
wire _7482_ ;
wire _7062_ ;
wire _11480_ ;
wire _11060_ ;
wire _8687_ ;
wire _8267_ ;
wire _1715_ ;
wire _4187_ ;
wire _626_ ;
wire _206_ ;
wire _6753_ ;
wire _6333_ ;
wire _10751_ ;
wire _10331_ ;
wire _7958_ ;
wire _7538_ ;
wire _7118_ ;
wire _2673_ ;
wire _2253_ ;
wire areg_16_bF$buf0 ;
wire areg_16_bF$buf1 ;
wire areg_16_bF$buf2 ;
wire areg_16_bF$buf3 ;
wire areg_16_bF$buf4 ;
wire areg_16_bF$buf5 ;
wire _11536_ ;
wire _11116_ ;
wire _3878_ ;
wire _3458_ ;
wire _3038_ ;
wire _7291_ ;
wire _5604_ ;
wire _8496_ ;
wire _8076_ ;
wire _6809_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _10807_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _6982_ ;
wire _6562_ ;
wire _6142_ ;
wire _10980_ ;
wire _10560_ ;
wire _10140_ ;
wire _7767_ ;
wire _7347_ ;
wire _2482_ ;
wire _2062_ ;
wire _11765_ ;
wire _11345_ ;
wire _3687_ ;
wire _3267_ ;
wire _9913_ ;
wire _5833_ ;
wire _5413_ ;
wire _6618_ ;
wire _1753_ ;
wire _1333_ ;
wire _10616_ ;
wire _664_ ;
wire _244_ ;
wire _2958_ ;
wire _2538_ ;
wire _2118_ ;
wire _6791_ ;
wire _6371_ ;
wire _7996_ ;
wire _7576_ ;
wire _7156_ ;
wire _2291_ ;
wire _11574_ ;
wire _11154_ ;
wire _3496_ ;
wire _3076_ ;
wire _9722_ ;
wire _9302_ ;
wire _1809_ ;
wire _5642_ ;
wire _5222_ ;
wire _6847_ ;
wire _6427_ ;
wire _6007_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _10845_ ;
wire _10425_ ;
wire _10005_ ;
wire _893_ ;
wire _473_ ;
wire _2767_ ;
wire _2347_ ;
wire _6180_ ;
wire _4913_ ;
wire _7385_ ;
wire _11383_ ;
wire _9951_ ;
wire _9531_ ;
wire _9111_ ;
wire _1618_ ;
wire _5871_ ;
wire _5451_ ;
wire _5031_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _6656_ ;
wire _6236_ ;
wire _1791_ ;
wire _1371_ ;
wire _10654_ ;
wire _10234_ ;
wire _282_ ;
wire _2996_ ;
wire _2576_ ;
wire _2156_ ;
wire _8802_ ;
wire _11859_ ;
wire _11439_ ;
wire _11019_ ;
wire _4722_ ;
wire _4302_ ;
wire _7194_ ;
wire _11192_ ;
wire _5927_ ;
wire _5507_ ;
wire _8399_ ;
wire _9760_ ;
wire _9340_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _5680_ ;
wire _5260_ ;
wire _758_ ;
wire _338_ ;
wire _6885_ ;
wire _6465_ ;
wire _6045_ ;
wire _1180_ ;
wire _10883_ ;
wire _10463_ ;
wire _10043_ ;
wire _2385_ ;
wire _8611_ ;
wire _11668_ ;
wire _11248_ ;
wire _9816_ ;
wire _4951_ ;
wire _4531_ ;
wire _4111_ ;
wire _5736_ ;
wire _5316_ ;
wire _1656_ ;
wire _1236_ ;
wire _10939_ ;
wire _10519_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _3802_ ;
wire _6694_ ;
wire _6274_ ;
wire _10692_ ;
wire _10272_ ;
wire _7899_ ;
wire _7479_ ;
wire _7059_ ;
wire _2194_ ;
wire _8840_ ;
wire _8420_ ;
wire _8000_ ;
wire _11897_ ;
wire _11477_ ;
wire _11057_ ;
wire _3399_ ;
wire _9625_ ;
wire _9205_ ;
wire _4760_ ;
wire _4340_ ;
wire _5965_ ;
wire _5545_ ;
wire _5125_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _10748_ ;
wire _10328_ ;
wire _796_ ;
wire _376_ ;
wire _3611_ ;
wire _6083_ ;
wire _10081_ ;
wire _4816_ ;
wire _7288_ ;
wire _11286_ ;
wire _9854_ ;
wire _9434_ ;
wire _9014_ ;
wire _5774_ ;
wire _5354_ ;
wire _6979_ ;
wire _6559_ ;
wire _6139_ ;
wire _1694_ ;
wire _1274_ ;
wire _7920_ ;
wire _7500_ ;
wire _10977_ ;
wire _10557_ ;
wire _10137_ ;
wire _185_ ;
wire _2899_ ;
wire _2479_ ;
wire _2059_ ;
wire _8705_ ;
wire _3840_ ;
wire _3420_ ;
wire _3000_ ;
wire _4625_ ;
wire _4205_ ;
wire _7097_ ;
wire _11095_ ;
wire _9663_ ;
wire _9243_ ;
wire _5583_ ;
wire _5163_ ;
wire _6788_ ;
wire _6368_ ;
wire _1083_ ;
wire _10786_ ;
wire _10366_ ;
wire _2288_ ;
wire _8934_ ;
wire _8514_ ;
wire _9719_ ;
wire _4854_ ;
wire _4434_ ;
wire _4014_ ;
wire _5639_ ;
wire _5219_ ;
wire _9892_ ;
wire _9472_ ;
wire _9052_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2920_ ;
wire _2500_ ;
wire _5392_ ;
wire _3705_ ;
wire _6597_ ;
wire _6177_ ;
wire _10595_ ;
wire _10175_ ;
wire _2097_ ;
wire _8743_ ;
wire _8323_ ;
wire _9948_ ;
wire _9528_ ;
wire _9108_ ;
wire _4663_ ;
wire _4243_ ;
wire _5868_ ;
wire _5448_ ;
wire _5028_ ;
wire _9281_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _3934_ ;
wire _3514_ ;
wire _4719_ ;
wire _8972_ ;
wire _8552_ ;
wire _8132_ ;
wire _11189_ ;
wire _9757_ ;
wire _9337_ ;
wire _4892_ ;
wire _4472_ ;
wire _4052_ ;
wire _911_ ;
wire _5677_ ;
wire _5257_ ;
wire _9090_ ;
wire _1597_ ;
wire _1177_ ;
wire _7823_ ;
wire _7403_ ;
wire _11821_ ;
wire _11401_ ;
wire _8608_ ;
wire _3743_ ;
wire _3323_ ;
wire _4948_ ;
wire _4528_ ;
wire _4108_ ;
wire _8781_ ;
wire _8361_ ;
wire _9986_ ;
wire _9566_ ;
wire _9146_ ;
wire _4281_ ;
wire _720_ ;
wire _300_ ;
wire _5486_ ;
wire _5066_ ;
wire _7632_ ;
wire _7212_ ;
wire _10689_ ;
wire _10269_ ;
wire _11630_ ;
wire _11210_ ;
wire _8837_ ;
wire _8417_ ;
wire _3972_ ;
wire _3552_ ;
wire _3132_ ;
wire _4757_ ;
wire _4337_ ;
wire _8590_ ;
wire _8170_ ;
wire _36_ ;
wire _6903_ ;
wire _9795_ ;
wire _9375_ ;
wire _4090_ ;
wire _10901_ ;
wire _2823_ ;
wire _2403_ ;
wire _5295_ ;
wire _3608_ ;
wire _7861_ ;
wire _7441_ ;
wire _7021_ ;
wire _10498_ ;
wire _10078_ ;
wire _8646_ ;
wire _8226_ ;
wire _3781_ ;
wire _3361_ ;
wire _4986_ ;
wire _4566_ ;
wire _4146_ ;
wire _6712_ ;
wire _9184_ ;
wire _10710_ ;
wire _7917_ ;
wire _2632_ ;
wire _2212_ ;
wire _3837_ ;
wire _3417_ ;
wire _7670_ ;
wire _7250_ ;
wire _8875_ ;
wire _8455_ ;
wire _8035_ ;
wire _3590_ ;
wire _3170_ ;
wire _1903_ ;
wire _4795_ ;
wire _4375_ ;
wire _814_ ;
wire _74_ ;
wire _6941_ ;
wire _6521_ ;
wire _6101_ ;
wire _7726_ ;
wire _7306_ ;
wire _2861_ ;
wire _2441_ ;
wire _2021_ ;
wire _11724_ ;
wire _11304_ ;
wire _3646_ ;
wire _3226_ ;
wire _2376__bF$buf0 ;
wire _2376__bF$buf1 ;
wire _2376__bF$buf2 ;
wire _2376__bF$buf3 ;
wire _8684_ ;
wire _8264_ ;
wire _1712_ ;
wire _9889_ ;
wire _9469_ ;
wire _9049_ ;
wire _4184_ ;
wire _623_ ;
wire _203_ ;
wire _2917_ ;
wire _5389_ ;
wire _6750_ ;
wire _6330_ ;
wire _7955_ ;
wire _7535_ ;
wire _7115_ ;
wire _2670_ ;
wire _2250_ ;
wire _11533_ ;
wire _11113_ ;
wire _3875_ ;
wire _3455_ ;
wire _3035_ ;
wire _5601_ ;
wire _8493_ ;
wire _8073_ ;
wire _6806_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _9698_ ;
wire _9278_ ;
wire _10804_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _5198_ ;
wire _7764_ ;
wire _7344_ ;
wire _11762_ ;
wire _11342_ ;
wire _8969_ ;
wire _8549_ ;
wire _8129_ ;
wire _3684_ ;
wire _3264_ ;
wire _9910_ ;
wire _4889_ ;
wire _4469_ ;
wire _4049_ ;
wire _5830_ ;
wire _5410_ ;
wire _908_ ;
wire _6615_ ;
wire _1750_ ;
wire _1330_ ;
wire _9087_ ;
wire _10613_ ;
wire _661_ ;
wire _241_ ;
wire _2955_ ;
wire _2535_ ;
wire _2115_ ;
wire _11818_ ;
wire _7993_ ;
wire _7573_ ;
wire _7153_ ;
wire _11571_ ;
wire _11151_ ;
wire _8778_ ;
wire _8358_ ;
wire _3493_ ;
wire _3073_ ;
wire _1806_ ;
wire _4698_ ;
wire _4278_ ;
wire _717_ ;
wire _6844_ ;
wire _6424_ ;
wire _6004_ ;
wire _10842_ ;
wire _10422_ ;
wire _10002_ ;
wire _890_ ;
wire _470_ ;
wire _7629_ ;
wire _7209_ ;
wire _2764_ ;
wire _2344_ ;
wire _11627_ ;
wire _11207_ ;
wire _3969_ ;
wire _3549_ ;
wire _3129_ ;
wire _4910_ ;
wire areg_27_bF$buf0 ;
wire areg_27_bF$buf1 ;
wire areg_27_bF$buf2 ;
wire areg_27_bF$buf3 ;
wire areg_27_bF$buf4 ;
wire areg_27_bF$buf5 ;
wire _7382_ ;
wire _11380_ ;
wire _8587_ ;
wire _8167_ ;
wire _1615_ ;
wire _4087_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _6653_ ;
wire _6233_ ;
wire _10651_ ;
wire _10231_ ;
wire _7858_ ;
wire _7438_ ;
wire _7018_ ;
wire _2993_ ;
wire _2573_ ;
wire _2153_ ;
wire _11856_ ;
wire _11436_ ;
wire _11016_ ;
wire _3778_ ;
wire _3358_ ;
wire _7191_ ;
wire _5924_ ;
wire _5504_ ;
wire _8396_ ;
wire _6709_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _10707_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _6882_ ;
wire _6462_ ;
wire _6042_ ;
wire _10880_ ;
wire _10460_ ;
wire _10040_ ;
wire _7667_ ;
wire _7247_ ;
wire _2382_ ;
wire _11665_ ;
wire _11245_ ;
wire _3587_ ;
wire _3167_ ;
wire _9813_ ;
wire _5733_ ;
wire _5313_ ;
wire _6938_ ;
wire _6518_ ;
wire _1653_ ;
wire _1233_ ;
wire _10936_ ;
wire _10516_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2858_ ;
wire _2438_ ;
wire _2018_ ;
wire _6691_ ;
wire _6271_ ;
wire _7896_ ;
wire _7476_ ;
wire _7056_ ;
wire _2191_ ;
wire _11894_ ;
wire _11474_ ;
wire _11054_ ;
wire _3396_ ;
wire _9622_ ;
wire _9202_ ;
wire _1709_ ;
wire _5962_ ;
wire _5542_ ;
wire _5122_ ;
wire _6747_ ;
wire _6327_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _10745_ ;
wire _10325_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _6080_ ;
wire _4813_ ;
wire _7285_ ;
wire _11283_ ;
wire _9851_ ;
wire _9431_ ;
wire _9011_ ;
wire areg_9_bF$buf0 ;
wire areg_9_bF$buf1 ;
wire areg_9_bF$buf2 ;
wire areg_9_bF$buf3 ;
wire areg_9_bF$buf4 ;
wire _1938_ ;
wire _1518_ ;
wire _5771_ ;
wire _5351_ ;
wire _849_ ;
wire _429_ ;
wire _6976_ ;
wire _6556_ ;
wire _6136_ ;
wire _1691_ ;
wire _1271_ ;
wire _10974_ ;
wire _10554_ ;
wire _10134_ ;
wire _182_ ;
wire _2896_ ;
wire _2476_ ;
wire _2056_ ;
wire _8702_ ;
wire _11759_ ;
wire _11339_ ;
wire _9907_ ;
wire _4622_ ;
wire _4202_ ;
wire _7094_ ;
wire _11092_ ;
wire _5827_ ;
wire _5407_ ;
wire _8299_ ;
wire _9660_ ;
wire _9240_ ;
wire _1747_ ;
wire _1327_ ;
wire _5580_ ;
wire _5160_ ;
wire _658_ ;
wire _238_ ;
wire _6785_ ;
wire _6365_ ;
wire _1080_ ;
wire _10783_ ;
wire _10363_ ;
wire _2285_ ;
wire _8931_ ;
wire _8511_ ;
wire _11568_ ;
wire _11148_ ;
wire _9716_ ;
wire _4851_ ;
wire _4431_ ;
wire _4011_ ;
wire _5636_ ;
wire _5216_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _10839_ ;
wire _10419_ ;
wire _887_ ;
wire _467_ ;
wire _3702_ ;
wire _6594_ ;
wire _6174_ ;
wire _10592_ ;
wire _10172_ ;
wire _4907_ ;
wire _7799_ ;
wire _7379_ ;
wire _2094_ ;
wire _8740_ ;
wire _8320_ ;
wire _11797_ ;
wire _11377_ ;
wire _3299_ ;
wire _9945_ ;
wire _9525_ ;
wire _9105_ ;
wire _4660_ ;
wire _4240_ ;
wire areg_11_bF$buf0 ;
wire areg_11_bF$buf1 ;
wire areg_11_bF$buf2 ;
wire _5865_ ;
wire areg_11_bF$buf3 ;
wire _5445_ ;
wire areg_11_bF$buf4 ;
wire _5025_ ;
wire _1785_ ;
wire _1365_ ;
wire _10648_ ;
wire _10228_ ;
wire _696_ ;
wire _276_ ;
wire _3931_ ;
wire _3511_ ;
wire _4716_ ;
wire _7188_ ;
wire _11186_ ;
wire _9754_ ;
wire _9334_ ;
wire _5674_ ;
wire _5254_ ;
wire _6879_ ;
wire _6459_ ;
wire _6039_ ;
wire _1594_ ;
wire _1174_ ;
wire _7820_ ;
wire _7400_ ;
wire _10877_ ;
wire _10457_ ;
wire _10037_ ;
wire _2799_ ;
wire _2379_ ;
wire _8605_ ;
wire _3740_ ;
wire _3320_ ;
wire _4945_ ;
wire _4525_ ;
wire _4105_ ;
wire _9983_ ;
wire _9563_ ;
wire _9143_ ;
wire _5483_ ;
wire _5063_ ;
wire _6688_ ;
wire _6268_ ;
wire _10686_ ;
wire _10266_ ;
wire _2188_ ;
wire _8834_ ;
wire _8414_ ;
wire _9619_ ;
wire _4754_ ;
wire _4334_ ;
wire _5959_ ;
wire _5539_ ;
wire _5119_ ;
wire _33_ ;
wire _6900_ ;
wire _9792_ ;
wire _9372_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2820_ ;
wire _2400_ ;
wire _5292_ ;
wire _3605_ ;
wire _6497_ ;
wire _6077_ ;
wire _10495_ ;
wire _10075_ ;
wire _8643_ ;
wire _8223_ ;
wire _9848_ ;
wire _9428_ ;
wire _9008_ ;
wire _4983_ ;
wire _4563_ ;
wire _4143_ ;
wire _5768_ ;
wire _5348_ ;
wire _9181_ ;
wire _1688_ ;
wire _1268_ ;
wire _7914_ ;
wire _599_ ;
wire _179_ ;
wire _3834_ ;
wire _3414_ ;
wire _4619_ ;
wire _8872_ ;
wire _8452_ ;
wire _8032_ ;
wire _11089_ ;
wire _1900_ ;
wire _9657_ ;
wire _9237_ ;
wire _4792_ ;
wire _4372_ ;
wire _811_ ;
wire _5997_ ;
wire _5577_ ;
wire _5157_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _7723_ ;
wire _7303_ ;
wire _11721_ ;
wire _11301_ ;
wire _8928_ ;
wire _8508_ ;
wire _3643_ ;
wire _3223_ ;
wire _4848_ ;
wire _4428_ ;
wire _4008_ ;
wire _8681_ ;
wire _8261_ ;
wire _9886_ ;
wire _9466_ ;
wire _9046_ ;
wire _4181_ ;
wire _620_ ;
wire _200_ ;
wire _2914_ ;
wire _5386_ ;
wire _7952_ ;
wire _7532_ ;
wire _7112_ ;
wire _10589_ ;
wire _10169_ ;
wire _11530_ ;
wire _11110_ ;
wire _8737_ ;
wire _8317_ ;
wire _3872_ ;
wire _3452_ ;
wire _3032_ ;
wire _4657_ ;
wire _4237_ ;
wire _8490_ ;
wire _8070_ ;
wire _6803_ ;
wire _9695_ ;
wire _9275_ ;
wire _10801_ ;
wire _2723_ ;
wire _2303_ ;
wire _5195_ ;
wire _3928_ ;
wire _3508_ ;
wire _7761_ ;
wire _7341_ ;
wire _10398_ ;
wire _8966_ ;
wire _8546_ ;
wire _8126_ ;
wire _3681_ ;
wire _3261_ ;
wire _4886_ ;
wire _4466_ ;
wire _4046_ ;
wire _905_ ;
wire _6612_ ;
wire _9084_ ;
wire _10610_ ;
wire _7817_ ;
wire _2952_ ;
wire _2532_ ;
wire _2112_ ;
wire _11815_ ;
wire _3737_ ;
wire _3317_ ;
wire breg_29_bF$buf0 ;
wire breg_29_bF$buf1 ;
wire breg_29_bF$buf2 ;
wire breg_29_bF$buf3 ;
wire breg_29_bF$buf4 ;
wire _7990_ ;
wire _7570_ ;
wire _7150_ ;
wire _8775_ ;
wire _8355_ ;
wire _3490_ ;
wire _3070_ ;
wire _1803_ ;
wire _4695_ ;
wire _4275_ ;
wire _714_ ;
wire _6841_ ;
wire _6421_ ;
wire _6001_ ;
wire breg_7_bF$buf0 ;
wire breg_7_bF$buf1 ;
wire breg_7_bF$buf2 ;
wire breg_7_bF$buf3 ;
wire breg_7_bF$buf4 ;
wire breg_7_bF$buf5 ;
wire _7626_ ;
wire _7206_ ;
wire _2761_ ;
wire _2341_ ;
wire _11624_ ;
wire _11204_ ;
wire _3966_ ;
wire _3546_ ;
wire _3126_ ;
wire _8584_ ;
wire _8164_ ;
wire _1612_ ;
wire _9789_ ;
wire _9369_ ;
wire _4084_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2817_ ;
wire _5289_ ;
wire _6650_ ;
wire _6230_ ;
wire _7855_ ;
wire _7435_ ;
wire _7015_ ;
wire _2990_ ;
wire _2570_ ;
wire _2150_ ;
wire _11853_ ;
wire _11433_ ;
wire _11013_ ;
wire _3775_ ;
wire _3355_ ;
wire _5921_ ;
wire _5501_ ;
wire _8393_ ;
wire _6706_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _9598_ ;
wire _9178_ ;
wire _10704_ ;
wire _5190__bF$buf0 ;
wire _5190__bF$buf1 ;
wire _5190__bF$buf2 ;
wire _5190__bF$buf3 ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _5098_ ;
wire [63:0] _11909_ ;
wire _7664_ ;
wire _7244_ ;
wire _11662_ ;
wire _11242_ ;
wire _8869_ ;
wire _8449_ ;
wire _8029_ ;
wire _3584_ ;
wire _3164_ ;
wire _9810_ ;
wire _4789_ ;
wire _4369_ ;
wire _5730_ ;
wire _5310_ ;
wire _808_ ;
wire _68_ ;
wire _6935_ ;
wire _6515_ ;
wire _1650_ ;
wire _1230_ ;
wire _10933_ ;
wire _10513_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2855_ ;
wire _2435_ ;
wire _2015_ ;
wire _11718_ ;
wire _7893_ ;
wire _7473_ ;
wire _7053_ ;
wire _11891_ ;
wire _11471_ ;
wire _11051_ ;
wire _8678_ ;
wire _8258_ ;
wire _3393_ ;
wire _1706_ ;
wire _4598_ ;
wire _4178_ ;
wire _617_ ;
wire _6744_ ;
wire _6324_ ;
wire _10742_ ;
wire _10322_ ;
wire _790_ ;
wire _370_ ;
wire _7949_ ;
wire _7529_ ;
wire _7109_ ;
wire _2664_ ;
wire _2244_ ;
wire _11527_ ;
wire _11107_ ;
wire _3869_ ;
wire _3449_ ;
wire _3029_ ;
wire _4810_ ;
wire _7282_ ;
wire _11280_ ;
wire _8487_ ;
wire _8067_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _6973_ ;
wire _6553_ ;
wire _6133_ ;
wire _10971_ ;
wire _10551_ ;
wire _10131_ ;
wire _7758_ ;
wire _7338_ ;
wire _2893_ ;
wire _2473_ ;
wire _2053_ ;
wire _11756_ ;
wire _11336_ ;
wire _3678_ ;
wire _3258_ ;
wire _9904_ ;
wire _7091_ ;
wire _5824_ ;
wire _5404_ ;
wire _8296_ ;
wire _6609_ ;
wire _1744_ ;
wire _1324_ ;
wire _10607_ ;
wire _655_ ;
wire _235_ ;
wire _2949_ ;
wire _2529_ ;
wire _2109_ ;
wire _6782_ ;
wire _6362_ ;
wire _10780_ ;
wire _10360_ ;
wire _7987_ ;
wire _7567_ ;
wire _7147_ ;
wire _2282_ ;
wire _11565_ ;
wire _11145_ ;
wire _3487_ ;
wire _3067_ ;
wire _9713_ ;
wire _5633_ ;
wire _5213_ ;
wire _6838_ ;
wire _6418_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _10836_ ;
wire _10416_ ;
wire _884_ ;
wire _464_ ;
wire _2758_ ;
wire _2338_ ;
wire _6591_ ;
wire _6171_ ;
wire _4904_ ;
wire _7796_ ;
wire _7376_ ;
wire _2091_ ;
wire _11794_ ;
wire _11374_ ;
wire _3296_ ;
wire _9942_ ;
wire _9522_ ;
wire _9102_ ;
wire _1609_ ;
wire _5862_ ;
wire _5442_ ;
wire _5022_ ;
wire _6647_ ;
wire _6227_ ;
wire _1782_ ;
wire _1362_ ;
wire _10645_ ;
wire _10225_ ;
wire _693_ ;
wire _273_ ;
wire _2987_ ;
wire _2567_ ;
wire _2147_ ;
wire _4713_ ;
wire _7185_ ;
wire _11183_ ;
wire _5918_ ;
wire _9751_ ;
wire _9331_ ;
wire _1838_ ;
wire _1418_ ;
wire _5671_ ;
wire _5251_ ;
wire _749_ ;
wire _329_ ;
wire _6876_ ;
wire _6456_ ;
wire _6036_ ;
wire _1591_ ;
wire _1171_ ;
wire _10874_ ;
wire _10454_ ;
wire _10034_ ;
wire _2796_ ;
wire _2376_ ;
wire _8602_ ;
wire _11659_ ;
wire _11239_ ;
wire _9807_ ;
wire _4942_ ;
wire _4522_ ;
wire _4102_ ;
wire _5727_ ;
wire _5307_ ;
wire _8199_ ;
wire _9980_ ;
wire _9560_ ;
wire _9140_ ;
wire _1647_ ;
wire _1227_ ;
wire _5480_ ;
wire _5060_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _6685_ ;
wire _6265_ ;
wire _10683_ ;
wire _10263_ ;
wire _2185_ ;
wire _8831_ ;
wire _8411_ ;
wire _11888_ ;
wire _11468_ ;
wire _11048_ ;
wire _9616_ ;
wire _4751_ ;
wire _4331_ ;
wire _5956_ ;
wire _5536_ ;
wire _5116_ ;
wire _30_ ;
wire areg_22_bF$buf0 ;
wire _1876_ ;
wire areg_22_bF$buf1 ;
wire _1456_ ;
wire areg_22_bF$buf2 ;
wire _1036_ ;
wire areg_22_bF$buf3 ;
wire areg_22_bF$buf4 ;
wire _10739_ ;
wire _10319_ ;
wire _787_ ;
wire _367_ ;
wire _3602_ ;
wire _6494_ ;
wire _6074_ ;
wire _10492_ ;
wire _10072_ ;
wire _4807_ ;
wire _7699_ ;
wire _7279_ ;
wire _8640_ ;
wire _8220_ ;
wire _11697_ ;
wire _11277_ ;
wire _3199_ ;
wire _9845_ ;
wire _9425_ ;
wire _9005_ ;
wire _4980_ ;
wire _4560_ ;
wire _4140_ ;
wire _5765_ ;
wire _5345_ ;
wire _1685_ ;
wire _1265_ ;
wire _7911_ ;
wire _10968_ ;
wire _10548_ ;
wire _10128_ ;
wire _596_ ;
wire _176_ ;
wire _3831_ ;
wire _3411_ ;
wire _4616_ ;
wire _7088_ ;
wire _11086_ ;
wire _9654_ ;
wire _9234_ ;
wire _5994_ ;
wire _5574_ ;
wire _5154_ ;
wire _6779_ ;
wire _6359_ ;
wire _1494_ ;
wire _1074_ ;
wire _7720_ ;
wire _7300_ ;
wire _10777_ ;
wire _10357_ ;
wire _2699_ ;
wire _2279_ ;
wire _8925_ ;
wire _8505_ ;
wire _3640_ ;
wire _3220_ ;
wire _4845_ ;
wire _4425_ ;
wire _4005_ ;
wire _9883_ ;
wire _9463_ ;
wire _9043_ ;
wire _2911_ ;
wire _5383_ ;
wire _6588_ ;
wire _6168_ ;
wire _10586_ ;
wire _10166_ ;
wire _2088_ ;
wire _8734_ ;
wire _8314_ ;
wire _9939_ ;
wire _9519_ ;
wire _4654_ ;
wire _4234_ ;
wire _5859_ ;
wire _5439_ ;
wire _5019_ ;
wire _6800_ ;
wire _9692_ ;
wire _9272_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire _5192_ ;
wire _3925_ ;
wire _3505_ ;
wire _6397_ ;
wire areg_4_bF$buf0 ;
wire areg_4_bF$buf1 ;
wire areg_4_bF$buf2 ;
wire areg_4_bF$buf3 ;
wire areg_4_bF$buf4 ;
wire _10395_ ;
wire _8963_ ;
wire _8543_ ;
wire _8123_ ;
wire _9748_ ;
wire _9328_ ;
wire _4883_ ;
wire _4463_ ;
wire _4043_ ;
wire _902_ ;
wire _5668_ ;
wire _5248_ ;
wire _9081_ ;
wire _1588_ ;
wire _1168_ ;
wire _7814_ ;
wire _499_ ;
wire _11812_ ;
wire _3734_ ;
wire _3314_ ;
wire _4939_ ;
wire _4519_ ;
wire _8772_ ;
wire _8352_ ;
wire _1800_ ;
wire _9977_ ;
wire _9557_ ;
wire _9137_ ;
wire _4692_ ;
wire _4272_ ;
wire _711_ ;
wire _5897_ ;
wire _5477_ ;
wire _5057_ ;
wire _1397_ ;
wire _7623_ ;
wire _7203_ ;
wire _11621_ ;
wire _11201_ ;
wire _8828_ ;
wire _8408_ ;
wire _3963_ ;
wire _3543_ ;
wire _3123_ ;
wire _4748_ ;
wire _4328_ ;
wire _8581_ ;
wire _8161_ ;
wire _27_ ;
wire _9786_ ;
wire _9366_ ;
wire _4081_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2814_ ;
wire _5286_ ;
wire _7852_ ;
wire _7432_ ;
wire _7012_ ;
wire _10489_ ;
wire _10069_ ;
wire _11850_ ;
wire _11430_ ;
wire _11010_ ;
wire _8637_ ;
wire _8217_ ;
wire _3772_ ;
wire _3352_ ;
wire _4977_ ;
wire _4557_ ;
wire _4137_ ;
wire _8390_ ;
wire _6703_ ;
wire _9595_ ;
wire _9175_ ;
wire _10701_ ;
wire _7908_ ;
wire _2623_ ;
wire _2203_ ;
wire _5095_ ;
wire _11906_ ;
wire _3828_ ;
wire _3408_ ;
wire _7661_ ;
wire _7241_ ;
wire _10298_ ;
wire _8866_ ;
wire _8446_ ;
wire _8026_ ;
wire _3581_ ;
wire _3161_ ;
wire _4786_ ;
wire _4366_ ;
wire _805_ ;
wire _65_ ;
wire _6932_ ;
wire _6512_ ;
wire _10930_ ;
wire _10510_ ;
wire _7717_ ;
wire _2852_ ;
wire _2432_ ;
wire _2012_ ;
wire _11715_ ;
wire _3637_ ;
wire _3217_ ;
wire _7890_ ;
wire _7470_ ;
wire _7050_ ;
wire _8675_ ;
wire _8255_ ;
wire _3390_ ;
wire _1703_ ;
wire _4595_ ;
wire _4175_ ;
wire _614_ ;
wire _2908_ ;
wire _6741_ ;
wire _6321_ ;
wire _7946_ ;
wire _7526_ ;
wire _7106_ ;
wire _2661_ ;
wire _2241_ ;
wire _11524_ ;
wire _11104_ ;
wire _3866_ ;
wire _3446_ ;
wire _3026_ ;
wire _8484_ ;
wire _8064_ ;
wire _1932_ ;
wire _1512_ ;
wire _9689_ ;
wire _9269_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _5189_ ;
wire _6970_ ;
wire _6550_ ;
wire _6130_ ;
wire _7755_ ;
wire _7335_ ;
wire _2890_ ;
wire _2470_ ;
wire _2050_ ;
wire _11753_ ;
wire _11333_ ;
wire _3675_ ;
wire _3255_ ;
wire _9901_ ;
wire _5821_ ;
wire _5401_ ;
wire _8293_ ;
wire _6606_ ;
wire _1741_ ;
wire _1321_ ;
wire _9498_ ;
wire _9078_ ;
wire _10604_ ;
wire _652_ ;
wire _232_ ;
wire _2946_ ;
wire _2526_ ;
wire _2106_ ;
wire _11809_ ;
wire _7984_ ;
wire _7564_ ;
wire _7144_ ;
wire _11562_ ;
wire _11142_ ;
wire _8769_ ;
wire _8349_ ;
wire _3484_ ;
wire _3064_ ;
wire _9710_ ;
wire _4689_ ;
wire _4269_ ;
wire _5630_ ;
wire _5210_ ;
wire _708_ ;
wire _6835_ ;
wire _6415_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _10833_ ;
wire _10413_ ;
wire _881_ ;
wire _461_ ;
wire _2755_ ;
wire _2335_ ;
wire _11618_ ;
wire _4901_ ;
wire _7793_ ;
wire _7373_ ;
wire _11791_ ;
wire _11371_ ;
wire _8998_ ;
wire _8578_ ;
wire _8158_ ;
wire _3293_ ;
wire _1606_ ;
wire _4498_ ;
wire _4078_ ;
wire _937_ ;
wire _517_ ;
wire _6644_ ;
wire _6224_ ;
wire _10642_ ;
wire _10222_ ;
wire _690_ ;
wire _270_ ;
wire _7849_ ;
wire _7429_ ;
wire _7009_ ;
wire _2984_ ;
wire _2564_ ;
wire _2144_ ;
wire _11847_ ;
wire _11427_ ;
wire _11007_ ;
wire _3769_ ;
wire _3349_ ;
wire _4710_ ;
wire _7182_ ;
wire _11180_ ;
wire _5915_ ;
wire _8387_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _6873_ ;
wire _6453_ ;
wire _6033_ ;
wire _10871_ ;
wire _10451_ ;
wire _10031_ ;
wire _7658_ ;
wire _7238_ ;
wire _2793_ ;
wire _2373_ ;
wire _11656_ ;
wire _11236_ ;
wire _3998_ ;
wire _3578_ ;
wire _3158_ ;
wire _9804_ ;
wire _5724_ ;
wire _5304_ ;
wire _8196_ ;
wire _6929_ ;
wire _6509_ ;
wire breg_24_bF$buf0 ;
wire _1644_ ;
wire breg_24_bF$buf1 ;
wire _1224_ ;
wire breg_24_bF$buf2 ;
wire breg_24_bF$buf3 ;
wire breg_24_bF$buf4 ;
wire breg_24_bF$buf5 ;
wire _10927_ ;
wire _10507_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2849_ ;
wire _2429_ ;
wire _2009_ ;
wire _6682_ ;
wire _6262_ ;
wire _10680_ ;
wire _10260_ ;
wire _7887_ ;
wire _7467_ ;
wire _7047_ ;
wire _2182_ ;
wire _11885_ ;
wire _11465_ ;
wire _11045_ ;
wire _3387_ ;
wire breg_2_bF$buf0 ;
wire _9613_ ;
wire breg_2_bF$buf1 ;
wire breg_2_bF$buf2 ;
wire breg_2_bF$buf3 ;
wire breg_2_bF$buf4 ;
wire _5953_ ;
wire _5533_ ;
wire _5113_ ;
wire _6738_ ;
wire _6318_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _10736_ ;
wire _10316_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _6491_ ;
wire _6071_ ;
wire _4804_ ;
wire _7696_ ;
wire _7276_ ;
wire _11694_ ;
wire _11274_ ;
wire _3196_ ;
wire _9842_ ;
wire _9422_ ;
wire _9002_ ;
wire _1929_ ;
wire _1509_ ;
wire _5762_ ;
wire _5342_ ;
wire _6967_ ;
wire _6547_ ;
wire _6127_ ;
wire _1682_ ;
wire _1262_ ;
wire _10965_ ;
wire _10545_ ;
wire _10125_ ;
wire _593_ ;
wire _173_ ;
wire _2887_ ;
wire _2467_ ;
wire _2047_ ;
wire _4613_ ;
wire _7085_ ;
wire _11083_ ;
wire _5818_ ;
wire _9651_ ;
wire _9231_ ;
wire _1738_ ;
wire _1318_ ;
wire _5991_ ;
wire _5571_ ;
wire _5151_ ;
wire _649_ ;
wire _229_ ;
wire _6776_ ;
wire _6356_ ;
wire _1491_ ;
wire _1071_ ;
wire _10774_ ;
wire _10354_ ;
wire _2696_ ;
wire _2276_ ;
wire _8922_ ;
wire _8502_ ;
wire _11559_ ;
wire _11139_ ;
wire _9707_ ;
wire _4842_ ;
wire _4422_ ;
wire _4002_ ;
wire _5627_ ;
wire _5207_ ;
wire _8099_ ;
wire _9880_ ;
wire _9460_ ;
wire _9040_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _5380_ ;
wire _878_ ;
wire _458_ ;
wire _6585_ ;
wire _6165_ ;
wire _10583_ ;
wire _10163_ ;
wire _2085_ ;
wire _8731_ ;
wire _8311_ ;
wire _11788_ ;
wire _11368_ ;
wire _9936_ ;
wire _9516_ ;
wire _4651_ ;
wire _4231_ ;
wire _5856_ ;
wire _5436_ ;
wire _5016_ ;
wire _1776_ ;
wire _1356_ ;
wire _10639_ ;
wire _10219_ ;
wire _687_ ;
wire _267_ ;
wire _3922_ ;
wire _3502_ ;
wire _6394_ ;
wire _10392_ ;
wire _4707_ ;
wire _7599_ ;
wire _7179_ ;
wire _8960_ ;
wire _8540_ ;
wire _8120_ ;
wire _11597_ ;
wire _11177_ ;
wire _3099_ ;
wire _9745_ ;
wire _9325_ ;
wire _4880_ ;
wire _4460_ ;
wire _4040_ ;
wire _5665_ ;
wire _5245_ ;
wire _1585_ ;
wire _1165_ ;
wire _7811_ ;
wire _10868_ ;
wire _10448_ ;
wire _10028_ ;
wire _496_ ;
wire _3731_ ;
wire _3311_ ;
wire _4936_ ;
wire _4516_ ;
wire _9974_ ;
wire _9554_ ;
wire _9134_ ;
wire _5894_ ;
wire _5474_ ;
wire _5054_ ;
wire _6679_ ;
wire _6259_ ;
wire _1394_ ;
wire _7620_ ;
wire _7200_ ;
wire _10677_ ;
wire _10257_ ;
wire _2599_ ;
wire _2179_ ;
wire _8825_ ;
wire _8405_ ;
wire _3960_ ;
wire _3540_ ;
wire _3120_ ;
wire _4745_ ;
wire _4325_ ;
wire _24_ ;
wire _9783_ ;
wire _9363_ ;
wire _2811_ ;
wire _5283_ ;
wire _6488_ ;
wire _6068_ ;
wire _10486_ ;
wire _10066_ ;
wire _8634_ ;
wire _8214_ ;
wire _9839_ ;
wire _9419_ ;
wire _4974_ ;
wire _4554_ ;
wire _4134_ ;
wire _5759_ ;
wire _5339_ ;
wire _6700_ ;
wire _9592_ ;
wire _9172_ ;
wire _1679_ ;
wire _1259_ ;
wire _7905_ ;
wire _2620_ ;
wire _2200_ ;
wire _5092_ ;
wire _11903_ ;
wire _3825_ ;
wire _3405_ ;
wire _6297_ ;
wire _10295_ ;
wire _8863_ ;
wire _8443_ ;
wire _8023_ ;
wire _9648_ ;
wire _9228_ ;
wire _4783_ ;
wire _4363_ ;
wire _802_ ;
wire _5988_ ;
wire _5568_ ;
wire _5148_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _7714_ ;
wire _399_ ;
wire _11712_ ;
wire _8919_ ;
wire _3634_ ;
wire _3214_ ;
wire _4839_ ;
wire _4419_ ;
wire _8672_ ;
wire _8252_ ;
wire _1700_ ;
wire _9877_ ;
wire _9457_ ;
wire _9037_ ;
wire _4592_ ;
wire _4172_ ;
wire _611_ ;
wire _2905_ ;
wire _5797_ ;
wire _5377_ ;
wire _1297_ ;
wire _7943_ ;
wire _7523_ ;
wire _7103_ ;
wire _11521_ ;
wire _11101_ ;
wire _8728_ ;
wire _8308_ ;
wire _3863_ ;
wire _3443_ ;
wire _3023_ ;
wire _4648_ ;
wire _4228_ ;
wire _8481_ ;
wire _8061_ ;
wire _9686_ ;
wire _9266_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _5186_ ;
wire _3919_ ;
wire _7752_ ;
wire _7332_ ;
wire _10389_ ;
wire _11750_ ;
wire _11330_ ;
wire _8957_ ;
wire _8537_ ;
wire _8117_ ;
wire _3672_ ;
wire _3252_ ;
wire _4877_ ;
wire _4457_ ;
wire _4037_ ;
wire _8290_ ;
wire _6603_ ;
wire _9495_ ;
wire _9075_ ;
wire _10601_ ;
wire _7808_ ;
wire _2943_ ;
wire _2523_ ;
wire _2103_ ;
wire _11806_ ;
wire _3728_ ;
wire _3308_ ;
wire _7981_ ;
wire _7561_ ;
wire _7141_ ;
wire _10198_ ;
wire _8766_ ;
wire _8346_ ;
wire _3481_ ;
wire _3061_ ;
wire _4686_ ;
wire _4266_ ;
wire _705_ ;
wire _6832_ ;
wire _6412_ ;
wire _10830_ ;
wire _10410_ ;
wire _7617_ ;
wire _2752_ ;
wire _2332_ ;
wire _11615_ ;
wire _3957_ ;
wire _3537_ ;
wire _3117_ ;
wire _7790_ ;
wire _7370_ ;
wire _8995_ ;
wire _8575_ ;
wire _8155_ ;
wire _3290_ ;
wire _1603_ ;
wire _4495_ ;
wire _4075_ ;
wire _934_ ;
wire _514_ ;
wire _2808_ ;
wire _6641_ ;
wire _6221_ ;
wire _7846_ ;
wire _7426_ ;
wire _7006_ ;
wire _2981_ ;
wire _2561_ ;
wire _2141_ ;
wire _11844_ ;
wire _11424_ ;
wire _11004_ ;
wire _3766_ ;
wire _3346_ ;
wire _5912_ ;
wire _8384_ ;
wire _1832_ ;
wire _1412_ ;
wire _9589_ ;
wire _9169_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _5089_ ;
wire _6870_ ;
wire _6450_ ;
wire _6030_ ;
wire _7655_ ;
wire _7235_ ;
wire _2790_ ;
wire _2370_ ;
wire _11653_ ;
wire _11233_ ;
wire _3995_ ;
wire _3575_ ;
wire _3155_ ;
wire _9801_ ;
wire _5721_ ;
wire _5301_ ;
wire _8193_ ;
wire _59_ ;
wire _6926_ ;
wire _6506_ ;
wire _1641_ ;
wire _1221_ ;
wire _9398_ ;
wire _10924_ ;
wire _10504_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2846_ ;
wire _2426_ ;
wire _2006_ ;
wire _11709_ ;
wire _7884_ ;
wire _7464_ ;
wire _7044_ ;
wire _11882_ ;
wire _11462_ ;
wire _11042_ ;
wire _8669_ ;
wire _8249_ ;
wire _3384_ ;
wire _9610_ ;
wire _4589_ ;
wire _4169_ ;
wire _5950_ ;
wire _5530_ ;
wire _5110_ ;
wire _608_ ;
wire _6735_ ;
wire _6315_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _10733_ ;
wire _10313_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _11518_ ;
wire _2669__bF$buf0 ;
wire _2669__bF$buf1 ;
wire _2669__bF$buf2 ;
wire _2669__bF$buf3 ;
wire _4801_ ;
wire _7693_ ;
wire _7273_ ;
wire _11691_ ;
wire _11271_ ;
wire _8898_ ;
wire _8478_ ;
wire _8058_ ;
wire _3193_ ;
wire _1926_ ;
wire _1506_ ;
wire _4398_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _6964_ ;
wire _6544_ ;
wire _6124_ ;
wire _10962_ ;
wire _10542_ ;
wire _10122_ ;
wire _590_ ;
wire _170_ ;
wire _7749_ ;
wire _7329_ ;
wire _2884_ ;
wire _2464_ ;
wire _2044_ ;
wire _11747_ ;
wire _11327_ ;
wire _3669_ ;
wire _3249_ ;
wire _4610_ ;
wire _7082_ ;
wire _11080_ ;
wire _5815_ ;
wire _8287_ ;
wire _1735_ ;
wire _1315_ ;
wire breg_16_bF$buf0 ;
wire breg_16_bF$buf1 ;
wire breg_16_bF$buf2 ;
wire breg_16_bF$buf3 ;
wire breg_16_bF$buf4 ;
wire breg_16_bF$buf5 ;
wire _646_ ;
wire _226_ ;
wire _6773_ ;
wire _6353_ ;
wire _10771_ ;
wire _10351_ ;
wire _7978_ ;
wire _7558_ ;
wire _7138_ ;
wire _2693_ ;
wire _2273_ ;
wire _11556_ ;
wire _11136_ ;
wire _3898_ ;
wire _3478_ ;
wire _3058_ ;
wire _9704_ ;
wire _5624_ ;
wire _5204_ ;
wire _8096_ ;
wire _6829_ ;
wire _6409_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _10827_ ;
wire _10407_ ;
wire _875_ ;
wire _455_ ;
wire _2749_ ;
wire _2329_ ;
wire _6582_ ;
wire _6162_ ;
wire _10580_ ;
wire _10160_ ;
wire _7787_ ;
wire _7367_ ;
wire _2082_ ;
wire _11785_ ;
wire _11365_ ;
wire _3287_ ;
wire _9933_ ;
wire _9513_ ;
wire _5853_ ;
wire _5433_ ;
wire _5013_ ;
wire _6638_ ;
wire _6218_ ;
wire _1773_ ;
wire _1353_ ;
wire _10636_ ;
wire _10216_ ;
wire _684_ ;
wire _264_ ;
wire _2978_ ;
wire _2558_ ;
wire _2138_ ;
wire _6391_ ;
wire _4704_ ;
wire _7596_ ;
wire _7176_ ;
wire _11594_ ;
wire _11174_ ;
wire _5909_ ;
wire _3096_ ;
wire _9742_ ;
wire _9322_ ;
wire _1829_ ;
wire _1409_ ;
wire _5662_ ;
wire _5242_ ;
wire _6867_ ;
wire _6447_ ;
wire _6027_ ;
wire _1582_ ;
wire _1162_ ;
wire _10865_ ;
wire _10445_ ;
wire _10025_ ;
wire _493_ ;
wire _2787_ ;
wire _2367_ ;
wire _4933_ ;
wire _4513_ ;
wire _5718_ ;
wire _9971_ ;
wire _9551_ ;
wire _9131_ ;
wire _1638_ ;
wire _1218_ ;
wire _5891_ ;
wire _5471_ ;
wire _5051_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _6676_ ;
wire _6256_ ;
wire _1391_ ;
wire _10674_ ;
wire _10254_ ;
wire _2596_ ;
wire _2176_ ;
wire _8822_ ;
wire _8402_ ;
wire _11879_ ;
wire _11459_ ;
wire _11039_ ;
wire _9607_ ;
wire _4742_ ;
wire _4322_ ;
wire _5947_ ;
wire _5527_ ;
wire _5107_ ;
wire _21_ ;
wire _9780_ ;
wire _9360_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _5280_ ;
wire _778_ ;
wire _358_ ;
wire _6485_ ;
wire _6065_ ;
wire _10483_ ;
wire _10063_ ;
wire _8631_ ;
wire _8211_ ;
wire _11688_ ;
wire _11268_ ;
wire _9836_ ;
wire _9416_ ;
wire _4971_ ;
wire _4551_ ;
wire _4131_ ;
wire _5756_ ;
wire _5336_ ;
wire _1676_ ;
wire _1256_ ;
wire _7902_ ;
wire _10959_ ;
wire _10539_ ;
wire _10119_ ;
wire _587_ ;
wire _167_ ;
wire _11900_ ;
wire _3822_ ;
wire _3402_ ;
wire _6294_ ;
wire _10292_ ;
wire _4607_ ;
wire _7499_ ;
wire _7079_ ;
wire _8860_ ;
wire _8440_ ;
wire _8020_ ;
wire _11497_ ;
wire _11077_ ;
wire _9645_ ;
wire _9225_ ;
wire _4780_ ;
wire _4360_ ;
wire _5985_ ;
wire _5565_ ;
wire _5145_ ;
wire _2519__bF$buf0 ;
wire _2519__bF$buf1 ;
wire _2519__bF$buf2 ;
wire _2519__bF$buf3 ;
wire _1485_ ;
wire _1065_ ;
wire _7711_ ;
wire _10768_ ;
wire _10348_ ;
wire _396_ ;
wire _8916_ ;
wire _3631_ ;
wire _3211_ ;
wire _4836_ ;
wire _4416_ ;
wire _9874_ ;
wire _9454_ ;
wire _9034_ ;
wire _2902_ ;
wire _5794_ ;
wire _5374_ ;
wire _6999_ ;
wire _6579_ ;
wire _6159_ ;
wire _1294_ ;
wire _7940_ ;
wire _7520_ ;
wire _7100_ ;
wire _10997_ ;
wire _10577_ ;
wire _10157_ ;
wire _2499_ ;
wire _2079_ ;
wire _8725_ ;
wire _8305_ ;
wire _3860_ ;
wire _3440_ ;
wire _3020_ ;
wire _4645_ ;
wire _4225_ ;
wire _9683_ ;
wire _9263_ ;
wire _2711_ ;
wire _5183_ ;
wire _3916_ ;
wire _6388_ ;
wire _10386_ ;
wire _8954_ ;
wire _8534_ ;
wire _8114_ ;
wire _9739_ ;
wire _9319_ ;
wire _4874_ ;
wire _4454_ ;
wire _4034_ ;
wire _5659_ ;
wire _5239_ ;
wire _6600_ ;
wire _9492_ ;
wire _9072_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _7805_ ;
wire _2940_ ;
wire _2520_ ;
wire _2100_ ;
wire _11803_ ;
wire _3725_ ;
wire _3305_ ;
wire _6197_ ;
wire _10195_ ;
wire _8763_ ;
wire _8343_ ;
wire _9968_ ;
wire _9548_ ;
wire _9128_ ;
wire _4683_ ;
wire _4263_ ;
wire _702_ ;
wire _5888_ ;
wire _5468_ ;
wire _5048_ ;
wire _5921__bF$buf0 ;
wire _5921__bF$buf1 ;
wire _5921__bF$buf2 ;
wire _5921__bF$buf3 ;
wire _1388_ ;
wire _7614_ ;
wire _299_ ;
wire _11612_ ;
wire _8819_ ;
wire _3954_ ;
wire _3534_ ;
wire _3114_ ;
wire _4739_ ;
wire _4319_ ;
wire _8992_ ;
wire _8572_ ;
wire _8152_ ;
wire areg_18_bF$buf0 ;
wire areg_18_bF$buf1 ;
wire areg_18_bF$buf2 ;
wire areg_18_bF$buf3 ;
wire areg_18_bF$buf4 ;
wire areg_18_bF$buf5 ;
wire _18_ ;
wire _1600_ ;
wire _9777_ ;
wire _9357_ ;
wire _4492_ ;
wire _4072_ ;
wire _931_ ;
wire _511_ ;
wire _2805_ ;
wire _5697_ ;
wire _5277_ ;
wire _1197_ ;
wire _7843_ ;
wire _7423_ ;
wire _7003_ ;
wire _11841_ ;
wire _11421_ ;
wire _11001_ ;
wire _8628_ ;
wire _8208_ ;
wire _3763_ ;
wire _3343_ ;
wire _4968_ ;
wire _4548_ ;
wire _4128_ ;
wire _8381_ ;
wire _9586_ ;
wire _9166_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _5086_ ;
wire _3819_ ;
wire _7652_ ;
wire _7232_ ;
wire _10289_ ;
wire _11650_ ;
wire _11230_ ;
wire _8857_ ;
wire _8437_ ;
wire _8017_ ;
wire _3992_ ;
wire _3572_ ;
wire _3152_ ;
wire _4777_ ;
wire _4357_ ;
wire _8190_ ;
wire _56_ ;
wire _6923_ ;
wire _6503_ ;
wire _9395_ ;
wire _10921_ ;
wire _10501_ ;
wire _7708_ ;
wire _2843_ ;
wire _2423_ ;
wire _2003_ ;
wire _11706_ ;
wire _3628_ ;
wire _3208_ ;
wire _7881_ ;
wire _7461_ ;
wire _7041_ ;
wire _10098_ ;
wire _8666_ ;
wire _8246_ ;
wire _3381_ ;
wire _4586_ ;
wire _4166_ ;
wire _605_ ;
wire _6732_ ;
wire _6312_ ;
wire _10730_ ;
wire _10310_ ;
wire _7937_ ;
wire _7517_ ;
wire _2652_ ;
wire _2232_ ;
wire _11515_ ;
wire _3857_ ;
wire _3437_ ;
wire _3017_ ;
wire _7690_ ;
wire _7270_ ;
wire _8895_ ;
wire _8475_ ;
wire _8055_ ;
wire _3190_ ;
wire _1923_ ;
wire _1503_ ;
wire _4395_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _6961_ ;
wire _6541_ ;
wire _6121_ ;
wire _7746_ ;
wire _7326_ ;
wire _2881_ ;
wire _2461_ ;
wire _2041_ ;
wire _11744_ ;
wire _11324_ ;
wire _3666_ ;
wire _3246_ ;
wire _5812_ ;
wire _8284_ ;
wire _1732_ ;
wire _1312_ ;
wire _9489_ ;
wire _9069_ ;
wire _643_ ;
wire _223_ ;
wire _2937_ ;
wire _2517_ ;
wire _6770_ ;
wire _6350_ ;
wire _7975_ ;
wire _7555_ ;
wire _7135_ ;
wire _2690_ ;
wire _2270_ ;
wire _11553_ ;
wire _11133_ ;
wire _3895_ ;
wire _3475_ ;
wire _3055_ ;
wire _9701_ ;
wire _5621_ ;
wire _5201_ ;
wire _8093_ ;
wire _6826_ ;
wire _6406_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _9298_ ;
wire _10824_ ;
wire _10404_ ;
wire _872_ ;
wire _452_ ;
wire _2746_ ;
wire _2326_ ;
wire _11609_ ;
wire _7784_ ;
wire _7364_ ;
wire _11782_ ;
wire _11362_ ;
wire _8989_ ;
wire _8569_ ;
wire _8149_ ;
wire _3284_ ;
wire _9930_ ;
wire _9510_ ;
wire _4489_ ;
wire _4069_ ;
wire _5850_ ;
wire _5430_ ;
wire _5010_ ;
wire _928_ ;
wire _508_ ;
wire _6635_ ;
wire _6215_ ;
wire _1770_ ;
wire _1350_ ;
wire _10633_ ;
wire _10213_ ;
wire _681_ ;
wire _261_ ;
wire _2975_ ;
wire _2555_ ;
wire _2135_ ;
wire _11838_ ;
wire _11418_ ;
wire _4701_ ;
wire _7593_ ;
wire _7173_ ;
wire _11591_ ;
wire _11171_ ;
wire _5906_ ;
wire _8798_ ;
wire _8378_ ;
wire _3093_ ;
wire _1826_ ;
wire _1406_ ;
wire _4298_ ;
wire _737_ ;
wire _317_ ;
wire _6864_ ;
wire _6444_ ;
wire _6024_ ;
wire _10862_ ;
wire _10442_ ;
wire _10022_ ;
wire _490_ ;
wire _7649_ ;
wire _7229_ ;
wire _2784_ ;
wire _2364_ ;
wire _11647_ ;
wire _11227_ ;
wire _3989_ ;
wire _3569_ ;
wire _3149_ ;
wire _4930_ ;
wire _4510_ ;
wire _5715_ ;
wire _8187_ ;
wire _1635_ ;
wire _1215_ ;
wire _10918_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _6673_ ;
wire _6253_ ;
wire _10671_ ;
wire _10251_ ;
wire _7878_ ;
wire _7458_ ;
wire _7038_ ;
wire _2593_ ;
wire _2173_ ;
wire _11876_ ;
wire _11456_ ;
wire _11036_ ;
wire _3798_ ;
wire _3378_ ;
wire _9604_ ;
wire _5944_ ;
wire _5524_ ;
wire _5104_ ;
wire _6729_ ;
wire _6309_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _10727_ ;
wire _10307_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _6482_ ;
wire _6062_ ;
wire _10480_ ;
wire _10060_ ;
wire _7687_ ;
wire _7267_ ;
wire _11685_ ;
wire _11265_ ;
wire _3187_ ;
wire _9833_ ;
wire _9413_ ;
wire _5753_ ;
wire _5333_ ;
wire _6958_ ;
wire _6538_ ;
wire _6118_ ;
wire _1673_ ;
wire _1253_ ;
wire _10956_ ;
wire _10536_ ;
wire _10116_ ;
wire _584_ ;
wire _164_ ;
wire _2878_ ;
wire _2458_ ;
wire _2038_ ;
wire _6291_ ;
wire _4604_ ;
wire _7496_ ;
wire _7076_ ;
wire _11494_ ;
wire _11074_ ;
wire _5809_ ;
wire _9642_ ;
wire _9222_ ;
wire _1729_ ;
wire _1309_ ;
wire _5982_ ;
wire _5562_ ;
wire _5142_ ;
wire _6767_ ;
wire _6347_ ;
wire _1482_ ;
wire _1062_ ;
wire _10765_ ;
wire _10345_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _8913_ ;
wire _4833_ ;
wire _4413_ ;
wire _5618_ ;
wire _9871_ ;
wire _9451_ ;
wire _9031_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _5791_ ;
wire _5371_ ;
wire _869_ ;
wire _449_ ;
wire _6996_ ;
wire _6576_ ;
wire _6156_ ;
wire _1291_ ;
wire _10994_ ;
wire _10574_ ;
wire _10154_ ;
wire _2496_ ;
wire _2076_ ;
wire _8722_ ;
wire _8302_ ;
wire _11779_ ;
wire _11359_ ;
wire _9927_ ;
wire _9507_ ;
wire _4642_ ;
wire _4222_ ;
wire _5847_ ;
wire _5427_ ;
wire _5007_ ;
wire _9680_ ;
wire _9260_ ;
wire _1767_ ;
wire _1347_ ;
wire _5180_ ;
wire _678_ ;
wire _258_ ;
wire _3913_ ;
wire _6385_ ;
wire _10383_ ;
wire _8951_ ;
wire _8531_ ;
wire _8111_ ;
wire _11588_ ;
wire _11168_ ;
wire _9736_ ;
wire _9316_ ;
wire _4871_ ;
wire _4451_ ;
wire _4031_ ;
wire _5656_ ;
wire _5236_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _7802_ ;
wire _10859_ ;
wire _10439_ ;
wire _10019_ ;
wire _487_ ;
wire _11800_ ;
wire _3722_ ;
wire _3302_ ;
wire _6194_ ;
wire breg_11_bF$buf0 ;
wire breg_11_bF$buf1 ;
wire breg_11_bF$buf2 ;
wire _10192_ ;
wire breg_11_bF$buf3 ;
wire breg_11_bF$buf4 ;
wire _4927_ ;
wire _4507_ ;
wire _7399_ ;
wire _8760_ ;
wire _8340_ ;
wire _11397_ ;
wire _9965_ ;
wire _9545_ ;
wire _9125_ ;
wire _4680_ ;
wire _4260_ ;
wire _5885_ ;
wire _5465_ ;
wire _5045_ ;
wire _1385_ ;
wire _7611_ ;
wire _10668_ ;
wire _10248_ ;
wire _296_ ;
wire _8816_ ;
wire _3951_ ;
wire _3531_ ;
wire _3111_ ;
wire _4736_ ;
wire _4316_ ;
wire _15_ ;
wire _9774_ ;
wire _9354_ ;
wire _2802_ ;
wire _5694_ ;
wire _5274_ ;
wire _6899_ ;
wire _6479_ ;
wire _6059_ ;
wire _1194_ ;
wire _7840_ ;
wire _7420_ ;
wire _7000_ ;
wire _10897_ ;
wire _10477_ ;
wire _10057_ ;
wire _2399_ ;
wire _8625_ ;
wire _8205_ ;
wire _3760_ ;
wire _3340_ ;
wire _4965_ ;
wire _4545_ ;
wire _4125_ ;
wire _9583_ ;
wire _9163_ ;
wire _2611_ ;
wire _5083_ ;
wire _3816_ ;
wire _6288_ ;
wire _10286_ ;
wire _8854_ ;
wire _8434_ ;
wire _8014_ ;
wire _9639_ ;
wire _9219_ ;
wire _4774_ ;
wire _4354_ ;
wire _5979_ ;
wire _5559_ ;
wire _5139_ ;
wire _53_ ;
wire _6920_ ;
wire _6500_ ;
wire _9392_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _7705_ ;
wire _2840_ ;
wire _2420_ ;
wire _2000_ ;
wire _11703_ ;
wire _3625_ ;
wire _3205_ ;
wire _6097_ ;
wire _10095_ ;
wire _8663_ ;
wire _8243_ ;
wire _9868_ ;
wire _9448_ ;
wire _9028_ ;
wire _4583_ ;
wire _4163_ ;
wire areg_29_bF$buf0 ;
wire areg_29_bF$buf1 ;
wire areg_29_bF$buf2 ;
wire areg_29_bF$buf3 ;
wire areg_29_bF$buf4 ;
wire areg_29_bF$buf5 ;
wire _602_ ;
wire _5788_ ;
wire _5368_ ;
wire [31:0] breg ;
wire _1288_ ;
wire _7934_ ;
wire _7514_ ;
wire _199_ ;
wire _11512_ ;
wire _8719_ ;
wire _3854_ ;
wire _3434_ ;
wire _3014_ ;
wire _4639_ ;
wire _4219_ ;
wire _8892_ ;
wire _8472_ ;
wire _8052_ ;
wire _1920_ ;
wire _1500_ ;
wire _9677_ ;
wire _9257_ ;
wire _4392_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _6300__bF$buf0 ;
wire _6300__bF$buf1 ;
wire _6300__bF$buf2 ;
wire _5597_ ;
wire _6300__bF$buf3 ;
wire _5177_ ;
wire _91_ ;
wire _1097_ ;
wire _7743_ ;
wire _7323_ ;
wire _11741_ ;
wire _11321_ ;
wire _8948_ ;
wire _8528_ ;
wire _8108_ ;
wire _3663_ ;
wire _3243_ ;
wire _4868_ ;
wire _4448_ ;
wire _4028_ ;
wire _8281_ ;
wire _9486_ ;
wire _9066_ ;
wire _640_ ;
wire _220_ ;
wire _2934_ ;
wire _2514_ ;
wire _3719_ ;
wire _7972_ ;
wire _7552_ ;
wire _7132_ ;
wire _10189_ ;
wire _11550_ ;
wire _11130_ ;
wire _8757_ ;
wire _8337_ ;
wire _3892_ ;
wire _3472_ ;
wire _3052_ ;
wire _4677_ ;
wire _4257_ ;
wire _8090_ ;
wire _6823_ ;
wire _6403_ ;
wire _9295_ ;
wire _10821_ ;
wire _10401_ ;
wire _7608_ ;
wire _2743_ ;
wire _2323_ ;
wire _11606_ ;
wire _3948_ ;
wire _3528_ ;
wire _3108_ ;
wire _9_ ;
wire _7781_ ;
wire _7361_ ;
wire _8986_ ;
wire _8566_ ;
wire _8146_ ;
wire _3281_ ;
wire _4486_ ;
wire _4066_ ;
wire _925_ ;
wire _505_ ;
wire _6632_ ;
wire _6212_ ;
wire _10630_ ;
wire _10210_ ;
wire _7837_ ;
wire _7417_ ;
wire _2972_ ;
wire _2552_ ;
wire _2132_ ;
wire _11835_ ;
wire _11415_ ;
wire _3757_ ;
wire _3337_ ;
wire _7590_ ;
wire _7170_ ;
wire _5903_ ;
wire _8795_ ;
wire _8375_ ;
wire _3090_ ;
wire _1823_ ;
wire _1403_ ;
wire _4295_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _6861_ ;
wire _6441_ ;
wire _6021_ ;
wire _7646_ ;
wire _7226_ ;
wire _2781_ ;
wire _2361_ ;
wire _11644_ ;
wire _11224_ ;
wire _3986_ ;
wire _3566_ ;
wire _3146_ ;
wire _5712_ ;
wire _8184_ ;
wire _6917_ ;
wire _1632_ ;
wire _1212_ ;
wire _9389_ ;
wire _10915_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2837_ ;
wire _2417_ ;
wire _6670_ ;
wire _6250_ ;
wire _7875_ ;
wire _7455_ ;
wire _7035_ ;
wire _2590_ ;
wire _2170_ ;
wire _11873_ ;
wire _11453_ ;
wire _11033_ ;
wire _3795_ ;
wire _3375_ ;
wire _9601_ ;
wire _5941_ ;
wire _5521_ ;
wire _5101_ ;
wire _6726_ ;
wire _6306_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _9198_ ;
wire _10724_ ;
wire _10304_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire areg_13_bF$buf0 ;
wire _11509_ ;
wire areg_13_bF$buf1 ;
wire areg_13_bF$buf2 ;
wire areg_13_bF$buf3 ;
wire areg_13_bF$buf4 ;
wire _7684_ ;
wire _7264_ ;
wire _11682_ ;
wire _11262_ ;
wire _8889_ ;
wire _8469_ ;
wire _8049_ ;
wire _3184_ ;
wire _9830_ ;
wire _9410_ ;
wire _1917_ ;
wire _4389_ ;
wire _5750_ ;
wire _5330_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _6955_ ;
wire _2825__bF$buf0 ;
wire _6535_ ;
wire _2825__bF$buf1 ;
wire _6115_ ;
wire _2825__bF$buf2 ;
wire _2825__bF$buf3 ;
wire _2825__bF$buf4 ;
wire _1670_ ;
wire _1250_ ;
wire _10953_ ;
wire _10533_ ;
wire _10113_ ;
wire _581_ ;
wire _161_ ;
wire _2875_ ;
wire _2455_ ;
wire _2035_ ;
wire _11738_ ;
wire _11318_ ;
wire _4601_ ;
wire _7493_ ;
wire _7073_ ;
wire _11491_ ;
wire _11071_ ;
wire _5806_ ;
wire _8698_ ;
wire _8278_ ;
wire _1726_ ;
wire _1306_ ;
wire _4198_ ;
wire _637_ ;
wire _217_ ;
wire _6764_ ;
wire _6344_ ;
wire _10762_ ;
wire _10342_ ;
wire _390_ ;
wire _7969_ ;
wire _7549_ ;
wire _7129_ ;
wire _2684_ ;
wire _2264_ ;
wire _8910_ ;
wire _11547_ ;
wire _11127_ ;
wire _3889_ ;
wire _3469_ ;
wire _3049_ ;
wire _4830_ ;
wire _4410_ ;
wire _5615_ ;
wire _8087_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _10818_ ;
wire _866_ ;
wire _446_ ;
wire _6993_ ;
wire _6573_ ;
wire _6153_ ;
wire _10991_ ;
wire _10571_ ;
wire _10151_ ;
wire _7778_ ;
wire _7358_ ;
wire _2493_ ;
wire _2073_ ;
wire _11776_ ;
wire _11356_ ;
wire _3698_ ;
wire _3278_ ;
wire _9924_ ;
wire _9504_ ;
wire _5844_ ;
wire _5424_ ;
wire _5004_ ;
wire _3961__bF$buf0 ;
wire _3961__bF$buf1 ;
wire _3961__bF$buf2 ;
wire _3961__bF$buf3 ;
wire _3961__bF$buf4 ;
wire _6629_ ;
wire _6209_ ;
wire _1764_ ;
wire _1344_ ;
wire _10627_ ;
wire _10207_ ;
wire _675_ ;
wire _255_ ;
wire _2969_ ;
wire _2549_ ;
wire _2129_ ;
wire _3910_ ;
wire _6382_ ;
wire _10380_ ;
wire _7587_ ;
wire _7167_ ;
wire _11585_ ;
wire _11165_ ;
wire _3087_ ;
wire _3646__bF$buf0 ;
wire _3646__bF$buf1 ;
wire _9733_ ;
wire _3646__bF$buf2 ;
wire _9313_ ;
wire _3646__bF$buf3 ;
wire _5653_ ;
wire _5233_ ;
wire _6858_ ;
wire _6438_ ;
wire _6018_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _10856_ ;
wire _10436_ ;
wire _10016_ ;
wire _484_ ;
wire _2778_ ;
wire _2358_ ;
wire _6191_ ;
wire _4924_ ;
wire _4504_ ;
wire _7396_ ;
wire _11394_ ;
wire _5709_ ;
wire _9962_ ;
wire _9542_ ;
wire _9122_ ;
wire _1629_ ;
wire _1209_ ;
wire _5882_ ;
wire _5462_ ;
wire _5042_ ;
wire _6667_ ;
wire _6247_ ;
wire _1382_ ;
wire _10665_ ;
wire _10245_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _8813_ ;
wire _4733_ ;
wire _4313_ ;
wire _5938_ ;
wire _5518_ ;
wire _12_ ;
wire _9771_ ;
wire _9351_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _5691_ ;
wire _5271_ ;
wire _769_ ;
wire _349_ ;
wire _6896_ ;
wire _6476_ ;
wire _6056_ ;
wire _1191_ ;
wire _10894_ ;
wire _10474_ ;
wire _10054_ ;
wire _2396_ ;
wire _8622_ ;
wire _8202_ ;
wire _11679_ ;
wire _11259_ ;
wire _9827_ ;
wire _9407_ ;
wire _4962_ ;
wire _4542_ ;
wire _4122_ ;
wire _5747_ ;
wire _5327_ ;
wire _9580_ ;
wire _9160_ ;
wire _1667_ ;
wire _1247_ ;
wire _5080_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _3813_ ;
wire _6285_ ;
wire _10283_ ;
wire _8851_ ;
wire _8431_ ;
wire _8011_ ;
wire _11488_ ;
wire _11068_ ;
wire _9636_ ;
wire _9216_ ;
wire _4771_ ;
wire _4351_ ;
wire _5976_ ;
wire _5556_ ;
wire _5136_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _7702_ ;
wire _10759_ ;
wire _10339_ ;
wire _387_ ;
wire _11700_ ;
wire _8907_ ;
wire _3622_ ;
wire _3202_ ;
wire _6094_ ;
wire breg_9_bF$buf0 ;
wire _10092_ ;
wire breg_9_bF$buf1 ;
wire breg_9_bF$buf2 ;
wire breg_9_bF$buf3 ;
wire _4827_ ;
wire breg_9_bF$buf4 ;
wire _4407_ ;
wire breg_9_bF$buf5 ;
wire _7299_ ;
wire _8660_ ;
wire _8240_ ;
wire _11297_ ;
wire _9865_ ;
wire _9445_ ;
wire _9025_ ;
wire _4580_ ;
wire _4160_ ;
wire _5785_ ;
wire _5365_ ;
wire _1285_ ;
wire _7931_ ;
wire _7511_ ;
wire _10988_ ;
wire _10568_ ;
wire _10148_ ;
wire _196_ ;
wire _8716_ ;
wire _3851_ ;
wire _3431_ ;
wire _3011_ ;
wire _4636_ ;
wire _4216_ ;
wire _9674_ ;
wire _9254_ ;
wire _2702_ ;
wire _5594_ ;
wire _5174_ ;
wire _3907_ ;
wire _6799_ ;
wire _6379_ ;
wire _1094_ ;
wire _7740_ ;
wire _7320_ ;
wire _10797_ ;
wire _10377_ ;
wire _2299_ ;
wire _8945_ ;
wire _8525_ ;
wire _8105_ ;
wire _3660_ ;
wire _3240_ ;
wire _4865_ ;
wire _4445_ ;
wire _4025_ ;
wire _9483_ ;
wire _9063_ ;
wire _2931_ ;
wire _2511_ ;
wire _3716_ ;
wire _6188_ ;
wire _10186_ ;
wire _8754_ ;
wire _8334_ ;
wire _9959_ ;
wire _9539_ ;
wire _9119_ ;
wire _4674_ ;
wire _4254_ ;
wire _5879_ ;
wire _5459_ ;
wire _5039_ ;
wire _6820_ ;
wire _6400_ ;
wire _9292_ ;
wire _1799_ ;
wire _1379_ ;
wire _7605_ ;
wire _2740_ ;
wire _2320_ ;
wire _11603_ ;
wire _3945_ ;
wire _3525_ ;
wire _3105_ ;
wire _6_ ;
wire _8983_ ;
wire _8563_ ;
wire _8143_ ;
wire _9768_ ;
wire _9348_ ;
wire _4483_ ;
wire _4063_ ;
wire _922_ ;
wire _502_ ;
wire _5688_ ;
wire _5268_ ;
wire [31:0] areg ;
wire _1188_ ;
wire _7834_ ;
wire _7414_ ;
wire _11832_ ;
wire _11412_ ;
wire _8619_ ;
wire _3754_ ;
wire _3334_ ;
wire _4959_ ;
wire _4539_ ;
wire _4119_ ;
wire _5900_ ;
wire _8792_ ;
wire _8372_ ;
wire _1820_ ;
wire _1400_ ;
wire _9997_ ;
wire _9577_ ;
wire _9157_ ;
wire _4292_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _5497_ ;
wire _5077_ ;
wire _7643_ ;
wire _7223_ ;
wire _11641_ ;
wire _11221_ ;
wire _8848_ ;
wire _8428_ ;
wire _8008_ ;
wire _3983_ ;
wire _3563_ ;
wire _3143_ ;
wire _4768_ ;
wire _4348_ ;
wire _8181_ ;
wire _47_ ;
wire _6914_ ;
wire _9386_ ;
wire _10912_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2834_ ;
wire _2414_ ;
wire _3619_ ;
wire _7872_ ;
wire _7452_ ;
wire _7032_ ;
wire _10089_ ;
wire _11870_ ;
wire _11450_ ;
wire _11030_ ;
wire _8657_ ;
wire _8237_ ;
wire _3792_ ;
wire _3372_ ;
wire _4997_ ;
wire _4577_ ;
wire _4157_ ;
wire _6723_ ;
wire _6303_ ;
wire _9195_ ;
wire _10721_ ;
wire _10301_ ;
wire _7928_ ;
wire _7508_ ;
wire _2643_ ;
wire _2223_ ;
wire _11506_ ;
wire _3848_ ;
wire _3428_ ;
wire _3008_ ;
wire _7681_ ;
wire _7261_ ;
wire _8886_ ;
wire _8466_ ;
wire _8046_ ;
wire _3181_ ;
wire _1914_ ;
wire _4386_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _6952_ ;
wire _6532_ ;
wire _6112_ ;
wire _10950_ ;
wire _10530_ ;
wire _10110_ ;
wire _7737_ ;
wire _7317_ ;
wire _2872_ ;
wire _2452_ ;
wire _2032_ ;
wire _11735_ ;
wire _11315_ ;
wire _3657_ ;
wire _3237_ ;
wire _7490_ ;
wire _7070_ ;
wire _5803_ ;
wire _8695_ ;
wire _8275_ ;
wire _1723_ ;
wire _1303_ ;
wire _4195_ ;
wire _634_ ;
wire _214_ ;
wire _2928_ ;
wire _2508_ ;
wire _6761_ ;
wire _6341_ ;
wire _7966_ ;
wire _7546_ ;
wire _7126_ ;
wire _2681_ ;
wire _2261_ ;
wire _11544_ ;
wire _11124_ ;
wire _3886_ ;
wire _3466_ ;
wire _3046_ ;
wire _5612_ ;
wire _8084_ ;
wire _6817_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _9289_ ;
wire _10815_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _6990_ ;
wire _6570_ ;
wire _6150_ ;
wire _7775_ ;
wire _7355_ ;
wire areg_24_bF$buf0 ;
wire areg_24_bF$buf1 ;
wire areg_24_bF$buf2 ;
wire _2490_ ;
wire areg_24_bF$buf3 ;
wire _2070_ ;
wire areg_24_bF$buf4 ;
wire _11773_ ;
wire _11353_ ;
wire _3695_ ;
wire _3275_ ;
wire _9921_ ;
wire _9501_ ;
wire _5841_ ;
wire _5421_ ;
wire _5001_ ;
wire _919_ ;
wire _6626_ ;
wire _6206_ ;
wire _1761_ ;
wire _1341_ ;
wire _9098_ ;
wire _10624_ ;
wire _10204_ ;
wire _672_ ;
wire _252_ ;
wire _2966_ ;
wire _2546_ ;
wire _2126_ ;
wire _11829_ ;
wire _11409_ ;
wire _7584_ ;
wire _7164_ ;
wire _11582_ ;
wire _11162_ ;
wire _8789_ ;
wire _8369_ ;
wire _3084_ ;
wire _9730_ ;
wire _9310_ ;
wire _1817_ ;
wire _4289_ ;
wire _5650_ ;
wire _5230_ ;
wire _728_ ;
wire _308_ ;
wire _6855_ ;
wire _6435_ ;
wire _6015_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _10853_ ;
wire _10433_ ;
wire _10013_ ;
wire _481_ ;
wire _2775_ ;
wire _2355_ ;
wire _11638_ ;
wire _11218_ ;
wire _4921_ ;
wire _4501_ ;
wire _7393_ ;
wire _11391_ ;
wire _5706_ ;
wire _8598_ ;
wire _8178_ ;
wire _1626_ ;
wire _1206_ ;
wire _4098_ ;
wire _10909_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _6815__bF$buf0 ;
wire _6815__bF$buf1 ;
wire _6815__bF$buf2 ;
wire _6815__bF$buf3 ;
wire _6815__bF$buf4 ;
wire _6664_ ;
wire _6244_ ;
wire _10662_ ;
wire _10242_ ;
wire _290_ ;
wire _7869_ ;
wire _7449_ ;
wire _7029_ ;
wire _2584_ ;
wire _2164_ ;
wire _8810_ ;
wire _11867_ ;
wire _11447_ ;
wire _11027_ ;
wire _3789_ ;
wire _3369_ ;
wire _4730_ ;
wire _4310_ ;
wire _5935_ ;
wire _5515_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _10718_ ;
wire _766_ ;
wire _346_ ;
wire _6893_ ;
wire _6473_ ;
wire _6053_ ;
wire _10891_ ;
wire _10471_ ;
wire _10051_ ;
wire _7678_ ;
wire _7258_ ;
wire _2393_ ;
wire _11676_ ;
wire _11256_ ;
wire _3598_ ;
wire _3178_ ;
wire _9824_ ;
wire _9404_ ;
wire areg_6_bF$buf0 ;
wire areg_6_bF$buf1 ;
wire areg_6_bF$buf2 ;
wire areg_6_bF$buf3 ;
wire areg_6_bF$buf4 ;
wire _5744_ ;
wire _5324_ ;
wire _6949_ ;
wire _6529_ ;
wire _6109_ ;
wire _1664_ ;
wire _1244_ ;
wire _10947_ ;
wire _10527_ ;
wire _10107_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2869_ ;
wire _2449_ ;
wire _2029_ ;
wire _3810_ ;
wire _6282_ ;
wire _10280_ ;
wire _7487_ ;
wire _7067_ ;
wire _11485_ ;
wire _11065_ ;
wire _9633_ ;
wire _9213_ ;
wire _5973_ ;
wire _5553_ ;
wire _5133_ ;
wire _6758_ ;
wire _6338_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _10756_ ;
wire _10336_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _8904_ ;
wire _6091_ ;
wire _4824_ ;
wire _4404_ ;
wire _7296_ ;
wire _11294_ ;
wire _5609_ ;
wire _9862_ ;
wire _9442_ ;
wire _9022_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _5782_ ;
wire _5362_ ;
wire _6987_ ;
wire _6567_ ;
wire _6147_ ;
wire _1282_ ;
wire _10985_ ;
wire _10565_ ;
wire _10145_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _8713_ ;
wire _9918_ ;
wire _4633_ ;
wire _4213_ ;
wire _5838_ ;
wire _5418_ ;
wire _9671_ ;
wire _9251_ ;
wire _1758_ ;
wire _1338_ ;
wire _5591_ ;
wire _5171_ ;
wire _669_ ;
wire _249_ ;
wire _3904_ ;
wire _6796_ ;
wire _6376_ ;
wire _1091_ ;
wire _10794_ ;
wire _10374_ ;
wire _2296_ ;
wire _8942_ ;
wire _8522_ ;
wire _8102_ ;
wire _11579_ ;
wire _11159_ ;
wire _9727_ ;
wire _9307_ ;
wire _4862_ ;
wire _4442_ ;
wire _4022_ ;
wire _5647_ ;
wire _5227_ ;
wire _9480_ ;
wire _9060_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _3713_ ;
wire _6185_ ;
wire _10183_ ;
wire _4918_ ;
wire _8751_ ;
wire _8331_ ;
wire _11388_ ;
wire _9956_ ;
wire _9536_ ;
wire _9116_ ;
wire _4671_ ;
wire _4251_ ;
wire _5876_ ;
wire _5456_ ;
wire _5036_ ;
wire _1796_ ;
wire _1376_ ;
wire _7602_ ;
wire _10659_ ;
wire _10239_ ;
wire _287_ ;
wire _11600_ ;
wire _8807_ ;
wire _3942_ ;
wire _3522_ ;
wire _3102_ ;
wire _3_ ;
wire _4727_ ;
wire _4307_ ;
wire _7199_ ;
wire _8980_ ;
wire _8560_ ;
wire _8140_ ;
wire _11197_ ;
wire _9765_ ;
wire _9345_ ;
wire _4480_ ;
wire _4060_ ;
wire _5685_ ;
wire _5265_ ;
wire _1185_ ;
wire _7831_ ;
wire _7411_ ;
wire _10888_ ;
wire _10468_ ;
wire _10048_ ;
wire _8616_ ;
wire _3751_ ;
wire _3331_ ;
wire _4956_ ;
wire _4536_ ;
wire _4116_ ;
wire _9994_ ;
wire _9574_ ;
wire _9154_ ;
wire _2602_ ;
wire _5494_ ;
wire _5074_ ;
wire _3807_ ;
wire _6699_ ;
wire _6279_ ;
wire _7640_ ;
wire _7220_ ;
wire _10697_ ;
wire _10277_ ;
wire _2199_ ;
wire _8845_ ;
wire _8425_ ;
wire _8005_ ;
wire _3980_ ;
wire _3560_ ;
wire _3140_ ;
wire _4765_ ;
wire _4345_ ;
wire _44_ ;
wire _6911_ ;
wire _9383_ ;
wire _2831_ ;
wire _2411_ ;
wire _3616_ ;
wire _6088_ ;
wire _10086_ ;
wire _8654_ ;
wire _8234_ ;
wire _9859_ ;
wire _9439_ ;
wire _9019_ ;
wire _4994_ ;
wire _4574_ ;
wire _4154_ ;
wire _5779_ ;
wire _5359_ ;
wire _6720_ ;
wire _6300_ ;
wire _9192_ ;
wire _1699_ ;
wire _1279_ ;
wire _7925_ ;
wire _7505_ ;
wire _2640_ ;
wire _2220_ ;
wire _11503_ ;
wire _3845_ ;
wire _3425_ ;
wire _3005_ ;
wire _8883_ ;
wire _8463_ ;
wire _8043_ ;
wire _1911_ ;
wire _9668_ ;
wire _9248_ ;
wire _4383_ ;
wire _822_ ;
wire _402_ ;
wire _5588_ ;
wire _5168_ ;
wire _82_ ;
wire _1088_ ;
wire _7734_ ;
wire _7314_ ;
wire _11732_ ;
wire _11312_ ;
wire _8939_ ;
wire _8519_ ;
wire _3654_ ;
wire _3234_ ;
wire _4859_ ;
wire _4439_ ;
wire _4019_ ;
wire _5800_ ;
wire _8692_ ;
wire _8272_ ;
wire _1720_ ;
wire _1300_ ;
wire _9897_ ;
wire _9477_ ;
wire _9057_ ;
wire _4192_ ;
wire _631_ ;
wire _211_ ;
wire _2925_ ;
wire _2505_ ;
wire _5397_ ;
wire _7963_ ;
wire _7543_ ;
wire _7123_ ;
wire breg_26_bF$buf0 ;
wire breg_26_bF$buf1 ;
wire breg_26_bF$buf2 ;
wire breg_26_bF$buf3 ;
wire _4541__bF$buf0 ;
wire breg_26_bF$buf4 ;
wire _4541__bF$buf1 ;
wire _4541__bF$buf2 ;
wire _4541__bF$buf3 ;
wire _4541__bF$buf4 ;
wire _11541_ ;
wire _11121_ ;
wire _8748_ ;
wire _8328_ ;
wire _3883_ ;
wire _3463_ ;
wire _3043_ ;
wire _4668_ ;
wire _4248_ ;
wire _8081_ ;
wire _6814_ ;
wire _9286_ ;
wire breg_4_bF$buf0 ;
wire breg_4_bF$buf1 ;
wire _10812_ ;
wire breg_4_bF$buf2 ;
wire breg_4_bF$buf3 ;
wire breg_4_bF$buf4 ;
wire breg_4_bF$buf5 ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _3939_ ;
wire _3519_ ;
wire _7772_ ;
wire _7352_ ;
wire _11770_ ;
wire _11350_ ;
wire _8977_ ;
wire _8557_ ;
wire _8137_ ;
wire _3692_ ;
wire _3272_ ;
wire _4897_ ;
wire _4477_ ;
wire _4057_ ;
wire _916_ ;
wire _6623_ ;
wire _6203_ ;
wire _9095_ ;
wire _10621_ ;
wire _10201_ ;
wire _7828_ ;
wire _7408_ ;
wire _2963_ ;
wire _2543_ ;
wire _2123_ ;
wire _11826_ ;
wire _11406_ ;
wire _3748_ ;
wire _3328_ ;
wire _7581_ ;
wire _7161_ ;
wire _8786_ ;
wire _8366_ ;
wire _3081_ ;
wire _1814_ ;
wire _4286_ ;
wire _725_ ;
wire _305_ ;
wire _6852_ ;
wire _6432_ ;
wire _6012_ ;
wire _10850_ ;
wire _10430_ ;
wire _10010_ ;
wire _7637_ ;
wire _7217_ ;
wire _2772_ ;
wire _2352_ ;
wire _11635_ ;
wire _11215_ ;
wire _3977_ ;
wire _3557_ ;
wire _3137_ ;
wire _7390_ ;
wire _5703_ ;
wire _8595_ ;
wire _8175_ ;
wire _6908_ ;
wire _1623_ ;
wire _1203_ ;
wire _4095_ ;
wire _10906_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2828_ ;
wire _2408_ ;
wire _6661_ ;
wire _6241_ ;
wire _7866_ ;
wire _7446_ ;
wire _7026_ ;
wire _2581_ ;
wire _2161_ ;
wire _11864_ ;
wire _11444_ ;
wire _11024_ ;
wire _3786_ ;
wire _3366_ ;
wire _5932_ ;
wire _5512_ ;
wire _6717_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _9189_ ;
wire _10715_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _6890_ ;
wire _6470_ ;
wire _6050_ ;
wire _7675_ ;
wire _7255_ ;
wire _2390_ ;
wire _11673_ ;
wire _11253_ ;
wire _3595_ ;
wire _3175_ ;
wire _9821_ ;
wire _9401_ ;
wire _1908_ ;
wire _5741_ ;
wire _5321_ ;
wire _819_ ;
wire _79_ ;
wire _6946_ ;
wire _6526_ ;
wire _6106_ ;
wire _1661_ ;
wire _1241_ ;
wire _10944_ ;
wire _10524_ ;
wire _10104_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2866_ ;
wire _2446_ ;
wire _2026_ ;
wire _11729_ ;
wire _11309_ ;
wire _7484_ ;
wire _7064_ ;
wire _11482_ ;
wire _11062_ ;
wire _8689_ ;
wire _8269_ ;
wire _9630_ ;
wire _9210_ ;
wire _1717_ ;
wire _4189_ ;
wire _5970_ ;
wire _5550_ ;
wire _5130_ ;
wire _628_ ;
wire _208_ ;
wire _6755_ ;
wire _6335_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _10753_ ;
wire _10333_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _8901_ ;
wire _11538_ ;
wire _11118_ ;
wire _4821_ ;
wire _4401_ ;
wire _7293_ ;
wire _11291_ ;
wire _5606_ ;
wire _8498_ ;
wire _8078_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _10809_ ;
wire _857_ ;
wire _437_ ;
wire _6984_ ;
wire _6564_ ;
wire _6144_ ;
wire _10982_ ;
wire _10562_ ;
wire _10142_ ;
wire _190_ ;
wire _7769_ ;
wire _7349_ ;
wire _2484_ ;
wire _2064_ ;
wire _8710_ ;
wire _11767_ ;
wire _11347_ ;
wire _3689_ ;
wire _3269_ ;
wire _9915_ ;
wire _4630_ ;
wire _4210_ ;
wire _5835_ ;
wire _5415_ ;
wire _1755_ ;
wire _1335_ ;
wire _10618_ ;
wire _666_ ;
wire _246_ ;
wire _3901_ ;
wire _6793_ ;
wire _6373_ ;
wire _10791_ ;
wire _10371_ ;
wire _7998_ ;
wire _7578_ ;
wire _7158_ ;
wire _2293_ ;
wire _11576_ ;
wire _11156_ ;
wire _3498_ ;
wire _3078_ ;
wire _9724_ ;
wire _9304_ ;
wire _5644_ ;
wire _5224_ ;
wire _6849_ ;
wire _6429_ ;
wire _6009_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _10847_ ;
wire _10427_ ;
wire _10007_ ;
wire _895_ ;
wire _475_ ;
wire _2769_ ;
wire _2349_ ;
wire _3710_ ;
wire _6182_ ;
wire _10180_ ;
wire _4915_ ;
wire _7387_ ;
wire _11385_ ;
wire _9953_ ;
wire _9533_ ;
wire _9113_ ;
wire _5873_ ;
wire _5453_ ;
wire _5033_ ;
wire _6658_ ;
wire _6238_ ;
wire _1793_ ;
wire _1373_ ;
wire _10656_ ;
wire _10236_ ;
wire _284_ ;
wire _2998_ ;
wire _2578_ ;
wire _2158_ ;
wire _8804_ ;
wire [63:0] _0_ ;
wire _4724_ ;
wire _4304_ ;
wire _7196_ ;
wire _11194_ ;
wire _5929_ ;
wire _5509_ ;
wire _9762_ ;
wire _9342_ ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _5682_ ;
wire _5262_ ;
wire _6887_ ;
wire _6467_ ;
wire _6047_ ;
wire _1182_ ;
wire _10885_ ;
wire _10465_ ;
wire _10045_ ;
wire _2387_ ;
wire _8613_ ;
wire _9818_ ;
wire _4953_ ;
wire _4533_ ;
wire _4113_ ;
wire _5738_ ;
wire _5318_ ;
wire _9991_ ;
wire _9571_ ;
wire _9151_ ;
wire _1658_ ;
wire _1238_ ;
wire _5491_ ;
wire _5071_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _3804_ ;
wire _6696_ ;
wire _6276_ ;
wire _10694_ ;
wire _10274_ ;
wire _2196_ ;
wire _8842_ ;
wire _8422_ ;
wire _8002_ ;
wire _11899_ ;
wire _11479_ ;
wire _11059_ ;
wire _9627_ ;
wire _9207_ ;
wire _4762_ ;
wire _4342_ ;
wire _5967_ ;
wire _5547_ ;
wire _5127_ ;
wire _41_ ;
wire _9380_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _3613_ ;
wire _6085_ ;
wire _10083_ ;
wire _4818_ ;
wire _8651_ ;
wire _8231_ ;
wire _11288_ ;
wire _9856_ ;
wire _9436_ ;
wire _9016_ ;
wire _4991_ ;
wire _4571_ ;
wire _4151_ ;
wire _5776_ ;
wire _5356_ ;
wire _1696_ ;
wire _1276_ ;
wire _7922_ ;
wire _7502_ ;
wire _10979_ ;
wire _10559_ ;
wire _10139_ ;
wire _187_ ;
wire _11500_ ;
wire _8707_ ;
wire _3842_ ;
wire _3422_ ;
wire _3002_ ;
wire _4627_ ;
wire _4207_ ;
wire _7099_ ;
wire _8880_ ;
wire _8460_ ;
wire _8040_ ;
wire _11097_ ;
wire _9665_ ;
wire _9245_ ;
wire _4380_ ;
wire _5585_ ;
wire _5165_ ;
wire _1085_ ;
wire _7731_ ;
wire _7311_ ;
wire areg_1_bF$buf0 ;
wire areg_1_bF$buf1 ;
wire areg_1_bF$buf2 ;
wire areg_1_bF$buf3 ;
wire areg_1_bF$buf4 ;
wire _10788_ ;
wire _10368_ ;
wire _8936_ ;
wire _8516_ ;
wire _3651_ ;
wire _3231_ ;
wire _4856_ ;
wire _4436_ ;
wire _4016_ ;
wire _9894_ ;
wire _9474_ ;
wire _9054_ ;
wire _2922_ ;
wire _2502_ ;
wire _5394_ ;
wire _3707_ ;
wire _6599_ ;
wire _6179_ ;
wire _7960_ ;
wire _7540_ ;
wire _7120_ ;
wire _10597_ ;
wire _10177_ ;
wire _2099_ ;
wire _8745_ ;
wire _8325_ ;
wire _3880_ ;
wire _3460_ ;
wire _3040_ ;
wire _4665_ ;
wire _4245_ ;
wire _6811_ ;
wire _9283_ ;
wire _2731_ ;
wire _2311_ ;
wire _3936_ ;
wire _3516_ ;
wire _8974_ ;
wire _8554_ ;
wire _8134_ ;
wire _9759_ ;
wire _9339_ ;
wire _4894_ ;
wire _4474_ ;
wire _4054_ ;
wire _913_ ;
wire _5679_ ;
wire _5259_ ;
wire _6620_ ;
wire _6200_ ;
wire _9092_ ;
wire _1599_ ;
wire _1179_ ;
wire _7825_ ;
wire _7405_ ;
wire _2960_ ;
wire _2540_ ;
wire _2120_ ;
wire _11823_ ;
wire _11403_ ;
wire _3745_ ;
wire _3325_ ;
wire _8783_ ;
wire _8363_ ;
wire _1811_ ;
wire _9988_ ;
wire _9568_ ;
wire _9148_ ;
wire _4283_ ;
wire _722_ ;
wire _302_ ;
wire _5488_ ;
wire _5068_ ;
wire _7634_ ;
wire _7214_ ;
wire breg_18_bF$buf0 ;
wire breg_18_bF$buf1 ;
wire breg_18_bF$buf2 ;
wire breg_18_bF$buf3 ;
wire breg_18_bF$buf4 ;
wire breg_18_bF$buf5 ;
wire _11632_ ;
wire _11212_ ;
wire _8839_ ;
wire _8419_ ;
wire _3974_ ;
wire _3554_ ;
wire _3134_ ;
wire _4759_ ;
wire _4339_ ;
wire _5700_ ;
wire _8592_ ;
wire _8172_ ;
wire _38_ ;
wire _6905_ ;
wire _1620_ ;
wire _1200_ ;
wire _9797_ ;
wire _9377_ ;
wire _4092_ ;
wire _10903_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2825_ ;
wire _2405_ ;
wire _5297_ ;
wire _7863_ ;
wire _7443_ ;
wire _7023_ ;
wire _11861_ ;
wire _11441_ ;
wire _11021_ ;
wire _8648_ ;
wire _8228_ ;
wire _3783_ ;
wire _3363_ ;
wire _4988_ ;
wire _4568_ ;
wire _4148_ ;
wire _6714_ ;
wire _9186_ ;
wire _10712_ ;
wire _760_ ;
wire _340_ ;
wire _7919_ ;
wire _2634_ ;
wire _2214_ ;
wire _3839_ ;
wire _3419_ ;
wire _7672_ ;
wire _7252_ ;
wire _11670_ ;
wire _11250_ ;
wire _8877_ ;
wire _8457_ ;
wire _8037_ ;
wire _3592_ ;
wire _3172_ ;
wire _1905_ ;
wire _4797_ ;
wire _4377_ ;
wire _816_ ;
wire _76_ ;
wire _6943_ ;
wire _6523_ ;
wire _6103_ ;
wire _10941_ ;
wire _10521_ ;
wire _10101_ ;
wire _7728_ ;
wire _7308_ ;
wire _2863_ ;
wire _2443_ ;
wire _2023_ ;
wire _11726_ ;
wire _11306_ ;
wire _3648_ ;
wire _3228_ ;
wire _7481_ ;
wire _7061_ ;
wire _8686_ ;
wire _8266_ ;
wire _1714_ ;
wire _4186_ ;
wire _625_ ;
wire _205_ ;
wire _2919_ ;
wire _6752_ ;
wire _6332_ ;
wire _10750_ ;
wire _10330_ ;
wire _7957_ ;
wire _7537_ ;
wire _7117_ ;
wire _2562__bF$buf0 ;
wire _2562__bF$buf1 ;
wire _2562__bF$buf2 ;
wire _2672_ ;
wire _2562__bF$buf3 ;
wire _2252_ ;
wire _2562__bF$buf4 ;
wire clk_bF$buf10 ;
wire _11535_ ;
wire _11115_ ;
wire _3877_ ;
wire _3457_ ;
wire _3037_ ;
wire _7290_ ;
wire _5603_ ;
wire _8495_ ;
wire _8075_ ;
wire _6808_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _10806_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _6981_ ;
wire _6561_ ;
wire _6141_ ;
wire _7766_ ;
wire _7346_ ;
wire _2481_ ;
wire _2061_ ;
wire _11764_ ;
wire _11344_ ;
wire _3686_ ;
wire _3266_ ;
wire _9912_ ;
wire _5832_ ;
wire _5412_ ;
wire _6617_ ;
wire _1752_ ;
wire _1332_ ;
wire _9089_ ;
wire _10615_ ;
wire _663_ ;
wire _243_ ;
wire _2957_ ;
wire _2537_ ;
wire _2117_ ;
wire _6790_ ;
wire _6370_ ;
wire _7995_ ;
wire _7575_ ;
wire _7155_ ;
wire _2290_ ;
wire _11573_ ;
wire _11153_ ;
wire _3495_ ;
wire _3075_ ;
wire _9721_ ;
wire _9301_ ;
wire _1808_ ;
wire _5641_ ;
wire _5221_ ;
wire _719_ ;
wire _6846_ ;
wire _6426_ ;
wire _6006_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _10844_ ;
wire _10424_ ;
wire _10004_ ;
wire _892_ ;
wire _472_ ;
wire _2766_ ;
wire _2346_ ;
wire _11629_ ;
wire _11209_ ;
wire _4912_ ;
wire _7384_ ;
wire _11382_ ;
wire _8589_ ;
wire _8169_ ;
wire _9950_ ;
wire _9530_ ;
wire _9110_ ;
wire _1617_ ;
wire breg_21_bF$buf0 ;
wire breg_21_bF$buf1 ;
wire _4089_ ;
wire breg_21_bF$buf2 ;
wire breg_21_bF$buf3 ;
wire breg_21_bF$buf4 ;
wire _5870_ ;
wire _5450_ ;
wire _5030_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _6655_ ;
wire _6235_ ;
wire _1790_ ;
wire _1370_ ;
wire _10653_ ;
wire _10233_ ;
wire _281_ ;
wire _2995_ ;
wire _2575_ ;
wire _2155_ ;
wire _8801_ ;
wire _11858_ ;
wire _11438_ ;
wire _11018_ ;
wire _4721_ ;
wire _4301_ ;
wire _7193_ ;
wire _11191_ ;
wire _5926_ ;
wire _5506_ ;
wire _8398_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _10709_ ;
wire _757_ ;
wire _337_ ;
wire _6884_ ;
wire _6464_ ;
wire _6044_ ;
wire _10882_ ;
wire _10462_ ;
wire _10042_ ;
wire _7669_ ;
wire _7249_ ;
wire _2384_ ;
wire _8610_ ;
wire _11667_ ;
wire _11247_ ;
wire _3589_ ;
wire _3169_ ;
wire _9815_ ;
wire _4950_ ;
wire _4530_ ;
wire _4110_ ;
wire _5735_ ;
wire _5315_ ;
wire _1655_ ;
wire _1235_ ;
wire _10938_ ;
wire _10518_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _3801_ ;
wire _6693_ ;
wire _6273_ ;
wire _10691_ ;
wire _10271_ ;
wire _7898_ ;
wire _7478_ ;
wire _7058_ ;
wire _2193_ ;
wire _11896_ ;
wire _11476_ ;
wire _11056_ ;
wire _3398_ ;
wire _9624_ ;
wire _9204_ ;
wire _5964_ ;
wire _5544_ ;
wire _5124_ ;
wire _6749_ ;
wire _6329_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _10747_ ;
wire _10327_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _3610_ ;
wire _6082_ ;
wire _10080_ ;
wire _4815_ ;
wire _7287_ ;
wire _11285_ ;
wire _9853_ ;
wire _9433_ ;
wire _9013_ ;
wire _5773_ ;
wire _5353_ ;
wire areg_30_bF$buf0 ;
wire areg_30_bF$buf1 ;
wire areg_30_bF$buf2 ;
wire areg_30_bF$buf3 ;
wire areg_30_bF$buf4 ;
wire areg_30_bF$buf5 ;
wire _6978_ ;
wire _6558_ ;
wire _6138_ ;
wire _1693_ ;
wire _1273_ ;
wire _10976_ ;
wire _10556_ ;
wire _10136_ ;
wire _184_ ;
wire _2898_ ;
wire _2478_ ;
wire _2058_ ;
wire _8704_ ;
wire _9909_ ;
wire _4624_ ;
wire _4204_ ;
wire _7096_ ;
wire _11094_ ;
wire _5829_ ;
wire _5409_ ;
wire _9662_ ;
wire _9242_ ;
wire _1749_ ;
wire _1329_ ;
wire _5582_ ;
wire _5162_ ;
wire _6787_ ;
wire _6367_ ;
wire _1082_ ;
wire _10785_ ;
wire _10365_ ;
wire _2287_ ;
wire _8933_ ;
wire _8513_ ;
wire _9718_ ;
wire _4853_ ;
wire _4433_ ;
wire _4013_ ;
wire _5638_ ;
wire _5218_ ;
wire _9891_ ;
wire _9471_ ;
wire _9051_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _5391_ ;
wire _889_ ;
wire _469_ ;
wire _3704_ ;
wire _6596_ ;
wire _6176_ ;
wire _10594_ ;
wire _10174_ ;
wire _4909_ ;
wire _2096_ ;
wire _8742_ ;
wire _8322_ ;
wire _11799_ ;
wire _11379_ ;
wire _9947_ ;
wire _9527_ ;
wire _9107_ ;
wire _4662_ ;
wire _4242_ ;
wire _5867_ ;
wire _5447_ ;
wire _5027_ ;
wire _9280_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _3933_ ;
wire _3513_ ;
wire _4718_ ;
wire _8971_ ;
wire _8551_ ;
wire _8131_ ;
wire _11188_ ;
wire _9756_ ;
wire _9336_ ;
wire _4891_ ;
wire _4471_ ;
wire _4051_ ;
wire _910_ ;
wire _5676_ ;
wire _5256_ ;
wire _1596_ ;
wire _1176_ ;
wire _7822_ ;
wire _7402_ ;
wire _10879_ ;
wire _10459_ ;
wire _10039_ ;
wire _11820_ ;
wire _11400_ ;
wire _8607_ ;
wire _3742_ ;
wire _3322_ ;
wire _4947_ ;
wire _4527_ ;
wire _4107_ ;
wire _8780_ ;
wire _8360_ ;
wire _9985_ ;
wire _9565_ ;
wire _9145_ ;
wire _4280_ ;
wire _5485_ ;
wire _5065_ ;
wire _7631_ ;
wire _7211_ ;
wire _10688_ ;
wire _10268_ ;
wire _8836_ ;
wire _8416_ ;
wire _3971_ ;
wire _3551_ ;
wire _3131_ ;
wire _4756_ ;
wire _4336_ ;
wire _35_ ;
wire _6902_ ;
wire _9794_ ;
wire _9374_ ;
wire _10900_ ;
wire _2822_ ;
wire _2402_ ;
wire _5294_ ;
wire _3607_ ;
wire _6499_ ;
wire _6079_ ;
wire _7860_ ;
wire _7440_ ;
wire _7020_ ;
wire _10497_ ;
wire _10077_ ;
wire _8645_ ;
wire _8225_ ;
wire _3780_ ;
wire _3360_ ;
wire _4985_ ;
wire _4565_ ;
wire _4145_ ;
wire _6711_ ;
wire _9183_ ;
wire _7916_ ;
wire _2631_ ;
wire _2211_ ;
wire _3836_ ;
wire _3416_ ;
wire _8874_ ;
wire _8454_ ;
wire _8034_ ;
wire _1902_ ;
wire _9659_ ;
wire _9239_ ;
wire _4794_ ;
wire _4374_ ;
wire _813_ ;
wire _5999_ ;
wire _5579_ ;
wire _5159_ ;
wire _73_ ;
wire _6940_ ;
wire _6520_ ;
wire _6100_ ;
wire _1499_ ;
wire _1079_ ;
wire _7725_ ;
wire _7305_ ;
wire _2860_ ;
wire _2440_ ;
wire _2020_ ;
wire _11723_ ;
wire _11303_ ;
wire _3645_ ;
wire _3225_ ;
wire _8683_ ;
wire _8263_ ;
wire _1711_ ;
wire _9888_ ;
wire _9468_ ;
wire _9048_ ;
wire _4183_ ;
wire _622_ ;
wire _202_ ;
wire _2916_ ;
wire _5388_ ;
wire _7954_ ;
wire _7534_ ;
wire _7114_ ;
wire _11532_ ;
wire _11112_ ;
wire _8739_ ;
wire _8319_ ;
wire _3874_ ;
wire _3454_ ;
wire _3034_ ;
wire _4659_ ;
wire _4239_ ;
wire _5600_ ;
wire _8492_ ;
wire _8072_ ;
wire _6805_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _9697_ ;
wire _9277_ ;
wire _10803_ ;
wire _4551__bF$buf0 ;
wire _4551__bF$buf1 ;
wire _4551__bF$buf2 ;
wire _4551__bF$buf3 ;
wire _4551__bF$buf4 ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _5197_ ;
wire _3958__bF$buf0 ;
wire _3958__bF$buf1 ;
wire _7763_ ;
wire _3958__bF$buf2 ;
wire _7343_ ;
wire _3958__bF$buf3 ;
wire _11761_ ;
wire _11341_ ;
wire _8968_ ;
wire _8548_ ;
wire _8128_ ;
wire _3683_ ;
wire _3263_ ;
wire _4888_ ;
wire _4468_ ;
wire _4048_ ;
wire _907_ ;
wire _6614_ ;
wire _9086_ ;
wire _10612_ ;
wire _660_ ;
wire _240_ ;
wire _7819_ ;
wire _2954_ ;
wire _2534_ ;
wire _2114_ ;
wire _11817_ ;
wire _3739_ ;
wire _3319_ ;
wire _7992_ ;
wire _7572_ ;
wire _7152_ ;
wire _11570_ ;
wire _11150_ ;
wire _8777_ ;
wire _8357_ ;
wire _3492_ ;
wire _3072_ ;
wire _1805_ ;
wire _4697_ ;
wire _4277_ ;
wire _716_ ;
wire _6843_ ;
wire _6423_ ;
wire _6003_ ;
wire _10841_ ;
wire _10421_ ;
wire _10001_ ;
wire _7628_ ;
wire _7208_ ;
wire _2763_ ;
wire _2343_ ;
wire _11626_ ;
wire _11206_ ;
wire _3968_ ;
wire _3548_ ;
wire _3128_ ;
wire _7381_ ;
wire _8586_ ;
wire _8166_ ;
wire _1614_ ;
wire _4086_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2819_ ;
wire _6652_ ;
wire _6232_ ;
wire _10650_ ;
wire _10230_ ;
wire _7857_ ;
wire _7437_ ;
wire _7017_ ;
wire _2992_ ;
wire _2572_ ;
wire _2152_ ;
wire _11855_ ;
wire _11435_ ;
wire _11015_ ;
wire _3777_ ;
wire _3357_ ;
wire _7190_ ;
wire _5923_ ;
wire _5503_ ;
wire _8395_ ;
wire _6708_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _10706_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _6881_ ;
wire _6461_ ;
wire _6041_ ;
wire _7666_ ;
wire _7246_ ;
wire _2381_ ;
wire _11664_ ;
wire _11244_ ;
wire _3586_ ;
wire _3166_ ;
wire _9812_ ;
wire _5732_ ;
wire _5312_ ;
wire _6937_ ;
wire _6517_ ;
wire _1652_ ;
wire _1232_ ;
wire _10935_ ;
wire _10515_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2857_ ;
wire _2437_ ;
wire _2017_ ;
wire _6690_ ;
wire _6270_ ;
wire _7895_ ;
wire _7475_ ;
wire _7055_ ;
wire _2190_ ;
wire _11893_ ;
wire _11473_ ;
wire _11053_ ;
wire _3395_ ;
wire _9621_ ;
wire _9201_ ;
wire _1708_ ;
wire breg_13_bF$buf0 ;
wire breg_13_bF$buf1 ;
wire breg_13_bF$buf2 ;
wire breg_13_bF$buf3 ;
wire breg_13_bF$buf4 ;
wire _5961_ ;
wire _5541_ ;
wire _5121_ ;
wire _619_ ;
wire _6746_ ;
wire _6326_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _10744_ ;
wire _10324_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _11529_ ;
wire _11109_ ;
wire _4812_ ;
wire _7284_ ;
wire _11282_ ;
wire _8489_ ;
wire _8069_ ;
wire _9850_ ;
wire _9430_ ;
wire _9010_ ;
wire _1937_ ;
wire _1517_ ;
wire _5770_ ;
wire _5350_ ;
wire _848_ ;
wire _428_ ;
wire _6975_ ;
wire _6555_ ;
wire _6135_ ;
wire _1690_ ;
wire _1270_ ;
wire _10973_ ;
wire _10553_ ;
wire _10133_ ;
wire _181_ ;
wire _2895_ ;
wire _2475_ ;
wire _2055_ ;
wire _8701_ ;
wire _11758_ ;
wire _11338_ ;
wire _9906_ ;
wire _4621_ ;
wire _4201_ ;
wire _7093_ ;
wire _11091_ ;
wire _5826_ ;
wire _5406_ ;
wire _8298_ ;
wire _1746_ ;
wire _1326_ ;
wire _10609_ ;
wire _657_ ;
wire _237_ ;
wire _6686__bF$buf0 ;
wire _6686__bF$buf1 ;
wire _6686__bF$buf2 ;
wire _6686__bF$buf3 ;
wire _6784_ ;
wire _6364_ ;
wire _10782_ ;
wire _10362_ ;
wire _7989_ ;
wire _7569_ ;
wire _7149_ ;
wire _2284_ ;
wire _8930_ ;
wire _8510_ ;
wire _11567_ ;
wire _11147_ ;
wire _3489_ ;
wire _3069_ ;
wire _9715_ ;
wire _4850_ ;
wire _4430_ ;
wire _4010_ ;
wire _5635_ ;
wire _5215_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _10838_ ;
wire _10418_ ;
wire _886_ ;
wire _466_ ;
wire _3701_ ;
wire _6593_ ;
wire _6173_ ;
wire _10591_ ;
wire _10171_ ;
wire _4906_ ;
wire _7798_ ;
wire _7378_ ;
wire _2093_ ;
wire _11796_ ;
wire _11376_ ;
wire _3298_ ;
wire _9944_ ;
wire _9524_ ;
wire _9104_ ;
wire _5864_ ;
wire _5444_ ;
wire _5024_ ;
wire _6649_ ;
wire _6229_ ;
wire _1784_ ;
wire _1364_ ;
wire _10647_ ;
wire _10227_ ;
wire _695_ ;
wire _275_ ;
wire _2989_ ;
wire _2569_ ;
wire _2149_ ;
wire _3930_ ;
wire _3510_ ;
wire _4715_ ;
wire _7187_ ;
wire _11185_ ;
wire _9753_ ;
wire _9333_ ;
wire _5673_ ;
wire _5253_ ;
wire _6878_ ;
wire _6458_ ;
wire _6038_ ;
wire _1593_ ;
wire _1173_ ;
wire _10876_ ;
wire _10456_ ;
wire _10036_ ;
wire _2798_ ;
wire _2378_ ;
wire _8604_ ;
wire _9809_ ;
wire _4944_ ;
wire _4524_ ;
wire _4104_ ;
wire _5729_ ;
wire _5309_ ;
wire _9982_ ;
wire _9562_ ;
wire _9142_ ;
wire _1649_ ;
wire _1229_ ;
wire _5482_ ;
wire _5062_ ;
wire _6687_ ;
wire _6267_ ;
wire _10685_ ;
wire _10265_ ;
wire _2187_ ;
wire _8833_ ;
wire _8413_ ;
wire _9618_ ;
wire _4753_ ;
wire _4333_ ;
wire _5958_ ;
wire _5538_ ;
wire _5118_ ;
wire _32_ ;
wire _9791_ ;
wire _9371_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _5291_ ;
wire _789_ ;
wire _369_ ;
wire _3604_ ;
wire _6496_ ;
wire _6076_ ;
wire _10494_ ;
wire _10074_ ;
wire _4809_ ;
wire _8642_ ;
wire _8222_ ;
wire _11699_ ;
wire _11279_ ;
wire _9847_ ;
wire _9427_ ;
wire _9007_ ;
wire _4982_ ;
wire _4562_ ;
wire _4142_ ;
wire _5767_ ;
wire _5347_ ;
wire _9180_ ;
wire _1687_ ;
wire _1267_ ;
wire _7913_ ;
wire _598_ ;
wire _178_ ;
wire _3833_ ;
wire _3413_ ;
wire _4618_ ;
wire _8871_ ;
wire _8451_ ;
wire _8031_ ;
wire _11088_ ;
wire _9656_ ;
wire _9236_ ;
wire _4791_ ;
wire _4371_ ;
wire _810_ ;
wire _5996_ ;
wire _5576_ ;
wire _5156_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _7722_ ;
wire _7302_ ;
wire _10779_ ;
wire _10359_ ;
wire _11720_ ;
wire _11300_ ;
wire _8927_ ;
wire _8507_ ;
wire _3642_ ;
wire _3222_ ;
wire _4847_ ;
wire _4427_ ;
wire _4007_ ;
wire _8680_ ;
wire _8260_ ;
wire _9885_ ;
wire _9465_ ;
wire _9045_ ;
wire _4180_ ;
wire _2913_ ;
wire _5385_ ;
wire _7951_ ;
wire _7531_ ;
wire _7111_ ;
wire _10588_ ;
wire _10168_ ;
wire _8736_ ;
wire _8316_ ;
wire _3871_ ;
wire _3451_ ;
wire _3031_ ;
wire _4656_ ;
wire _4236_ ;
wire _6802_ ;
wire _9694_ ;
wire _9274_ ;
wire _10800_ ;
wire _2722_ ;
wire _2302_ ;
wire _5194_ ;
wire _3927_ ;
wire _3507_ ;
wire _6399_ ;
wire _7760_ ;
wire _7340_ ;
wire _10397_ ;
wire _8965_ ;
wire _8545_ ;
wire _8125_ ;
wire _3680_ ;
wire _3260_ ;
wire areg_15_bF$buf0 ;
wire areg_15_bF$buf1 ;
wire areg_15_bF$buf2 ;
wire areg_15_bF$buf3 ;
wire areg_15_bF$buf4 ;
wire _4885_ ;
wire _4465_ ;
wire _4045_ ;
wire _904_ ;
wire _6611_ ;
wire _9083_ ;
wire _7816_ ;
wire _2951_ ;
wire _2531_ ;
wire _2111_ ;
wire _11814_ ;
wire _3736_ ;
wire _3316_ ;
wire _8774_ ;
wire _8354_ ;
wire _1802_ ;
wire _9979_ ;
wire _9559_ ;
wire _9139_ ;
wire _4694_ ;
wire _4274_ ;
wire _713_ ;
wire _5899_ ;
wire _5479_ ;
wire _5059_ ;
wire _6840_ ;
wire _6420_ ;
wire _6000_ ;
wire _1399_ ;
wire _7625_ ;
wire _7205_ ;
wire _2760_ ;
wire _2340_ ;
wire _11623_ ;
wire _11203_ ;
wire _3965_ ;
wire _3545_ ;
wire _3125_ ;
wire _8583_ ;
wire _8163_ ;
wire _29_ ;
wire _1611_ ;
wire _9788_ ;
wire _9368_ ;
wire _4083_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _2816_ ;
wire _5288_ ;
wire _7854_ ;
wire _7434_ ;
wire _7014_ ;
wire _11852_ ;
wire _11432_ ;
wire _11012_ ;
wire _8639_ ;
wire _8219_ ;
wire _3774_ ;
wire _3354_ ;
wire _4979_ ;
wire _4559_ ;
wire _4139_ ;
wire _5920_ ;
wire _5500_ ;
wire _8392_ ;
wire _6705_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _9597_ ;
wire _9177_ ;
wire _10703_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _5097_ ;
wire _11908_ ;
wire _7663_ ;
wire _7243_ ;
wire _11661_ ;
wire _11241_ ;
wire _8868_ ;
wire _8448_ ;
wire _8028_ ;
wire _3583_ ;
wire _3163_ ;
wire _4788_ ;
wire _4368_ ;
wire _807_ ;
wire _67_ ;
wire _6934_ ;
wire _6514_ ;
wire _10932_ ;
wire _10512_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _7719_ ;
wire _2854_ ;
wire _2434_ ;
wire _2014_ ;
wire _11717_ ;
wire _3639_ ;
wire _3219_ ;
wire _7892_ ;
wire _7472_ ;
wire _7052_ ;
wire _11890_ ;
wire _11470_ ;
wire _11050_ ;
wire _8677_ ;
wire _8257_ ;
wire _3392_ ;
wire _1705_ ;
wire _4597_ ;
wire _4177_ ;
wire _616_ ;
wire _6743_ ;
wire _6323_ ;
wire _10741_ ;
wire _10321_ ;
wire _7948_ ;
wire _7528_ ;
wire _7108_ ;
wire _2663_ ;
wire _2243_ ;
wire _11526_ ;
wire _11106_ ;
wire _3868_ ;
wire _3448_ ;
wire _3028_ ;
wire _7281_ ;
wire _8486_ ;
wire _8066_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _6972_ ;
wire _6552_ ;
wire _6132_ ;
wire _10970_ ;
wire _10550_ ;
wire _10130_ ;
wire _7757_ ;
wire _7337_ ;
wire _2892_ ;
wire _2472_ ;
wire _2052_ ;
wire _11755_ ;
wire _11335_ ;
wire _3677_ ;
wire _3257_ ;
wire _9903_ ;
wire _7090_ ;
wire _5823_ ;
wire _5403_ ;
wire _8295_ ;
wire _6608_ ;
wire _1743_ ;
wire _1323_ ;
wire _10606_ ;
wire _654_ ;
wire _234_ ;
wire _2948_ ;
wire _2528_ ;
wire _2108_ ;
wire _6781_ ;
wire _6361_ ;
wire _7986_ ;
wire _7566_ ;
wire _7146_ ;
wire _2281_ ;
wire _11564_ ;
wire _11144_ ;
wire _3486_ ;
wire _3066_ ;
wire _9712_ ;
wire _5632_ ;
wire _5212_ ;
wire _6837_ ;
wire _6417_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _10835_ ;
wire _10415_ ;
wire _883_ ;
wire _463_ ;
wire _2757_ ;
wire _2337_ ;
wire _6590_ ;
wire _6170_ ;
wire _4903_ ;
wire _7795_ ;
wire _7375_ ;
wire _2090_ ;
wire _11793_ ;
wire _11373_ ;
wire _3295_ ;
wire _9941_ ;
wire _9521_ ;
wire _9101_ ;
wire _1608_ ;
wire _5861_ ;
wire _5441_ ;
wire _5021_ ;
wire _939_ ;
wire _519_ ;
wire _6646_ ;
wire _6226_ ;
wire _1781_ ;
wire _1361_ ;
wire _10644_ ;
wire _10224_ ;
wire _692_ ;
wire _272_ ;
wire _2986_ ;
wire _2566_ ;
wire _2146_ ;
wire _11849_ ;
wire _11429_ ;
wire _11009_ ;
wire _4712_ ;
wire _7184_ ;
wire _11182_ ;
wire _5917_ ;
wire _8389_ ;
wire _9750_ ;
wire _9330_ ;
wire _1837_ ;
wire _1417_ ;
wire _5670_ ;
wire _5250_ ;
wire _748_ ;
wire _328_ ;
wire _6875_ ;
wire _6455_ ;
wire _6035_ ;
wire _1590_ ;
wire _1170_ ;
wire _10873_ ;
wire _10453_ ;
wire _10033_ ;
wire _2795_ ;
wire _2375_ ;
wire _8601_ ;
wire _11658_ ;
wire _11238_ ;
wire _9806_ ;
wire _4941_ ;
wire _4521_ ;
wire _4101_ ;
wire _5726_ ;
wire _5306_ ;
wire _8198_ ;
wire _1646_ ;
wire _1226_ ;
wire _4258__bF$buf0 ;
wire _4258__bF$buf1 ;
wire _4258__bF$buf2 ;
wire _4258__bF$buf3 ;
wire _10929_ ;
wire _10509_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _6684_ ;
wire _6264_ ;
wire _10682_ ;
wire _10262_ ;
wire _7889_ ;
wire _7469_ ;
wire _7049_ ;
wire _2184_ ;
wire _8830_ ;
wire _8410_ ;
wire _11887_ ;
wire _11467_ ;
wire _11047_ ;
wire _3389_ ;
wire _9615_ ;
wire _4750_ ;
wire _4330_ ;
wire _5955_ ;
wire _5535_ ;
wire _5115_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _10738_ ;
wire _10318_ ;
wire _786_ ;
wire _366_ ;
wire _3601_ ;
wire _6493_ ;
wire _6073_ ;
wire _10491_ ;
wire _10071_ ;
wire _4806_ ;
wire _7698_ ;
wire _7278_ ;
wire _11696_ ;
wire _11276_ ;
wire _3198_ ;
wire _9844_ ;
wire _9424_ ;
wire _9004_ ;
wire _5764_ ;
wire _5344_ ;
wire _6969_ ;
wire _6549_ ;
wire _6129_ ;
wire _1684_ ;
wire _1264_ ;
wire _7910_ ;
wire _10967_ ;
wire _10547_ ;
wire _10127_ ;
wire _595_ ;
wire _175_ ;
wire _2889_ ;
wire _2469_ ;
wire _2049_ ;
wire _3830_ ;
wire _3410_ ;
wire _4615_ ;
wire _7087_ ;
wire _11085_ ;
wire _9653_ ;
wire _9233_ ;
wire _5993_ ;
wire _5573_ ;
wire _5153_ ;
wire _6778_ ;
wire _6358_ ;
wire _1493_ ;
wire _1073_ ;
wire _10776_ ;
wire _10356_ ;
wire _2698_ ;
wire _2278_ ;
wire _8924_ ;
wire _8504_ ;
wire _9709_ ;
wire _4844_ ;
wire _4424_ ;
wire _4004_ ;
wire _5629_ ;
wire _5209_ ;
wire _9882_ ;
wire _9462_ ;
wire _9042_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2910_ ;
wire _5382_ ;
wire _6587_ ;
wire _6167_ ;
wire _10585_ ;
wire _10165_ ;
wire _2087_ ;
wire _8733_ ;
wire _8313_ ;
wire _9938_ ;
wire _9518_ ;
wire _4653_ ;
wire _4233_ ;
wire _5858_ ;
wire _5438_ ;
wire _5018_ ;
wire _9691_ ;
wire _9271_ ;
wire _1778_ ;
wire _1358_ ;
wire _5191_ ;
wire _689_ ;
wire _269_ ;
wire _3924_ ;
wire _3504_ ;
wire _6396_ ;
wire _10394_ ;
wire _4709_ ;
wire _8962_ ;
wire _8542_ ;
wire _8122_ ;
wire _11599_ ;
wire _11179_ ;
wire _9747_ ;
wire _9327_ ;
wire _4882_ ;
wire _4462_ ;
wire _4042_ ;
wire _901_ ;
wire _5667_ ;
wire _5247_ ;
wire _9080_ ;
wire _1587_ ;
wire _1167_ ;
wire _7813_ ;
wire _498_ ;
wire _11811_ ;
wire _3733_ ;
wire _3313_ ;
wire _4938_ ;
wire _4518_ ;
wire _8771_ ;
wire _8351_ ;
wire _9976_ ;
wire _9556_ ;
wire _9136_ ;
wire _4691_ ;
wire _4271_ ;
wire _710_ ;
wire _5896_ ;
wire _5476_ ;
wire _5056_ ;
wire _1396_ ;
wire _7622_ ;
wire _7202_ ;
wire _10679_ ;
wire _10259_ ;
wire _11620_ ;
wire _11200_ ;
wire _8827_ ;
wire _8407_ ;
wire _3962_ ;
wire _3542_ ;
wire _3122_ ;
wire _4747_ ;
wire _4327_ ;
wire _8580_ ;
wire _8160_ ;
wire _26_ ;
wire _9785_ ;
wire _9365_ ;
wire _4080_ ;
wire _2813_ ;
wire _5285_ ;
wire _6050__bF$buf0 ;
wire _6050__bF$buf1 ;
wire _6050__bF$buf2 ;
wire _6050__bF$buf3 ;
wire _7851_ ;
wire _7431_ ;
wire _7011_ ;
wire _10488_ ;
wire _10068_ ;
wire _8636_ ;
wire _8216_ ;
wire _3771_ ;
wire _3351_ ;
wire _4976_ ;
wire _4556_ ;
wire _4136_ ;
wire areg_26_bF$buf0 ;
wire areg_26_bF$buf1 ;
wire areg_26_bF$buf2 ;
wire areg_26_bF$buf3 ;
wire areg_26_bF$buf4 ;
wire _6702_ ;
wire _9594_ ;
wire _9174_ ;
wire _10700_ ;
wire _7907_ ;
wire _2622_ ;
wire _2202_ ;
wire _5094_ ;
wire _11905_ ;
wire _3827_ ;
wire _3407_ ;
wire _6299_ ;
wire _7660_ ;
wire _7240_ ;
wire _10297_ ;
wire _8865_ ;
wire _8445_ ;
wire _8025_ ;
wire _3580_ ;
wire _3160_ ;
wire _4785_ ;
wire _4365_ ;
wire _804_ ;
wire _64_ ;
wire _6931_ ;
wire _6511_ ;
wire _7716_ ;
wire _2851_ ;
wire _2431_ ;
wire _2011_ ;
wire _11714_ ;
wire _3636_ ;
wire _3216_ ;
wire _8674_ ;
wire _8254_ ;
wire _1702_ ;
wire _9879_ ;
wire _9459_ ;
wire _9039_ ;
wire _4594_ ;
wire _4174_ ;
wire _613_ ;
wire _2907_ ;
wire _5799_ ;
wire _5379_ ;
wire _6740_ ;
wire _6320_ ;
wire _1299_ ;
wire _7945_ ;
wire _7525_ ;
wire _7105_ ;
wire _2660_ ;
wire _2240_ ;
wire _11523_ ;
wire _11103_ ;
wire _3865_ ;
wire _3445_ ;
wire _3025_ ;
wire _8483_ ;
wire _8063_ ;
wire _1931_ ;
wire _1511_ ;
wire _9688_ ;
wire _9268_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _5188_ ;
wire _7754_ ;
wire _7334_ ;
wire _11752_ ;
wire _11332_ ;
wire _8959_ ;
wire _8539_ ;
wire _8119_ ;
wire _3674_ ;
wire _3254_ ;
wire _9900_ ;
wire _4879_ ;
wire _4459_ ;
wire _4039_ ;
wire _5820_ ;
wire _5400_ ;
wire _8292_ ;
wire _6605_ ;
wire _1740_ ;
wire _1320_ ;
wire _9497_ ;
wire _9077_ ;
wire _10603_ ;
wire _651_ ;
wire _231_ ;
wire _2945_ ;
wire areg_8_bF$buf0 ;
wire _2525_ ;
wire areg_8_bF$buf1 ;
wire _2105_ ;
wire areg_8_bF$buf2 ;
wire areg_8_bF$buf3 ;
wire areg_8_bF$buf4 ;
wire _11808_ ;
wire _7983_ ;
wire _7563_ ;
wire _7143_ ;
wire _11561_ ;
wire _11141_ ;
wire _8768_ ;
wire _8348_ ;
wire _3483_ ;
wire _3063_ ;
wire _4688_ ;
wire _4268_ ;
wire _707_ ;
wire _6834_ ;
wire _6414_ ;
wire _10832_ ;
wire _10412_ ;
wire _880_ ;
wire _460_ ;
wire _7619_ ;
wire _2754_ ;
wire _2334_ ;
wire _11617_ ;
wire _3959_ ;
wire _3539_ ;
wire _3119_ ;
wire _4900_ ;
wire _7792_ ;
wire _7372_ ;
wire _11790_ ;
wire _11370_ ;
wire _8997_ ;
wire _8577_ ;
wire _8157_ ;
wire _3292_ ;
wire _1605_ ;
wire _4497_ ;
wire _4077_ ;
wire _936_ ;
wire _516_ ;
wire _6643_ ;
wire _6223_ ;
wire _10641_ ;
wire _10221_ ;
wire _7848_ ;
wire _7428_ ;
wire _7008_ ;
wire _2983_ ;
wire _2563_ ;
wire _2143_ ;
wire _11846_ ;
wire _11426_ ;
wire _11006_ ;
wire _3768_ ;
wire _3348_ ;
wire _7181_ ;
wire _5914_ ;
wire _8386_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _6872_ ;
wire _6452_ ;
wire _6032_ ;
wire areg_10_bF$buf0 ;
wire areg_10_bF$buf1 ;
wire areg_10_bF$buf2 ;
wire areg_10_bF$buf3 ;
wire areg_10_bF$buf4 ;
wire _10870_ ;
wire _10450_ ;
wire _10030_ ;
wire _7657_ ;
wire _7237_ ;
wire _2792_ ;
wire _2372_ ;
wire _11655_ ;
wire _11235_ ;
wire _3997_ ;
wire _3577_ ;
wire _3157_ ;
wire _9803_ ;
wire _5723_ ;
wire _5303_ ;
wire _8195_ ;
wire _6928_ ;
wire _6508_ ;
wire _1643_ ;
wire _1223_ ;
wire _10926_ ;
wire _10506_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2848_ ;
wire _2428_ ;
wire _2008_ ;
wire _6681_ ;
wire _6261_ ;
wire _7886_ ;
wire _7466_ ;
wire _7046_ ;
wire _2181_ ;
wire _11884_ ;
wire _11464_ ;
wire _11044_ ;
wire _3386_ ;
wire _9612_ ;
wire _5952_ ;
wire _5532_ ;
wire _5112_ ;
wire _6737_ ;
wire _6317_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _10735_ ;
wire _10315_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2362__bF$buf0 ;
wire _2237_ ;
wire _2362__bF$buf1 ;
wire _2362__bF$buf2 ;
wire _2362__bF$buf3 ;
wire _2362__bF$buf4 ;
wire _2362__bF$buf5 ;
wire _6490_ ;
wire _6070_ ;
wire _4803_ ;
wire _7695_ ;
wire _7275_ ;
wire _11693_ ;
wire _11273_ ;
wire _3195_ ;
wire _9841_ ;
wire _9421_ ;
wire _9001_ ;
wire _1928_ ;
wire _1508_ ;
wire _5761_ ;
wire _5341_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _6966_ ;
wire _6546_ ;
wire _6126_ ;
wire _1681_ ;
wire _1261_ ;
wire _10964_ ;
wire _10544_ ;
wire _10124_ ;
wire _592_ ;
wire _172_ ;
wire _2886_ ;
wire _2466_ ;
wire _2046_ ;
wire _11749_ ;
wire _11329_ ;
wire _4612_ ;
wire _7084_ ;
wire _11082_ ;
wire _5817_ ;
wire _8289_ ;
wire _9650_ ;
wire _9230_ ;
wire _1737_ ;
wire _1317_ ;
wire _5990_ ;
wire _5570_ ;
wire _5150_ ;
wire _648_ ;
wire _228_ ;
wire _6775_ ;
wire _6355_ ;
wire _1490_ ;
wire _1070_ ;
wire _10773_ ;
wire _10353_ ;
wire _2695_ ;
wire _2275_ ;
wire _8921_ ;
wire _8501_ ;
wire _11558_ ;
wire _11138_ ;
wire _9706_ ;
wire _4841_ ;
wire _4421_ ;
wire _4001_ ;
wire _5626_ ;
wire _5206_ ;
wire _8098_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _10829_ ;
wire _10409_ ;
wire _877_ ;
wire _457_ ;
wire _6584_ ;
wire _6164_ ;
wire _10582_ ;
wire _10162_ ;
wire _7789_ ;
wire _7369_ ;
wire _2084_ ;
wire _8730_ ;
wire _8310_ ;
wire _11787_ ;
wire _11367_ ;
wire _3289_ ;
wire _9935_ ;
wire _9515_ ;
wire _4650_ ;
wire _4230_ ;
wire _5855_ ;
wire _5435_ ;
wire _5015_ ;
wire _1775_ ;
wire _1355_ ;
wire _10638_ ;
wire _10218_ ;
wire _686_ ;
wire _266_ ;
wire _3921_ ;
wire _3501_ ;
wire _6393_ ;
wire _10391_ ;
wire _4706_ ;
wire _7598_ ;
wire _7178_ ;
wire _11596_ ;
wire _11176_ ;
wire _3098_ ;
wire _9744_ ;
wire _9324_ ;
wire _5664_ ;
wire _5244_ ;
wire _6869_ ;
wire _6449_ ;
wire _6029_ ;
wire _1584_ ;
wire _1164_ ;
wire _7810_ ;
wire _10867_ ;
wire _10447_ ;
wire _10027_ ;
wire _495_ ;
wire _2789_ ;
wire _2369_ ;
wire _3730_ ;
wire _3310_ ;
wire _4935_ ;
wire _4515_ ;
wire _9973_ ;
wire _9553_ ;
wire _9133_ ;
wire _5893_ ;
wire _5473_ ;
wire _5053_ ;
wire _6678_ ;
wire _6258_ ;
wire _1393_ ;
wire _10676_ ;
wire _10256_ ;
wire _2598_ ;
wire _2178_ ;
wire _8824_ ;
wire _8404_ ;
wire _9609_ ;
wire _4744_ ;
wire _4324_ ;
wire breg_28_bF$buf0 ;
wire breg_28_bF$buf1 ;
wire breg_28_bF$buf2 ;
wire breg_28_bF$buf3 ;
wire breg_28_bF$buf4 ;
wire breg_28_bF$buf5 ;
wire _5949_ ;
wire _5529_ ;
wire _5109_ ;
wire _23_ ;
wire _9782_ ;
wire _9362_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _2810_ ;
wire _5282_ ;
wire _6487_ ;
wire _6067_ ;
wire _10485_ ;
wire _10065_ ;
wire breg_6_bF$buf0 ;
wire breg_6_bF$buf1 ;
wire breg_6_bF$buf2 ;
wire breg_6_bF$buf3 ;
wire breg_6_bF$buf4 ;
wire breg_6_bF$buf5 ;
wire _8633_ ;
wire _8213_ ;
wire _9838_ ;
wire _9418_ ;
wire _4973_ ;
wire _4553_ ;
wire _4133_ ;
wire _5758_ ;
wire _5338_ ;
wire _9591_ ;
wire _9171_ ;
wire _1678_ ;
wire _1258_ ;
wire _7904_ ;
wire _5091_ ;
wire _589_ ;
wire _169_ ;
wire _11902_ ;
wire _3824_ ;
wire _3404_ ;
wire _6296_ ;
wire _10294_ ;
wire _4609_ ;
wire _8862_ ;
wire _8442_ ;
wire _8022_ ;
wire _11499_ ;
wire _11079_ ;
wire _9647_ ;
wire _9227_ ;
wire _4782_ ;
wire _4362_ ;
wire _801_ ;
wire _5987_ ;
wire _5567_ ;
wire _5147_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _7713_ ;
wire _398_ ;
wire _11711_ ;
wire _8918_ ;
wire _3633_ ;
wire _3213_ ;
wire _4838_ ;
wire _4418_ ;
wire _8671_ ;
wire _8251_ ;
wire _9876_ ;
wire _9456_ ;
wire _9036_ ;
wire _4591_ ;
wire _4171_ ;
wire _610_ ;
wire _2904_ ;
wire _5796_ ;
wire _5376_ ;
wire _1296_ ;
wire _7942_ ;
wire _7522_ ;
wire _7102_ ;
wire _10999_ ;
wire _10579_ ;
wire _10159_ ;
wire _11520_ ;
wire _11100_ ;
wire _8727_ ;
wire _8307_ ;
wire _3862_ ;
wire _3442_ ;
wire _3022_ ;
wire _4647_ ;
wire _4227_ ;
wire _8480_ ;
wire _8060_ ;
wire _9685_ ;
wire _9265_ ;
wire _2713_ ;
wire _5185_ ;
wire _3918_ ;
wire _7751_ ;
wire _7331_ ;
wire _10388_ ;
wire _8956_ ;
wire _8536_ ;
wire _8116_ ;
wire _3671_ ;
wire _3251_ ;
wire _4876_ ;
wire _4456_ ;
wire _4036_ ;
wire _6602_ ;
wire _9494_ ;
wire _9074_ ;
wire _10600_ ;
wire _7807_ ;
wire _2942_ ;
wire _2522_ ;
wire _2102_ ;
wire _11805_ ;
wire _3727_ ;
wire _3307_ ;
wire _6199_ ;
wire _7980_ ;
wire _7560_ ;
wire _7140_ ;
wire _10197_ ;
wire _8765_ ;
wire _8345_ ;
wire _3480_ ;
wire _3060_ ;
wire _4685_ ;
wire _4265_ ;
wire _704_ ;
wire _6831_ ;
wire _6411_ ;
wire _7616_ ;
wire _2751_ ;
wire _2331_ ;
wire _11614_ ;
wire _3956_ ;
wire _3536_ ;
wire _3116_ ;
wire _8994_ ;
wire _8574_ ;
wire _8154_ ;
wire _1602_ ;
wire _9779_ ;
wire _9359_ ;
wire _4494_ ;
wire _4074_ ;
wire _933_ ;
wire _513_ ;
wire _2807_ ;
wire _5699_ ;
wire _5279_ ;
wire _6640_ ;
wire _6220_ ;
wire _1199_ ;
wire _7845_ ;
wire _7425_ ;
wire _7005_ ;
wire _2980_ ;
wire _2560_ ;
wire _2140_ ;
wire _11843_ ;
wire _11423_ ;
wire _11003_ ;
wire _3765_ ;
wire _3345_ ;
wire _5911_ ;
wire _8383_ ;
wire _1831_ ;
wire _1411_ ;
wire _9588_ ;
wire _9168_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _5088_ ;
wire _7654_ ;
wire _7234_ ;
wire _11652_ ;
wire _11232_ ;
wire _8859_ ;
wire _8439_ ;
wire _8019_ ;
wire _3994_ ;
wire _3574_ ;
wire _3154_ ;
wire _9800_ ;
wire _4779_ ;
wire _4359_ ;
wire _5720_ ;
wire _5300_ ;
wire _8192_ ;
wire _58_ ;
wire _6925_ ;
wire _6505_ ;
wire _1640_ ;
wire _1220_ ;
wire _9397_ ;
wire _10923_ ;
wire _10503_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2845_ ;
wire _2425_ ;
wire _2005_ ;
wire _11708_ ;
wire _7883_ ;
wire _7463_ ;
wire _7043_ ;
wire _11881_ ;
wire _11461_ ;
wire _11041_ ;
wire _8668_ ;
wire _8248_ ;
wire _3383_ ;
wire _4588_ ;
wire _4168_ ;
wire _607_ ;
wire _6734_ ;
wire _6314_ ;
wire _10732_ ;
wire _10312_ ;
wire _780_ ;
wire _360_ ;
wire _7939_ ;
wire _7519_ ;
wire _2654_ ;
wire _2234_ ;
wire _11517_ ;
wire _3859_ ;
wire _3439_ ;
wire _3019_ ;
wire _4800_ ;
wire _7692_ ;
wire _7272_ ;
wire _11690_ ;
wire _11270_ ;
wire _8897_ ;
wire _8477_ ;
wire _8057_ ;
wire _3192_ ;
wire _1925_ ;
wire _1505_ ;
wire _4397_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _6963_ ;
wire _6543_ ;
wire _6123_ ;
wire _10961_ ;
wire _10541_ ;
wire _10121_ ;
wire _7748_ ;
wire _7328_ ;
wire _2883_ ;
wire _2463_ ;
wire _2043_ ;
wire areg_21_bF$buf0 ;
wire areg_21_bF$buf1 ;
wire areg_21_bF$buf2 ;
wire areg_21_bF$buf3 ;
wire areg_21_bF$buf4 ;
wire _11746_ ;
wire _11326_ ;
wire _3668_ ;
wire _3248_ ;
wire _7081_ ;
wire _5814_ ;
wire _8286_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2939_ ;
wire _2519_ ;
wire _6772_ ;
wire _6352_ ;
wire _10770_ ;
wire _10350_ ;
wire _7977_ ;
wire _7557_ ;
wire _7137_ ;
wire _2692_ ;
wire _2272_ ;
wire _11555_ ;
wire _11135_ ;
wire _3897_ ;
wire _3477_ ;
wire _3057_ ;
wire _9703_ ;
wire _5623_ ;
wire _5203_ ;
wire _8095_ ;
wire _6828_ ;
wire _6408_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _10826_ ;
wire _10406_ ;
wire _874_ ;
wire _454_ ;
wire _2748_ ;
wire _2328_ ;
wire _6581_ ;
wire _6161_ ;
wire _7786_ ;
wire _7366_ ;
wire _2081_ ;
wire _11784_ ;
wire _11364_ ;
wire _3286_ ;
wire _9932_ ;
wire _9512_ ;
wire _5852_ ;
wire _5432_ ;
wire _5012_ ;
wire _6637_ ;
wire _6217_ ;
wire _1772_ ;
wire _1352_ ;
wire _10635_ ;
wire _10215_ ;
wire _683_ ;
wire _263_ ;
wire _2977_ ;
wire _2557_ ;
wire _2137_ ;
wire _6390_ ;
wire _4703_ ;
wire _7595_ ;
wire _7175_ ;
wire _11593_ ;
wire _11173_ ;
wire _5908_ ;
wire _3095_ ;
wire _9741_ ;
wire _9321_ ;
wire _1828_ ;
wire _1408_ ;
wire _5661_ ;
wire _5241_ ;
wire _739_ ;
wire _319_ ;
wire _6866_ ;
wire _6446_ ;
wire _6026_ ;
wire _1581_ ;
wire _1161_ ;
wire _10864_ ;
wire _10444_ ;
wire _10024_ ;
wire _492_ ;
wire _2786_ ;
wire _2366_ ;
wire _11649_ ;
wire _11229_ ;
wire _4932_ ;
wire _4512_ ;
wire areg_3_bF$buf0 ;
wire areg_3_bF$buf1 ;
wire areg_3_bF$buf2 ;
wire areg_3_bF$buf3 ;
wire areg_3_bF$buf4 ;
wire _5717_ ;
wire _8189_ ;
wire _9970_ ;
wire _9550_ ;
wire _9130_ ;
wire _1637_ ;
wire _1217_ ;
wire _5890_ ;
wire _5470_ ;
wire _5050_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _6675_ ;
wire _6255_ ;
wire _1390_ ;
wire _10673_ ;
wire _10253_ ;
wire _2595_ ;
wire _2175_ ;
wire _8821_ ;
wire _8401_ ;
wire _11878_ ;
wire _11458_ ;
wire _11038_ ;
wire _9606_ ;
wire _4741_ ;
wire _4321_ ;
wire _7217__bF$buf0 ;
wire _7217__bF$buf1 ;
wire _7217__bF$buf2 ;
wire _7217__bF$buf3 ;
wire _7217__bF$buf4 ;
wire _5946_ ;
wire _5526_ ;
wire _5106_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _10729_ ;
wire _10309_ ;
wire _777_ ;
wire _357_ ;
wire _6484_ ;
wire _6064_ ;
wire _10482_ ;
wire _10062_ ;
wire _7689_ ;
wire _7269_ ;
wire _8630_ ;
wire _8210_ ;
wire _11687_ ;
wire _11267_ ;
wire _3189_ ;
wire _9835_ ;
wire _9415_ ;
wire _4970_ ;
wire _4550_ ;
wire _4130_ ;
wire _5755_ ;
wire _5335_ ;
wire _1675_ ;
wire _1255_ ;
wire _7901_ ;
wire _10958_ ;
wire _10538_ ;
wire _10118_ ;
wire _586_ ;
wire _166_ ;
wire _3821_ ;
wire _3401_ ;
wire _6293_ ;
wire _10291_ ;
wire _4606_ ;
wire _7498_ ;
wire _7078_ ;
wire _11496_ ;
wire _11076_ ;
wire _9644_ ;
wire _9224_ ;
wire _5984_ ;
wire _5564_ ;
wire _5144_ ;
wire _6769_ ;
wire _6349_ ;
wire _1484_ ;
wire _1064_ ;
wire _7710_ ;
wire _10767_ ;
wire _10347_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _8915_ ;
wire _3630_ ;
wire _3210_ ;
wire _4835_ ;
wire _4415_ ;
wire _9873_ ;
wire _9453_ ;
wire _9033_ ;
wire _2901_ ;
wire _5793_ ;
wire _5373_ ;
wire _3781__bF$buf0 ;
wire _6998_ ;
wire _3781__bF$buf1 ;
wire _6578_ ;
wire _3781__bF$buf2 ;
wire _6158_ ;
wire _3781__bF$buf3 ;
wire _1293_ ;
wire _10996_ ;
wire _10576_ ;
wire _10156_ ;
wire _2498_ ;
wire _2078_ ;
wire _8724_ ;
wire _8304_ ;
wire _9929_ ;
wire _9509_ ;
wire _4644_ ;
wire _4224_ ;
wire _5849_ ;
wire _5429_ ;
wire _5009_ ;
wire _9682_ ;
wire _9262_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _5182_ ;
wire _3915_ ;
wire _6387_ ;
wire _10385_ ;
wire _8953_ ;
wire _8533_ ;
wire _8113_ ;
wire _9738_ ;
wire _9318_ ;
wire _4873_ ;
wire _4453_ ;
wire _4033_ ;
wire _5658_ ;
wire _5238_ ;
wire _9491_ ;
wire _9071_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _7804_ ;
wire _489_ ;
wire _11802_ ;
wire _3724_ ;
wire _3304_ ;
wire _6196_ ;
wire _10194_ ;
wire _4929_ ;
wire _4509_ ;
wire _8762_ ;
wire _8342_ ;
wire _11399_ ;
wire _9967_ ;
wire _9547_ ;
wire _9127_ ;
wire _4682_ ;
wire _4262_ ;
wire _701_ ;
wire _5887_ ;
wire _5467_ ;
wire _5047_ ;
wire _1387_ ;
wire _7613_ ;
wire _298_ ;
wire _11611_ ;
wire _8818_ ;
wire _3953_ ;
wire _3533_ ;
wire _3113_ ;
wire _4738_ ;
wire _4318_ ;
wire _8991_ ;
wire _8571_ ;
wire _8151_ ;
wire _17_ ;
wire _9776_ ;
wire _9356_ ;
wire _4491_ ;
wire _4071_ ;
wire _3253__bF$buf0 ;
wire _3253__bF$buf1 ;
wire _3253__bF$buf2 ;
wire _3253__bF$buf3 ;
wire _930_ ;
wire _510_ ;
wire _2804_ ;
wire _5696_ ;
wire _5276_ ;
wire _1196_ ;
wire _7842_ ;
wire _7422_ ;
wire _7002_ ;
wire _10899_ ;
wire _10479_ ;
wire _10059_ ;
wire _11840_ ;
wire _11420_ ;
wire _11000_ ;
wire _8627_ ;
wire _8207_ ;
wire _3762_ ;
wire _3342_ ;
wire _4967_ ;
wire _4547_ ;
wire _4127_ ;
wire _8380_ ;
wire _9585_ ;
wire _9165_ ;
wire _2613_ ;
wire _5085_ ;
wire _3818_ ;
wire _7651_ ;
wire _7231_ ;
wire _10288_ ;
wire _8856_ ;
wire _8436_ ;
wire _8016_ ;
wire _3991_ ;
wire _3571_ ;
wire _3151_ ;
wire _4776_ ;
wire _4356_ ;
wire _55_ ;
wire _6922_ ;
wire _6502_ ;
wire _9394_ ;
wire _10920_ ;
wire _10500_ ;
wire _7707_ ;
wire _2842_ ;
wire _2422_ ;
wire _2002_ ;
wire _11705_ ;
wire _3627_ ;
wire _3207_ ;
wire _6099_ ;
wire _7880_ ;
wire _7460_ ;
wire _7040_ ;
wire _10097_ ;
wire _8665_ ;
wire _8245_ ;
wire _3380_ ;
wire _3529__bF$buf0 ;
wire _3529__bF$buf1 ;
wire _3529__bF$buf2 ;
wire _3529__bF$buf3 ;
wire _3529__bF$buf4 ;
wire _4585_ ;
wire _4165_ ;
wire _604_ ;
wire _6731_ ;
wire _6311_ ;
wire _7936_ ;
wire _7516_ ;
wire _2651_ ;
wire _2231_ ;
wire breg_23_bF$buf0 ;
wire breg_23_bF$buf1 ;
wire breg_23_bF$buf2 ;
wire breg_23_bF$buf3 ;
wire _11514_ ;
wire _3856_ ;
wire _3436_ ;
wire _3016_ ;
wire _8894_ ;
wire _8474_ ;
wire _8054_ ;
wire _1922_ ;
wire _1502_ ;
wire _9679_ ;
wire _9259_ ;
wire _4394_ ;
wire breg_1_bF$buf0 ;
wire breg_1_bF$buf1 ;
wire breg_1_bF$buf2 ;
wire breg_1_bF$buf3 ;
wire _833_ ;
wire breg_1_bF$buf4 ;
wire _413_ ;
wire breg_1_bF$buf5 ;
wire breg_1_bF$buf6 ;
wire _2707_ ;
wire _5599_ ;
wire _5179_ ;
wire _93_ ;
wire _6960_ ;
wire _6540_ ;
wire _6120_ ;
wire _1099_ ;
wire _7745_ ;
wire _7325_ ;
wire _2880_ ;
wire _2460_ ;
wire _2040_ ;
wire _11743_ ;
wire _11323_ ;
wire _3665_ ;
wire _3245_ ;
wire _5811_ ;
wire _8283_ ;
wire _1731_ ;
wire _1311_ ;
wire _9488_ ;
wire _9068_ ;
wire _642_ ;
wire _222_ ;
wire _2936_ ;
wire _2516_ ;
wire _7974_ ;
wire _7554_ ;
wire _7520__bF$buf0 ;
wire _7134_ ;
wire _7520__bF$buf1 ;
wire _7520__bF$buf2 ;
wire _7520__bF$buf3 ;
wire _11552_ ;
wire _11132_ ;
wire _8759_ ;
wire _8339_ ;
wire _3894_ ;
wire _3474_ ;
wire _3054_ ;
wire _9700_ ;
wire _4679_ ;
wire _4259_ ;
wire _5620_ ;
wire _5200_ ;
wire _8092_ ;
wire _6825_ ;
wire _6405_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _9297_ ;
wire _10823_ ;
wire _10403_ ;
wire _871_ ;
wire _451_ ;
wire _2745_ ;
wire _2325_ ;
wire _11608_ ;
wire _7783_ ;
wire _7363_ ;
wire _11781_ ;
wire _11361_ ;
wire _8988_ ;
wire _8568_ ;
wire _8148_ ;
wire _3283_ ;
wire _4488_ ;
wire _4068_ ;
wire _927_ ;
wire _507_ ;
wire _6634_ ;
wire _6214_ ;
wire _10632_ ;
wire _10212_ ;
wire _680_ ;
wire _260_ ;
wire _7839_ ;
wire _7419_ ;
wire _2974_ ;
wire _2554_ ;
wire _2134_ ;
wire _11837_ ;
wire _11417_ ;
wire _3759_ ;
wire _3339_ ;
wire _4700_ ;
wire _7592_ ;
wire _7172_ ;
wire _11590_ ;
wire _11170_ ;
wire _5905_ ;
wire _8797_ ;
wire _8377_ ;
wire _3092_ ;
wire _1825_ ;
wire _1405_ ;
wire _4297_ ;
wire _736_ ;
wire _316_ ;
wire _6863_ ;
wire _6443_ ;
wire _6023_ ;
wire _10861_ ;
wire _10441_ ;
wire _10021_ ;
wire _7648_ ;
wire _7228_ ;
wire _2783_ ;
wire _2363_ ;
wire _11646_ ;
wire _11226_ ;
wire _3988_ ;
wire _3568_ ;
wire _3148_ ;
wire _5714_ ;
wire _8186_ ;
wire _6919_ ;
wire _1634_ ;
wire _1214_ ;
wire _10917_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2839_ ;
wire _2419_ ;
wire _6672_ ;
wire _6252_ ;
wire _10670_ ;
wire _10250_ ;
wire _7877_ ;
wire _7457_ ;
wire _7037_ ;
wire _2592_ ;
wire _2172_ ;
wire _11875_ ;
wire _11455_ ;
wire _11035_ ;
wire _3797_ ;
wire _3377_ ;
wire _9603_ ;
wire _5943_ ;
wire _5523_ ;
wire _5103_ ;
wire _6728_ ;
wire _6308_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _10726_ ;
wire _10306_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _6481_ ;
wire _6061_ ;
wire _7686_ ;
wire _7266_ ;
wire _11684_ ;
wire _11264_ ;
wire _3186_ ;
wire _9832_ ;
wire _9412_ ;
wire _1919_ ;
wire _5752_ ;
wire _5332_ ;
wire _6957_ ;
wire _6537_ ;
wire _6117_ ;
wire _1672_ ;
wire _1252_ ;
wire _10955_ ;
wire _10535_ ;
wire _10115_ ;
wire _583_ ;
wire _163_ ;
wire _2877_ ;
wire _2457_ ;
wire _2037_ ;
wire _6290_ ;
wire _4603_ ;
wire _7495_ ;
wire _7075_ ;
wire _11493_ ;
wire _11073_ ;
wire _5808_ ;
wire _5668__bF$buf0 ;
wire _5668__bF$buf1 ;
wire _5668__bF$buf2 ;
wire _5668__bF$buf3 ;
wire _9641_ ;
wire _5668__bF$buf4 ;
wire _9221_ ;
wire _5668__bF$buf5 ;
wire _1728_ ;
wire _1308_ ;
wire _5981_ ;
wire _5561_ ;
wire _5141_ ;
wire _639_ ;
wire _219_ ;
wire _6766_ ;
wire _6346_ ;
wire _1481_ ;
wire _1061_ ;
wire _10764_ ;
wire _10344_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _8912_ ;
wire _11549_ ;
wire _11129_ ;
wire _4832_ ;
wire _4412_ ;
wire _5617_ ;
wire _8089_ ;
wire _9870_ ;
wire _9450_ ;
wire _9030_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _5790_ ;
wire _5370_ ;
wire _868_ ;
wire _448_ ;
wire _6995_ ;
wire _6575_ ;
wire _6155_ ;
wire _1290_ ;
wire _10993_ ;
wire _10573_ ;
wire _10153_ ;
wire _6044__bF$buf0 ;
wire _6044__bF$buf1 ;
wire _6044__bF$buf2 ;
wire _6044__bF$buf3 ;
wire _6044__bF$buf4 ;
wire _6044__bF$buf5 ;
wire _2495_ ;
wire _2075_ ;
wire _8721_ ;
wire _8301_ ;
wire _11778_ ;
wire _11358_ ;
wire _9926_ ;
wire _9506_ ;
wire _4641_ ;
wire _4221_ ;
wire _5846_ ;
wire _5426_ ;
wire _5006_ ;
wire _1766_ ;
wire _1346_ ;
wire _10629_ ;
wire _10209_ ;
wire _677_ ;
wire _257_ ;
wire _3912_ ;
wire _6384_ ;
wire _10382_ ;
wire _7589_ ;
wire _7169_ ;
wire _8950_ ;
wire _8530_ ;
wire _8110_ ;
wire _11587_ ;
wire _11167_ ;
wire _3089_ ;
wire _9735_ ;
wire _9315_ ;
wire _4870_ ;
wire _4450_ ;
wire _4030_ ;
wire _5655_ ;
wire _5235_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _7801_ ;
wire _10858_ ;
wire _10438_ ;
wire _10018_ ;
wire _486_ ;
wire _3721_ ;
wire _3301_ ;
wire _6193_ ;
wire _10191_ ;
wire _4926_ ;
wire _4506_ ;
wire _7398_ ;
wire _11396_ ;
wire _9964_ ;
wire _9544_ ;
wire _9124_ ;
wire _5884_ ;
wire _5464_ ;
wire _5044_ ;
wire _6669_ ;
wire _6249_ ;
wire _1384_ ;
wire _7610_ ;
wire _10667_ ;
wire _10247_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _8815_ ;
wire _3950_ ;
wire _3530_ ;
wire _3110_ ;
wire _4735_ ;
wire _4315_ ;
wire _14_ ;
wire _9773_ ;
wire _9353_ ;
wire _2801_ ;
wire _5693_ ;
wire _5273_ ;
wire _6898_ ;
wire _6478_ ;
wire _6058_ ;
wire _1193_ ;
wire _10896_ ;
wire _10476_ ;
wire _10056_ ;
wire _2398_ ;
wire _8624_ ;
wire _8204_ ;
wire _9829_ ;
wire _9409_ ;
wire _4964_ ;
wire _4544_ ;
wire _4124_ ;
wire _5749_ ;
wire _5329_ ;
wire _9582_ ;
wire _9162_ ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _5082_ ;
wire _3815_ ;
wire _6287_ ;
wire _10285_ ;
wire _8853_ ;
wire _8433_ ;
wire _8013_ ;
wire _9638_ ;
wire _9218_ ;
wire _4773_ ;
wire _4353_ ;
wire _5978_ ;
wire _5558_ ;
wire _5138_ ;
wire _52_ ;
wire _9391_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _7704_ ;
wire _389_ ;
wire _11702_ ;
wire _8909_ ;
wire _3624_ ;
wire _3204_ ;
wire _6096_ ;
wire _10094_ ;
wire _4829_ ;
wire _4409_ ;
wire _8662_ ;
wire _2884__bF$buf0 ;
wire _8242_ ;
wire _2884__bF$buf1 ;
wire _2884__bF$buf2 ;
wire _2884__bF$buf3 ;
wire _11299_ ;
wire _9867_ ;
wire _9447_ ;
wire _9027_ ;
wire _4582_ ;
wire _4162_ ;
wire _601_ ;
wire _5787_ ;
wire _5367_ ;
wire _1287_ ;
wire _3402__bF$buf0 ;
wire _3402__bF$buf1 ;
wire _3402__bF$buf2 ;
wire _3402__bF$buf3 ;
wire _7933_ ;
wire _7513_ ;
wire _198_ ;
wire _11511_ ;
wire _8718_ ;
wire _3853_ ;
wire _3433_ ;
wire _3013_ ;
wire _4638_ ;
wire _4218_ ;
wire _8891_ ;
wire _8471_ ;
wire _8051_ ;
wire _9676_ ;
wire _9256_ ;
wire _4391_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _5596_ ;
wire _5176_ ;
wire _90_ ;
wire _3909_ ;
wire _1096_ ;
wire _7742_ ;
wire _7322_ ;
wire _10799_ ;
wire _10379_ ;
wire _11740_ ;
wire _11320_ ;
wire _8947_ ;
wire _8527_ ;
wire _8107_ ;
wire _3662_ ;
wire _3242_ ;
wire _4867_ ;
wire _4447_ ;
wire _4027_ ;
wire _8280_ ;
wire _9485_ ;
wire _9065_ ;
wire _2933_ ;
wire _2513_ ;
wire _3718_ ;
wire _7971_ ;
wire _7551_ ;
wire _7131_ ;
wire _10188_ ;
wire _8756_ ;
wire _8336_ ;
wire _3891_ ;
wire _3471_ ;
wire _3051_ ;
wire _4676_ ;
wire _4256_ ;
wire _6822_ ;
wire _6402_ ;
wire _9294_ ;
wire _10820_ ;
wire _10400_ ;
wire _7607_ ;
wire _2742_ ;
wire _2322_ ;
wire breg_15_bF$buf0 ;
wire breg_15_bF$buf1 ;
wire breg_15_bF$buf2 ;
wire breg_15_bF$buf3 ;
wire breg_15_bF$buf4 ;
wire _11605_ ;
wire breg_15_bF$buf5 ;
wire _3947_ ;
wire _3527_ ;
wire _3107_ ;
wire _8_ ;
wire _7780_ ;
wire _7360_ ;
wire _8985_ ;
wire _8565_ ;
wire _8145_ ;
wire _3280_ ;
wire _4485_ ;
wire _4065_ ;
wire _924_ ;
wire _504_ ;
wire _6631_ ;
wire _6211_ ;
wire _7836_ ;
wire _7416_ ;
wire _2971_ ;
wire _2551_ ;
wire _2131_ ;
wire _11834_ ;
wire _11414_ ;
wire _3756_ ;
wire _3336_ ;
wire _5902_ ;
wire _8794_ ;
wire _8374_ ;
wire _1822_ ;
wire _1402_ ;
wire _9999_ ;
wire _9579_ ;
wire _9159_ ;
wire _4294_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _5499_ ;
wire _5079_ ;
wire _6860_ ;
wire _6440_ ;
wire _6020_ ;
wire _7645_ ;
wire _7225_ ;
wire _2780_ ;
wire _2360_ ;
wire _11643_ ;
wire _11223_ ;
wire _3985_ ;
wire _3565_ ;
wire _3145_ ;
wire _5711_ ;
wire _8183_ ;
wire _49_ ;
wire _6916_ ;
wire _1631_ ;
wire _1211_ ;
wire _9388_ ;
wire _10914_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2836_ ;
wire _2416_ ;
wire _7874_ ;
wire _7454_ ;
wire _7034_ ;
wire _11872_ ;
wire _11452_ ;
wire _11032_ ;
wire _8659_ ;
wire _8239_ ;
wire _3794_ ;
wire _3374_ ;
wire _9600_ ;
wire _4999_ ;
wire _4579_ ;
wire _4159_ ;
wire _5940_ ;
wire _5520_ ;
wire _5100_ ;
wire _6725_ ;
wire _6305_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _9197_ ;
wire _10723_ ;
wire _10303_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _11508_ ;
wire _7683_ ;
wire _7263_ ;
wire _11681_ ;
wire _11261_ ;
wire _8888_ ;
wire _8468_ ;
wire _8048_ ;
wire _3183_ ;
wire _1916_ ;
wire _4388_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _6954_ ;
wire _6534_ ;
wire _6114_ ;
wire _10952_ ;
wire _10532_ ;
wire _10112_ ;
wire _580_ ;
wire _160_ ;
wire _7739_ ;
wire _7319_ ;
wire _2874_ ;
wire _2454_ ;
wire _2034_ ;
wire _11737_ ;
wire _11317_ ;
wire _3659_ ;
wire _3239_ ;
wire _4600_ ;
wire _7492_ ;
wire _7072_ ;
wire _11490_ ;
wire _11070_ ;
wire _5805_ ;
wire _8697_ ;
wire _8277_ ;
wire _1725_ ;
wire _1305_ ;
wire _4197_ ;
wire _636_ ;
wire _216_ ;
wire _6763_ ;
wire _6343_ ;
wire _10761_ ;
wire _10341_ ;
wire _7968_ ;
wire _7548_ ;
wire _7128_ ;
wire _2683_ ;
wire _2263_ ;
wire _11546_ ;
wire _11126_ ;
wire _3888_ ;
wire _3468_ ;
wire _3048_ ;
wire _5614_ ;
wire _8086_ ;
wire _6819_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _10817_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _6992_ ;
wire _6572_ ;
wire _6152_ ;
wire _10990_ ;
wire _10570_ ;
wire _10150_ ;
wire _7777_ ;
wire _7357_ ;
wire _2492_ ;
wire _2072_ ;
wire _11775_ ;
wire _11355_ ;
wire _3697_ ;
wire _3277_ ;
wire _9923_ ;
wire _9503_ ;
wire _5843_ ;
wire _5423_ ;
wire _5003_ ;
wire _6628_ ;
wire _6208_ ;
wire _1763_ ;
wire _1343_ ;
wire _10626_ ;
wire _10206_ ;
wire _674_ ;
wire _254_ ;
wire _2968_ ;
wire _2548_ ;
wire _2128_ ;
wire _6381_ ;
wire _7586_ ;
wire _7166_ ;
wire _11584_ ;
wire _11164_ ;
wire _3086_ ;
wire _9732_ ;
wire _9312_ ;
wire _1819_ ;
wire _5652_ ;
wire _5232_ ;
wire _6857_ ;
wire _6437_ ;
wire _6017_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _10855_ ;
wire _10435_ ;
wire _10015_ ;
wire _483_ ;
wire _2777_ ;
wire _2357_ ;
wire _6190_ ;
wire _4923_ ;
wire _4503_ ;
wire _7395_ ;
wire _11393_ ;
wire _5708_ ;
wire _9961_ ;
wire _9541_ ;
wire _9121_ ;
wire _1628_ ;
wire _1208_ ;
wire _5881_ ;
wire _5461_ ;
wire _5041_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _6666_ ;
wire _6246_ ;
wire _1381_ ;
wire _10664_ ;
wire _10244_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _8812_ ;
wire _11869_ ;
wire _11449_ ;
wire _11029_ ;
wire _4732_ ;
wire _4312_ ;
wire _5937_ ;
wire _5517_ ;
wire _11_ ;
wire _9770_ ;
wire _9350_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _5690_ ;
wire _5270_ ;
wire _768_ ;
wire _348_ ;
wire _6895_ ;
wire _6475_ ;
wire _6055_ ;
wire _1190_ ;
wire _10893_ ;
wire _10473_ ;
wire _10053_ ;
wire _2395_ ;
wire _8621_ ;
wire _8201_ ;
wire _11678_ ;
wire _11258_ ;
wire _9826_ ;
wire _9406_ ;
wire _4961_ ;
wire _4541_ ;
wire _4121_ ;
wire _5746_ ;
wire _5326_ ;
wire _1666_ ;
wire areg_17_bF$buf0 ;
wire _1246_ ;
wire areg_17_bF$buf1 ;
wire areg_17_bF$buf2 ;
wire areg_17_bF$buf3 ;
wire areg_17_bF$buf4 ;
wire areg_17_bF$buf5 ;
wire _10949_ ;
wire _10529_ ;
wire _10109_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _3812_ ;
wire _6284_ ;
wire _10282_ ;
wire _7489_ ;
wire _7069_ ;
wire _8850_ ;
wire _8430_ ;
wire _8010_ ;
wire _11487_ ;
wire _11067_ ;
wire _9635_ ;
wire _9215_ ;
wire _4770_ ;
wire _4350_ ;
wire _5975_ ;
wire _5555_ ;
wire _5135_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _7701_ ;
wire _10758_ ;
wire _10338_ ;
wire _386_ ;
wire _8906_ ;
wire _3621_ ;
wire _3201_ ;
wire _6093_ ;
wire _10091_ ;
wire _4826_ ;
wire _4406_ ;
wire _7298_ ;
wire _11296_ ;
wire _9864_ ;
wire _9444_ ;
wire _9024_ ;
wire _5784_ ;
wire _5364_ ;
wire _6989_ ;
wire _6569_ ;
wire _6149_ ;
wire _1284_ ;
wire _7930_ ;
wire _7510_ ;
wire _10987_ ;
wire _10567_ ;
wire _10147_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _8715_ ;
wire _3850_ ;
wire _3430_ ;
wire _3010_ ;
wire _4635_ ;
wire _4215_ ;
wire _9673_ ;
wire _9253_ ;
wire _2701_ ;
wire _5593_ ;
wire _5173_ ;
wire _3906_ ;
wire _6798_ ;
wire _6378_ ;
wire _1093_ ;
wire _10796_ ;
wire _10376_ ;
wire _2298_ ;
wire _8944_ ;
wire _8524_ ;
wire _8104_ ;
wire _9729_ ;
wire _9309_ ;
wire _4864_ ;
wire _4444_ ;
wire _4024_ ;
wire _5649_ ;
wire _5229_ ;
wire _9482_ ;
wire _9062_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2930_ ;
wire _2510_ ;
wire _3715_ ;
wire _6187_ ;
wire _10185_ ;
wire _8753_ ;
wire _8333_ ;
wire _9958_ ;
wire _9538_ ;
wire _9118_ ;
wire _4673_ ;
wire _4253_ ;
wire _5878_ ;
wire _5458_ ;
wire _5038_ ;
wire _9291_ ;
wire _1798_ ;
wire _1378_ ;
wire _7604_ ;
wire _289_ ;
wire _11602_ ;
wire _8809_ ;
wire _3944_ ;
wire _3524_ ;
wire _3104_ ;
wire _5_ ;
wire _4729_ ;
wire _4309_ ;
wire _8982_ ;
wire _8562_ ;
wire _8142_ ;
wire _11199_ ;
wire _9767_ ;
wire _9347_ ;
wire _4482_ ;
wire _4062_ ;
wire _921_ ;
wire _501_ ;
wire _5687_ ;
wire _5267_ ;
wire _1187_ ;
wire _7833_ ;
wire _7413_ ;
wire _11831_ ;
wire _11411_ ;
wire _8618_ ;
wire _3753_ ;
wire _3333_ ;
wire _4958_ ;
wire _4538_ ;
wire _4118_ ;
wire _8791_ ;
wire _8371_ ;
wire _9996_ ;
wire _9576_ ;
wire _9156_ ;
wire _4291_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _5496_ ;
wire _5076_ ;
wire _3809_ ;
wire _7642_ ;
wire _7222_ ;
wire _10699_ ;
wire _10279_ ;
wire _11640_ ;
wire _11220_ ;
wire _8847_ ;
wire _8427_ ;
wire _8007_ ;
wire _3982_ ;
wire _3562_ ;
wire _3142_ ;
wire _4767_ ;
wire _4347_ ;
wire _8180_ ;
wire _46_ ;
wire _6913_ ;
wire _9385_ ;
wire _10911_ ;
wire _2833_ ;
wire _2413_ ;
wire _3618_ ;
wire _7871_ ;
wire _7451_ ;
wire _7031_ ;
wire _10088_ ;
wire _8656_ ;
wire _8236_ ;
wire _3791_ ;
wire _3371_ ;
wire _4996_ ;
wire _4576_ ;
wire _4156_ ;
wire _6722_ ;
wire _6302_ ;
wire _9194_ ;
wire _10720_ ;
wire _10300_ ;
wire _7927_ ;
wire _7507_ ;
wire _2642_ ;
wire _2222_ ;
wire _11505_ ;
wire _3847_ ;
wire _3427_ ;
wire _3007_ ;
wire _7680_ ;
wire _7260_ ;
wire _8885_ ;
wire _8465_ ;
wire _8045_ ;
wire _3180_ ;
wire _1913_ ;
wire _4385_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _6951_ ;
wire _6531_ ;
wire _6111_ ;
wire _7736_ ;
wire _7316_ ;
wire _2871_ ;
wire _2451_ ;
wire _2031_ ;
wire _11734_ ;
wire _11314_ ;
wire _3656_ ;
wire _3236_ ;
wire _5802_ ;
wire _8694_ ;
wire _8274_ ;
wire _1722_ ;
wire _1302_ ;
wire _9899_ ;
wire _9479_ ;
wire _9059_ ;
wire _4194_ ;
wire _633_ ;
wire _213_ ;
wire _2927_ ;
wire _2507_ ;
wire _5399_ ;
wire _6760_ ;
wire _6340_ ;
wire _7965_ ;
wire _7545_ ;
wire _7125_ ;
wire _2680_ ;
wire _2260_ ;
wire _11543_ ;
wire _11123_ ;
wire _3885_ ;
wire _3465_ ;
wire _3045_ ;
wire _5611_ ;
wire _8083_ ;
wire _6816_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _9288_ ;
wire _10814_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _7774_ ;
wire _7354_ ;
wire _11772_ ;
wire _11352_ ;
wire _8979_ ;
wire _8559_ ;
wire _8139_ ;
wire _3694_ ;
wire _3274_ ;
wire _9920_ ;
wire _9500_ ;
wire _4899_ ;
wire _4479_ ;
wire _4059_ ;
wire _5840_ ;
wire _5420_ ;
wire _5000_ ;
wire _918_ ;
wire _6625_ ;
wire _6205_ ;
wire _1760_ ;
wire _1340_ ;
wire _9097_ ;
wire _10623_ ;
wire _10203_ ;
wire _671_ ;
wire _251_ ;
wire _2965_ ;
wire _2545_ ;
wire _2125_ ;
wire _11828_ ;
wire _11408_ ;
wire _7583_ ;
wire _7163_ ;
wire _11581_ ;
wire _11161_ ;
wire _8788_ ;
wire _8368_ ;
wire _3083_ ;
wire _1816_ ;
wire _4288_ ;
wire _727_ ;
wire _307_ ;
wire _6854_ ;
wire _6434_ ;
wire _6014_ ;
wire _10852_ ;
wire _10432_ ;
wire _10012_ ;
wire _480_ ;
wire _7639_ ;
wire _7219_ ;
wire _2774_ ;
wire _2354_ ;
wire _11637_ ;
wire _11217_ ;
wire _3979_ ;
wire _3559_ ;
wire _3139_ ;
wire _4920_ ;
wire _4500_ ;
wire _7392_ ;
wire _11390_ ;
wire _5705_ ;
wire _8597_ ;
wire _8177_ ;
wire _1625_ ;
wire _1205_ ;
wire _4097_ ;
wire _10908_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _6663_ ;
wire _6243_ ;
wire _10661_ ;
wire _10241_ ;
wire _7868_ ;
wire _7448_ ;
wire _7028_ ;
wire _2583_ ;
wire _2163_ ;
wire _11866_ ;
wire _11446_ ;
wire _11026_ ;
wire _3788_ ;
wire _3368_ ;
wire _5934_ ;
wire _5514_ ;
wire breg_10_bF$buf0 ;
wire breg_10_bF$buf1 ;
wire breg_10_bF$buf2 ;
wire breg_10_bF$buf3 ;
wire breg_10_bF$buf4 ;
wire breg_10_bF$buf5 ;
wire _6719_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _10717_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _6892_ ;
wire _6472_ ;
wire _6052_ ;
wire _6582__bF$buf0 ;
wire _6582__bF$buf1 ;
wire _6582__bF$buf2 ;
wire _6582__bF$buf3 ;
wire _10890_ ;
wire _10470_ ;
wire _10050_ ;
wire _7677_ ;
wire _7257_ ;
wire _2392_ ;
wire _11675_ ;
wire _11255_ ;
wire _3597_ ;
wire _3177_ ;
wire _9823_ ;
wire _9403_ ;
wire _5743_ ;
wire _5323_ ;
wire _7100__bF$buf0 ;
wire _7100__bF$buf1 ;
wire _7100__bF$buf2 ;
wire _7100__bF$buf3 ;
wire _6948_ ;
wire _6528_ ;
wire _6108_ ;
wire _1663_ ;
wire _1243_ ;
wire _10946_ ;
wire _10526_ ;
wire _10106_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2868_ ;
wire _2448_ ;
wire _2028_ ;
wire _6281_ ;
wire _7486_ ;
wire _7066_ ;
wire _11484_ ;
wire _11064_ ;
wire _9632_ ;
wire _9212_ ;
wire _1719_ ;
wire _5972_ ;
wire _5552_ ;
wire _5132_ ;
wire _6757_ ;
wire _6337_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _10755_ ;
wire _10335_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _8903_ ;
wire _6090_ ;
wire _4823_ ;
wire _4403_ ;
wire _7295_ ;
wire _11293_ ;
wire _5608_ ;
wire _9861_ ;
wire _9441_ ;
wire _9021_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _5781_ ;
wire _5361_ ;
wire _859_ ;
wire _439_ ;
wire _6986_ ;
wire _6566_ ;
wire _6146_ ;
wire _1281_ ;
wire _10984_ ;
wire _10564_ ;
wire _10144_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _8712_ ;
wire _11769_ ;
wire _11349_ ;
wire _9917_ ;
wire _4632_ ;
wire _4212_ ;
wire _5837_ ;
wire _5417_ ;
wire _9670_ ;
wire _9250_ ;
wire _1757_ ;
wire _1337_ ;
wire _5590_ ;
wire _5170_ ;
wire _668_ ;
wire _248_ ;
wire areg_28_bF$buf0 ;
wire areg_28_bF$buf1 ;
wire areg_28_bF$buf2 ;
wire areg_28_bF$buf3 ;
wire areg_28_bF$buf4 ;
wire _3903_ ;
wire areg_28_bF$buf5 ;
wire _6795_ ;
wire _6375_ ;
wire _1090_ ;
wire _10793_ ;
wire _10373_ ;
wire _2295_ ;
wire _8941_ ;
wire _8521_ ;
wire _8101_ ;
wire _11578_ ;
wire _11158_ ;
wire _9726_ ;
wire _9306_ ;
wire _4861_ ;
wire _4441_ ;
wire _4021_ ;
wire _5646_ ;
wire _5226_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _10849_ ;
wire _10429_ ;
wire _10009_ ;
wire _897_ ;
wire _477_ ;
wire _3712_ ;
wire _6184_ ;
wire _10182_ ;
wire _4917_ ;
wire _7389_ ;
wire _8750_ ;
wire _8330_ ;
wire _11387_ ;
wire _9955_ ;
wire _9535_ ;
wire _9115_ ;
wire _4670_ ;
wire _4250_ ;
wire _5875_ ;
wire _5455_ ;
wire _5035_ ;
wire _1795_ ;
wire _1375_ ;
wire _7601_ ;
wire _10658_ ;
wire _10238_ ;
wire _286_ ;
wire _8806_ ;
wire _3941_ ;
wire _3521_ ;
wire _3101_ ;
wire _2_ ;
wire _4726_ ;
wire _4306_ ;
wire _7198_ ;
wire _11196_ ;
wire _9764_ ;
wire _9344_ ;
wire _5684_ ;
wire _5264_ ;
wire _6889_ ;
wire _6469_ ;
wire _6049_ ;
wire _1184_ ;
wire _7830_ ;
wire _7410_ ;
wire _10887_ ;
wire _10467_ ;
wire _10047_ ;
wire _2389_ ;
wire _8615_ ;
wire _3750_ ;
wire _3330_ ;
wire _4955_ ;
wire _4535_ ;
wire _4115_ ;
wire _9993_ ;
wire _9573_ ;
wire _9153_ ;
wire _2601_ ;
wire _5493_ ;
wire _5073_ ;
wire _3806_ ;
wire _6698_ ;
wire _6278_ ;
wire _10696_ ;
wire _10276_ ;
wire _2198_ ;
wire _8844_ ;
wire _8424_ ;
wire _8004_ ;
wire _9629_ ;
wire _9209_ ;
wire _4764_ ;
wire _4344_ ;
wire _5969_ ;
wire _5549_ ;
wire _5129_ ;
wire _43_ ;
wire _6910_ ;
wire _9382_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2830_ ;
wire _2410_ ;
wire _3615_ ;
wire _6087_ ;
wire _10085_ ;
wire _8653_ ;
wire _8233_ ;
wire _9858_ ;
wire _9438_ ;
wire _9018_ ;
wire _4993_ ;
wire _4573_ ;
wire _4153_ ;
wire _5778_ ;
wire _5358_ ;
wire _9191_ ;
wire _1698_ ;
wire _1278_ ;
wire _7924_ ;
wire _7504_ ;
wire _189_ ;
wire _11502_ ;
wire _8709_ ;
wire _3844_ ;
wire _3424_ ;
wire _3004_ ;
wire _4629_ ;
wire _4209_ ;
wire _8882_ ;
wire _8462_ ;
wire _8042_ ;
wire _11099_ ;
wire _1910_ ;
wire _9667_ ;
wire _9247_ ;
wire _4382_ ;
wire _821_ ;
wire _401_ ;
wire _5587_ ;
wire _5167_ ;
wire _81_ ;
wire _1087_ ;
wire _7733_ ;
wire _7313_ ;
wire _11731_ ;
wire _11311_ ;
wire _8938_ ;
wire _8518_ ;
wire _3653_ ;
wire _3233_ ;
wire areg_12_bF$buf0 ;
wire areg_12_bF$buf1 ;
wire areg_12_bF$buf2 ;
wire areg_12_bF$buf3 ;
wire areg_12_bF$buf4 ;
wire _4858_ ;
wire _4438_ ;
wire _4018_ ;
wire _8691_ ;
wire _8271_ ;
wire _9896_ ;
wire _9476_ ;
wire _9056_ ;
wire _4191_ ;
wire _630_ ;
wire _210_ ;
wire _2924_ ;
wire _2504_ ;
wire _5396_ ;
wire _3709_ ;
wire _7962_ ;
wire _7542_ ;
wire _7122_ ;
wire _10599_ ;
wire _10179_ ;
wire _11540_ ;
wire _11120_ ;
wire _8747_ ;
wire _8327_ ;
wire _3882_ ;
wire _3462_ ;
wire _3042_ ;
wire _4667_ ;
wire _4247_ ;
wire _8080_ ;
wire _6813_ ;
wire _9285_ ;
wire _10811_ ;
wire _2733_ ;
wire _2313_ ;
wire _3938_ ;
wire _3518_ ;
wire _7771_ ;
wire _7351_ ;
wire _8976_ ;
wire _8556_ ;
wire _8136_ ;
wire _3691_ ;
wire _3271_ ;
wire _4896_ ;
wire _4476_ ;
wire _4056_ ;
wire _915_ ;
wire _6622_ ;
wire _6202_ ;
wire _9094_ ;
wire _10620_ ;
wire _10200_ ;
wire _7827_ ;
wire _7407_ ;
wire _2962_ ;
wire _2542_ ;
wire _2122_ ;
wire _11825_ ;
wire _11405_ ;
wire _3747_ ;
wire _3327_ ;
wire _7580_ ;
wire _7160_ ;
wire _8785_ ;
wire _8365_ ;
wire _3080_ ;
wire _1813_ ;
wire _4285_ ;
wire _724_ ;
wire _304_ ;
wire _6851_ ;
wire _6431_ ;
wire _6011_ ;
wire _7636_ ;
wire _7216_ ;
wire _2771_ ;
wire _2351_ ;
wire _11634_ ;
wire _11214_ ;
wire _3976_ ;
wire _3556_ ;
wire _3136_ ;
wire _5702_ ;
wire _8594_ ;
wire _8174_ ;
wire _6907_ ;
wire _1622_ ;
wire _1202_ ;
wire _9799_ ;
wire _9379_ ;
wire _4094_ ;
wire _10905_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2827_ ;
wire _2407_ ;
wire _5299_ ;
wire _6660_ ;
wire _6240_ ;
wire _7865_ ;
wire _7445_ ;
wire _7025_ ;
wire _2580_ ;
wire _2160_ ;
wire _11863_ ;
wire _11443_ ;
wire _11023_ ;
wire _3785_ ;
wire _3365_ ;
wire _5931_ ;
wire _5511_ ;
wire _6716_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _9188_ ;
wire _10714_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _7674_ ;
wire _7254_ ;
wire _11672_ ;
wire _11252_ ;
wire _8879_ ;
wire _8459_ ;
wire _8039_ ;
wire _3594_ ;
wire _3174_ ;
wire _9820_ ;
wire _9400_ ;
wire _1907_ ;
wire _4799_ ;
wire _4379_ ;
wire _5740_ ;
wire _5320_ ;
wire _818_ ;
wire _78_ ;
wire _6945_ ;
wire _6525_ ;
wire _6105_ ;
wire _1660_ ;
wire _1240_ ;
wire _10943_ ;
wire _10523_ ;
wire _10103_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2865_ ;
wire _2445_ ;
wire _2025_ ;
wire _11728_ ;
wire _11308_ ;
wire _7483_ ;
wire _7063_ ;
wire _11481_ ;
wire _11061_ ;
wire _8688_ ;
wire _8268_ ;
wire _1716_ ;
wire _4188_ ;
wire _627_ ;
wire _207_ ;
wire _6754_ ;
wire _6334_ ;
wire _10752_ ;
wire _10332_ ;
wire _380_ ;
wire _7959_ ;
wire _7539_ ;
wire _7119_ ;
wire _2674_ ;
wire _2254_ ;
wire _8900_ ;
wire _11537_ ;
wire _11117_ ;
wire _3879_ ;
wire _3459_ ;
wire _3039_ ;
wire _4820_ ;
wire _4400_ ;
wire _7292_ ;
wire _11290_ ;
wire _5605_ ;
wire _8497_ ;
wire _8077_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _10808_ ;
wire _856_ ;
wire _436_ ;
wire _6983_ ;
wire _6563_ ;
wire _6143_ ;
wire _10981_ ;
wire _10561_ ;
wire _10141_ ;
wire _7768_ ;
wire _7348_ ;
wire _2483_ ;
wire _2063_ ;
wire _11766_ ;
wire _11346_ ;
wire _3688_ ;
wire _3268_ ;
wire _9914_ ;
wire _5834_ ;
wire _5414_ ;
wire _6619_ ;
wire _1754_ ;
wire _1334_ ;
wire _10617_ ;
wire _665_ ;
wire _245_ ;
wire _2959_ ;
wire _2539_ ;
wire _2119_ ;
wire _3900_ ;
wire _6792_ ;
wire _6372_ ;
wire _10790_ ;
wire _10370_ ;
wire _7997_ ;
wire _7577_ ;
wire _7157_ ;
wire _2292_ ;
wire _11575_ ;
wire _11155_ ;
wire _3497_ ;
wire _3077_ ;
wire _9723_ ;
wire _9303_ ;
wire _5643_ ;
wire _5223_ ;
wire _6848_ ;
wire _6428_ ;
wire _6008_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _10846_ ;
wire _10426_ ;
wire _10006_ ;
wire _894_ ;
wire _474_ ;
wire _2768_ ;
wire _2348_ ;
wire _6181_ ;
wire _4914_ ;
wire _7386_ ;
wire _11384_ ;
wire _9952_ ;
wire _9532_ ;
wire _9112_ ;
wire _1619_ ;
wire _5872_ ;
wire _5452_ ;
wire _5032_ ;
wire _6657_ ;
wire _6237_ ;
wire _1792_ ;
wire _1372_ ;
wire _10655_ ;
wire _10235_ ;
wire _283_ ;
wire _2997_ ;
wire _2577_ ;
wire _2157_ ;
wire _8803_ ;
wire _4723_ ;
wire _4303_ ;
wire _7195_ ;
wire _11193_ ;
wire _5928_ ;
wire _5508_ ;
wire _9761_ ;
wire _9341_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _5681_ ;
wire _5261_ ;
wire _759_ ;
wire _339_ ;
wire _6886_ ;
wire _6466_ ;
wire _6046_ ;
wire _1181_ ;
wire _10884_ ;
wire _10464_ ;
wire _10044_ ;
wire _2386_ ;
wire _8612_ ;
wire _11669_ ;
wire _11249_ ;
wire _9817_ ;
wire _4952_ ;
wire _4532_ ;
wire _4112_ ;
wire _5737_ ;
wire _5317_ ;
wire _9990_ ;
wire _9570_ ;
wire _9150_ ;
wire _1657_ ;
wire _1237_ ;
wire _5490_ ;
wire _5070_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _3803_ ;
wire _6695_ ;
wire _6275_ ;
wire _10693_ ;
wire _10273_ ;
wire _2195_ ;
wire _8841_ ;
wire _8421_ ;
wire _8001_ ;
wire _9104__bF$buf0 ;
wire _9104__bF$buf1 ;
wire _11898_ ;
wire _9104__bF$buf2 ;
wire _11478_ ;
wire _9104__bF$buf3 ;
wire _11058_ ;
wire _9626_ ;
wire _9206_ ;
wire _4761_ ;
wire _4341_ ;
wire _5966_ ;
wire _5546_ ;
wire _5126_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _10749_ ;
wire _10329_ ;
wire _797_ ;
wire _377_ ;
wire _3612_ ;
wire _6084_ ;
wire _10082_ ;
wire _4817_ ;
wire _7289_ ;
wire _8650_ ;
wire _8230_ ;
wire _11287_ ;
wire _9855_ ;
wire _9435_ ;
wire _9015_ ;
wire _4990_ ;
wire _4570_ ;
wire _4150_ ;
wire _5775_ ;
wire _5355_ ;
wire _1695_ ;
wire _1275_ ;
wire _7921_ ;
wire _7501_ ;
wire _10978_ ;
wire _10558_ ;
wire _10138_ ;
wire _186_ ;
wire _8706_ ;
wire _3841_ ;
wire _3421_ ;
wire _3001_ ;
wire _4626_ ;
wire _4206_ ;
wire _7098_ ;
wire _11096_ ;
wire _9664_ ;
wire _9244_ ;
wire _5584_ ;
wire _5164_ ;
wire _6789_ ;
wire _6369_ ;
wire _1084_ ;
wire _7730_ ;
wire _7310_ ;
wire _10787_ ;
wire _10367_ ;
wire _2289_ ;
wire _8935_ ;
wire _8515_ ;
wire _3650_ ;
wire _3230_ ;
wire _4855_ ;
wire _4435_ ;
wire _4015_ ;
wire _9893_ ;
wire _9473_ ;
wire _9053_ ;
wire _2921_ ;
wire _2501_ ;
wire _5393_ ;
wire _3706_ ;
wire _6598_ ;
wire _6178_ ;
wire _10596_ ;
wire _10176_ ;
wire _2098_ ;
wire _8744_ ;
wire _8324_ ;
wire _9949_ ;
wire _9529_ ;
wire _9109_ ;
wire _4664_ ;
wire _4244_ ;
wire _5869_ ;
wire _5449_ ;
wire _5029_ ;
wire _6810_ ;
wire _9282_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _3935_ ;
wire _3515_ ;
wire _8973_ ;
wire _8553_ ;
wire _8133_ ;
wire _9758_ ;
wire _9338_ ;
wire _4893_ ;
wire _4473_ ;
wire _4053_ ;
wire _912_ ;
wire _5678_ ;
wire _5258_ ;
wire _9091_ ;
wire _1598_ ;
wire _1178_ ;
wire _7824_ ;
wire _7404_ ;
wire _11822_ ;
wire _11402_ ;
wire _8609_ ;
wire _3744_ ;
wire _3324_ ;
wire _4949_ ;
wire _4529_ ;
wire _4109_ ;
wire _8782_ ;
wire _8362_ ;
wire areg_23_bF$buf0 ;
wire areg_23_bF$buf1 ;
wire areg_23_bF$buf2 ;
wire areg_23_bF$buf3 ;
wire areg_23_bF$buf4 ;
wire _1810_ ;
wire _9987_ ;
wire _9567_ ;
wire _9147_ ;
wire _4282_ ;
wire _721_ ;
wire _301_ ;
wire _5487_ ;
wire _5067_ ;
wire _7633_ ;
wire _7213_ ;
wire _11631_ ;
wire _11211_ ;
wire _8838_ ;
wire _8418_ ;
wire _3973_ ;
wire _3553_ ;
wire _3133_ ;
wire _4758_ ;
wire _4338_ ;
wire _8591_ ;
wire _8171_ ;
wire _37_ ;
wire _6904_ ;
wire _9796_ ;
wire _9376_ ;
wire _4091_ ;
wire _10902_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2824_ ;
wire _2404_ ;
wire _5296_ ;
wire _3609_ ;
wire _7862_ ;
wire _7442_ ;
wire _7022_ ;
wire _10499_ ;
wire _10079_ ;
wire _11860_ ;
wire _11440_ ;
wire _11020_ ;
wire _8647_ ;
wire _8227_ ;
wire _3782_ ;
wire _3362_ ;
wire _4987_ ;
wire _4567_ ;
wire _4147_ ;
wire _6713_ ;
wire _9185_ ;
wire _10711_ ;
wire _7918_ ;
wire _2633_ ;
wire _2213_ ;
wire _3838_ ;
wire _3418_ ;
wire _7671_ ;
wire _7251_ ;
wire _8876_ ;
wire _8456_ ;
wire _8036_ ;
wire _3591_ ;
wire _3171_ ;
wire _1904_ ;
wire _4796_ ;
wire _4376_ ;
wire _815_ ;
wire _75_ ;
wire _6942_ ;
wire _6522_ ;
wire _6102_ ;
wire _10940_ ;
wire _10520_ ;
wire _10100_ ;
wire _7727_ ;
wire _7307_ ;
wire _2862_ ;
wire _2442_ ;
wire _2022_ ;
wire _11725_ ;
wire _11305_ ;
wire _3647_ ;
wire _3227_ ;
wire _7480_ ;
wire _7060_ ;
wire _8685_ ;
wire _8265_ ;
wire _1713_ ;
wire _4185_ ;
wire _624_ ;
wire _204_ ;
wire _2918_ ;
wire areg_5_bF$buf0 ;
wire areg_5_bF$buf1 ;
wire areg_5_bF$buf2 ;
wire areg_5_bF$buf3 ;
wire areg_5_bF$buf4 ;
wire _6751_ ;
wire _6331_ ;
wire _7956_ ;
wire _7536_ ;
wire _7116_ ;
wire _2671_ ;
wire _2251_ ;
wire _11534_ ;
wire _11114_ ;
wire _3876_ ;
wire _3456_ ;
wire _3036_ ;
wire _5420__bF$buf0 ;
wire _5420__bF$buf1 ;
wire _5420__bF$buf2 ;
wire _5420__bF$buf3 ;
wire _5602_ ;
wire _8494_ ;
wire _8074_ ;
wire _6807_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _9699_ ;
wire _9279_ ;
wire _10805_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _5199_ ;
wire _6980_ ;
wire _6560_ ;
wire _6140_ ;
wire _7765_ ;
wire _7345_ ;
wire _2480_ ;
wire _2060_ ;
wire _11763_ ;
wire _11343_ ;
wire _3685_ ;
wire _3265_ ;
wire _9911_ ;
wire _5831_ ;
wire _5411_ ;
wire _909_ ;
wire _6616_ ;
wire _1751_ ;
wire _1331_ ;
wire _9088_ ;
wire _10614_ ;
wire _662_ ;
wire _242_ ;
wire _2956_ ;
wire _2536_ ;
wire _2116_ ;
wire _11819_ ;
wire _7994_ ;
wire _7574_ ;
wire _7154_ ;
wire _11572_ ;
wire _11152_ ;
wire _8779_ ;
wire _8359_ ;
wire _3494_ ;
wire _3074_ ;
wire _9720_ ;
wire _9300_ ;
wire _1807_ ;
wire _4699_ ;
wire _4279_ ;
wire _5640_ ;
wire _5220_ ;
wire _718_ ;
wire _6845_ ;
wire _6425_ ;
wire _6005_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _10843_ ;
wire _10423_ ;
wire _10003_ ;
wire _891_ ;
wire _471_ ;
wire _2765_ ;
wire _2345_ ;
wire _11628_ ;
wire _11208_ ;
wire _4911_ ;
wire _7383_ ;
wire _11381_ ;
wire _8588_ ;
wire _8168_ ;
wire _1616_ ;
wire _4088_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _6654_ ;
wire _6234_ ;
wire _10652_ ;
wire _10232_ ;
wire _280_ ;
wire _7859_ ;
wire _7439_ ;
wire _7019_ ;
wire _2994_ ;
wire _2574_ ;
wire _2154_ ;
wire _8800_ ;
wire _11857_ ;
wire _11437_ ;
wire _11017_ ;
wire _3779_ ;
wire _3359_ ;
wire _4720_ ;
wire _4300_ ;
wire _7192_ ;
wire _11190_ ;
wire _5925_ ;
wire _5505_ ;
wire _8397_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _10708_ ;
wire _756_ ;
wire _336_ ;
wire _6883_ ;
wire _6463_ ;
wire _6043_ ;
wire _10881_ ;
wire _10461_ ;
wire _10041_ ;
wire _7668_ ;
wire _7248_ ;
wire _2383_ ;
wire _11666_ ;
wire _11246_ ;
wire _3588_ ;
wire _3168_ ;
wire _9814_ ;
wire _5734_ ;
wire _5314_ ;
wire _6939_ ;
wire _6519_ ;
wire _1654_ ;
wire _1234_ ;
wire _10937_ ;
wire _10517_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2859_ ;
wire _2439_ ;
wire _2019_ ;
wire _3800_ ;
wire _6692_ ;
wire _6272_ ;
wire _10690_ ;
wire _10270_ ;
wire _7897_ ;
wire _7477_ ;
wire _7057_ ;
wire _2192_ ;
wire _11895_ ;
wire _11475_ ;
wire _11055_ ;
wire _3397_ ;
wire _9623_ ;
wire _9203_ ;
wire _5963_ ;
wire _5543_ ;
wire _5123_ ;
wire _6748_ ;
wire _6328_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _10746_ ;
wire _10326_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _6081_ ;
wire _4814_ ;
wire _7286_ ;
wire _11284_ ;
wire _9852_ ;
wire _9432_ ;
wire _9012_ ;
wire _1939_ ;
wire _1519_ ;
wire _5772_ ;
wire _5352_ ;
wire _6977_ ;
wire _6557_ ;
wire _6137_ ;
wire _1692_ ;
wire _1272_ ;
wire _10975_ ;
wire _10555_ ;
wire _10135_ ;
wire _183_ ;
wire _2897_ ;
wire _2477_ ;
wire _2057_ ;
wire _8703_ ;
wire _9908_ ;
wire _4623_ ;
wire _4203_ ;
wire _7095_ ;
wire _11093_ ;
wire _5828_ ;
wire _5408_ ;
wire _9661_ ;
wire _9241_ ;
wire _1748_ ;
wire _1328_ ;
wire _5581_ ;
wire _5161_ ;
wire _659_ ;
wire _239_ ;
wire _6786_ ;
wire _6366_ ;
wire _1081_ ;
wire _10784_ ;
wire _10364_ ;
wire _2286_ ;
wire _8932_ ;
wire _8512_ ;
wire _11569_ ;
wire _11149_ ;
wire _9717_ ;
wire _4852_ ;
wire _4432_ ;
wire _4012_ ;
wire _5637_ ;
wire _5217_ ;
wire _9890_ ;
wire _9470_ ;
wire _9050_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _5390_ ;
wire _888_ ;
wire _468_ ;
wire _3703_ ;
wire _6595_ ;
wire _6175_ ;
wire _10593_ ;
wire _10173_ ;
wire _4908_ ;
wire _2095_ ;
wire _8741_ ;
wire _8321_ ;
wire _11798_ ;
wire _11378_ ;
wire _9946_ ;
wire _9526_ ;
wire _9106_ ;
wire _4661_ ;
wire _4241_ ;
wire _5866_ ;
wire _5446_ ;
wire _5026_ ;
wire _1786_ ;
wire _1366_ ;
wire _10649_ ;
wire _10229_ ;
wire _697_ ;
wire _277_ ;
wire _3932_ ;
wire _3512_ ;
wire _4717_ ;
wire _7189_ ;
wire _8970_ ;
wire _8550_ ;
wire _8130_ ;
wire _11187_ ;
wire breg_25_bF$buf0 ;
wire breg_25_bF$buf1 ;
wire breg_25_bF$buf2 ;
wire breg_25_bF$buf3 ;
wire breg_25_bF$buf4 ;
wire breg_25_bF$buf5 ;
wire _9755_ ;
wire _9335_ ;
wire _4890_ ;
wire _4470_ ;
wire _4050_ ;
wire _5675_ ;
wire _5255_ ;
wire _1595_ ;
wire _1175_ ;
wire _7821_ ;
wire _7401_ ;
wire _10878_ ;
wire _10458_ ;
wire _10038_ ;
wire breg_3_bF$buf0 ;
wire breg_3_bF$buf1 ;
wire breg_3_bF$buf2 ;
wire breg_3_bF$buf3 ;
wire breg_3_bF$buf4 ;
wire breg_3_bF$buf5 ;
wire _8606_ ;
wire _3741_ ;
wire _3321_ ;
wire _4946_ ;
wire _4526_ ;
wire _4106_ ;
wire _9984_ ;
wire _9564_ ;
wire _9144_ ;
wire _5484_ ;
wire _5064_ ;
wire _6689_ ;
wire _6269_ ;
wire _7630_ ;
wire _7210_ ;
wire _10687_ ;
wire _10267_ ;
wire _2189_ ;
wire _8835_ ;
wire _8415_ ;
wire _3970_ ;
wire _3550_ ;
wire _3130_ ;
wire _4755_ ;
wire _4335_ ;
wire _34_ ;
wire _6901_ ;
wire _9793_ ;
wire _9373_ ;
wire _2821_ ;
wire _2401_ ;
wire _5293_ ;
wire _3606_ ;
wire _6498_ ;
wire _6078_ ;
wire _10496_ ;
wire _10076_ ;
wire _8644_ ;
wire _8224_ ;
wire _9849_ ;
wire _9429_ ;
wire _9009_ ;
wire _4984_ ;
wire _4564_ ;
wire _4144_ ;
wire _5769_ ;
wire _5349_ ;
wire _6710_ ;
wire _9182_ ;
wire _1689_ ;
wire _1269_ ;
wire _7915_ ;
wire _2630_ ;
wire _2210_ ;
wire _3835_ ;
wire _3415_ ;
wire _8873_ ;
wire _8453_ ;
wire _8033_ ;
wire _1901_ ;
wire _9658_ ;
wire _9238_ ;
wire _4793_ ;
wire _4373_ ;
wire _812_ ;
wire _5998_ ;
wire _5578_ ;
wire _5158_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _7724_ ;
wire _7304_ ;
wire _11722_ ;
wire _11302_ ;
wire _8929_ ;
wire _8509_ ;
wire _3644_ ;
wire _3224_ ;
wire _4849_ ;
wire _4429_ ;
wire _4009_ ;
wire _8682_ ;
wire _8262_ ;
wire _1710_ ;
wire _9887_ ;
wire _9467_ ;
wire _9047_ ;
wire _4182_ ;
wire _621_ ;
wire _201_ ;
wire _2915_ ;
wire _5387_ ;
wire _7953_ ;
wire _7533_ ;
wire _7113_ ;
wire _11531_ ;
wire _11111_ ;
wire _8738_ ;
wire _8318_ ;
wire _3873_ ;
wire _3453_ ;
wire _3033_ ;
wire _4658_ ;
wire _4238_ ;
wire _8491_ ;
wire _8071_ ;
wire _6804_ ;
wire _9696_ ;
wire _9276_ ;
wire _10802_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _5196_ ;
wire _3929_ ;
wire _3509_ ;
wire _7762_ ;
wire _7342_ ;
wire _10399_ ;
wire _11760_ ;
wire _11340_ ;
wire _8967_ ;
wire _8547_ ;
wire _8127_ ;
wire _3682_ ;
wire _3262_ ;
wire _4887_ ;
wire _4467_ ;
wire _4047_ ;
wire _906_ ;
wire _6613_ ;
wire _9085_ ;
wire _10611_ ;
wire _7818_ ;
wire _2953_ ;
wire _2533_ ;
wire _2113_ ;
wire _11816_ ;
wire _3738_ ;
wire _3318_ ;
wire _7991_ ;
wire _7571_ ;
wire _7151_ ;
wire _8776_ ;
wire _8356_ ;
wire _3491_ ;
wire _3071_ ;
wire _1804_ ;
wire _4696_ ;
wire _4276_ ;
wire _715_ ;
wire _6842_ ;
wire _6422_ ;
wire _6002_ ;
wire _10840_ ;
wire _10420_ ;
wire _10000_ ;
wire _7627_ ;
wire _7207_ ;
wire _2762_ ;
wire _2342_ ;
wire _11625_ ;
wire _11205_ ;
wire _3967_ ;
wire _3547_ ;
wire _3127_ ;
wire _7380_ ;
wire _8585_ ;
wire _8165_ ;
wire _1613_ ;
wire _4085_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2818_ ;
wire _6651_ ;
wire _6231_ ;
wire _7856_ ;
wire _7436_ ;
wire _7016_ ;
wire _2991_ ;
wire _2571_ ;
wire _2151_ ;
wire _11854_ ;
wire _11434_ ;
wire _11014_ ;
wire _3776_ ;
wire _3356_ ;
wire _5922_ ;
wire _5502_ ;
wire _8394_ ;
wire _6707_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _9599_ ;
wire _9179_ ;
wire _10705_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _5099_ ;
wire _6880_ ;
wire _6460_ ;
wire _6040_ ;
wire _7665_ ;
wire _7245_ ;
wire _2380_ ;
wire _11663_ ;
wire _11243_ ;
wire _3585_ ;
wire _3165_ ;
wire _9811_ ;
wire _5731_ ;
wire _5311_ ;
wire _809_ ;
wire _69_ ;
wire _6936_ ;
wire _6516_ ;
wire _1651_ ;
wire _1231_ ;
wire _10934_ ;
wire _10514_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2856_ ;
wire _2436_ ;
wire _2016_ ;
wire _11719_ ;
wire _7894_ ;
wire _7474_ ;
wire _7054_ ;
wire _11892_ ;
wire _11472_ ;
wire _11052_ ;
wire _8679_ ;
wire _8259_ ;
wire _3394_ ;
wire _9620_ ;
wire _9200_ ;
wire _1707_ ;
wire _4599_ ;
wire _4179_ ;
wire _5960_ ;
wire _5540_ ;
wire _5120_ ;
wire _618_ ;
wire _6745_ ;
wire _6325_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _10743_ ;
wire _10323_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _11528_ ;
wire _11108_ ;
wire _4811_ ;
wire _7283_ ;
wire _11281_ ;
wire _8488_ ;
wire _8068_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _6974_ ;
wire _6554_ ;
wire _6134_ ;
wire _10972_ ;
wire _10552_ ;
wire _10132_ ;
wire _180_ ;
wire _7759_ ;
wire _7339_ ;
wire _2894_ ;
wire _2474_ ;
wire _2054_ ;
wire _8700_ ;
wire _11757_ ;
wire _11337_ ;
wire _3679_ ;
wire _3259_ ;
wire _9905_ ;
wire _4620_ ;
wire _4200_ ;
wire _7092_ ;
wire _11090_ ;
wire _5825_ ;
wire _5405_ ;
wire _8297_ ;
wire _1745_ ;
wire _1325_ ;
wire _10608_ ;
wire _656_ ;
wire _236_ ;
wire _6783_ ;
wire _6363_ ;
wire _10781_ ;
wire _10361_ ;
wire _7988_ ;
wire _7568_ ;
wire _7148_ ;
wire _2283_ ;
wire _11566_ ;
wire _11146_ ;
wire _3488_ ;
wire _3068_ ;
wire _9714_ ;
wire _5634_ ;
wire _5214_ ;
wire _6839_ ;
wire _6419_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _10837_ ;
wire _10417_ ;
wire _885_ ;
wire _465_ ;
wire _2759_ ;
wire _2339_ ;
wire _3700_ ;
wire _6592_ ;
wire _6172_ ;
wire _10590_ ;
wire _10170_ ;
wire _4905_ ;
wire _7797_ ;
wire _7377_ ;
wire _2092_ ;
wire _11795_ ;
wire _11375_ ;
wire _3297_ ;
wire _9943_ ;
wire _9523_ ;
wire _9103_ ;
wire _5863_ ;
wire _5443_ ;
wire _5023_ ;
wire _6648_ ;
wire _6228_ ;
wire _1783_ ;
wire _1363_ ;
wire _10646_ ;
wire _10226_ ;
wire _694_ ;
wire _274_ ;
wire _2988_ ;
wire _2568_ ;
wire _2148_ ;
wire _4714_ ;
wire _7186_ ;
wire _11184_ ;
wire _5919_ ;
wire _9752_ ;
wire _9332_ ;
wire _1839_ ;
wire _1419_ ;
wire _5672_ ;
wire _5252_ ;
wire _6877_ ;
wire _6457_ ;
wire _6037_ ;
wire _1592_ ;
wire _1172_ ;
wire _10875_ ;
wire _10455_ ;
wire _10035_ ;
wire _2797_ ;
wire _2377_ ;
wire _549__bF$buf0 ;
wire _549__bF$buf1 ;
wire _549__bF$buf2 ;
wire _549__bF$buf3 ;
wire _549__bF$buf4 ;
wire _8603_ ;
wire _9808_ ;
wire _4943_ ;
wire _4523_ ;
wire _4103_ ;
wire _5728_ ;
wire _5308_ ;
wire _9981_ ;
wire _9561_ ;
wire _9141_ ;
wire _1648_ ;
wire _1228_ ;
wire _5481_ ;
wire _5061_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _6686_ ;
wire _6266_ ;
wire _10684_ ;
wire _10264_ ;
wire _2186_ ;
wire _8832_ ;
wire _8412_ ;
wire _11889_ ;
wire _11469_ ;
wire _11049_ ;
wire _9617_ ;
wire _4752_ ;
wire _4332_ ;
wire _5957_ ;
wire _5537_ ;
wire _5117_ ;
wire _31_ ;
wire _9790_ ;
wire _9370_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _5290_ ;
wire _788_ ;
wire _368_ ;
wire _3603_ ;
wire _6495_ ;
wire _6075_ ;
wire _10493_ ;
wire _10073_ ;
wire _4808_ ;
wire _8641_ ;
wire _8221_ ;
wire _11698_ ;
wire _11278_ ;
wire breg_17_bF$buf0 ;
wire breg_17_bF$buf1 ;
wire breg_17_bF$buf2 ;
wire breg_17_bF$buf3 ;
wire breg_17_bF$buf4 ;
wire _9846_ ;
wire _9426_ ;
wire _9006_ ;
wire _4981_ ;
wire _4561_ ;
wire _4141_ ;
wire _5766_ ;
wire _5346_ ;
wire _1686_ ;
wire _1266_ ;
wire _7912_ ;
wire _10969_ ;
wire _10549_ ;
wire _10129_ ;
wire _597_ ;
wire _177_ ;
wire _3832_ ;
wire _3412_ ;
wire _4617_ ;
wire _7089_ ;
wire _8870_ ;
wire _8450_ ;
wire _8030_ ;
wire _11087_ ;
wire _9655_ ;
wire _9235_ ;
wire _4790_ ;
wire _4370_ ;
wire _5995_ ;
wire _5575_ ;
wire _5155_ ;
wire _1495_ ;
wire _1075_ ;
wire _7721_ ;
wire _7301_ ;
wire _10778_ ;
wire _10358_ ;
wire _8926_ ;
wire _8506_ ;
wire _3641_ ;
wire _3221_ ;
wire _4846_ ;
wire _4426_ ;
wire _4006_ ;
wire _9884_ ;
wire _9464_ ;
wire _9044_ ;
wire _2912_ ;
wire _5384_ ;
wire _6589_ ;
wire _6169_ ;
wire _7950_ ;
wire _7530_ ;
wire _7110_ ;
wire _10587_ ;
wire _10167_ ;
wire _2089_ ;
wire _8735_ ;
wire _8315_ ;
wire _3870_ ;
wire _3450_ ;
wire _3030_ ;
wire _4655_ ;
wire _4235_ ;
wire _6801_ ;
wire _9693_ ;
wire _9273_ ;
wire _2721_ ;
wire _2301_ ;
wire _5193_ ;
wire _3926_ ;
wire _3506_ ;
wire _6398_ ;
wire _2560__bF$buf0 ;
wire _2560__bF$buf1 ;
wire _10396_ ;
wire _2560__bF$buf2 ;
wire _2560__bF$buf3 ;
wire _2560__bF$buf4 ;
wire _8964_ ;
wire _8544_ ;
wire _8124_ ;
wire _9749_ ;
wire _9329_ ;
wire _4884_ ;
wire _4464_ ;
wire _4044_ ;
wire _903_ ;
wire _5669_ ;
wire _5249_ ;
wire _6610_ ;
wire _9082_ ;
wire _1589_ ;
wire _1169_ ;
wire _7815_ ;
wire _2950_ ;
wire _2530_ ;
wire _2110_ ;
wire _11813_ ;
wire _3735_ ;
wire _3315_ ;
wire _8773_ ;
wire _8353_ ;
wire _1801_ ;
wire _9978_ ;
wire _9558_ ;
wire _9138_ ;
wire _4693_ ;
wire _4273_ ;
wire _712_ ;
wire _5898_ ;
wire _5478_ ;
wire _5058_ ;
wire _1398_ ;
wire _7624_ ;
wire _7204_ ;
wire _11622_ ;
wire _11202_ ;
wire _8829_ ;
wire _8409_ ;
wire _3964_ ;
wire _3544_ ;
wire _3124_ ;
wire _4749_ ;
wire _4329_ ;
wire _8582_ ;
wire _8162_ ;
wire _28_ ;
wire _1610_ ;
wire _9787_ ;
wire _9367_ ;
wire _4082_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _2815_ ;
wire _5287_ ;
wire _7853_ ;
wire _7433_ ;
wire _7013_ ;
wire _11851_ ;
wire _11431_ ;
wire _11011_ ;
wire _8638_ ;
wire _8218_ ;
wire _3773_ ;
wire _3353_ ;
wire _4978_ ;
wire _4558_ ;
wire _4138_ ;
wire _8391_ ;
wire _6704_ ;
wire _9596_ ;
wire _9176_ ;
wire _10702_ ;
wire _750_ ;
wire _330_ ;
wire _7909_ ;
wire _2624_ ;
wire _2204_ ;
wire _5096_ ;
wire breg_20_bF$buf0 ;
wire _11907_ ;
wire breg_20_bF$buf1 ;
wire breg_20_bF$buf2 ;
wire breg_20_bF$buf3 ;
wire breg_20_bF$buf4 ;
wire _3829_ ;
wire _3409_ ;
wire _7662_ ;
wire _7242_ ;
wire _10299_ ;
wire _11660_ ;
wire _11240_ ;
wire _8867_ ;
wire _8447_ ;
wire _8027_ ;
wire _3582_ ;
wire _3162_ ;
wire _4787_ ;
wire _4367_ ;
wire _806_ ;
wire _66_ ;
wire _6933_ ;
wire _6513_ ;
wire _10931_ ;
wire _10511_ ;
wire _7718_ ;
wire _2853_ ;
wire _2433_ ;
wire _2013_ ;
wire _11716_ ;
wire _3638_ ;
wire _3218_ ;
wire _7891_ ;
wire _7471_ ;
wire _7051_ ;
wire _8676_ ;
wire _8256_ ;
wire _3391_ ;
wire _1704_ ;
wire _4596_ ;
wire _4176_ ;
wire _615_ ;
wire _2909_ ;
wire _6742_ ;
wire _6322_ ;
wire _10740_ ;
wire _10320_ ;
wire _7947_ ;
wire _7527_ ;
wire _7107_ ;
wire _2662_ ;
wire _2242_ ;
wire _11525_ ;
wire _11105_ ;
wire _3867_ ;
wire _3447_ ;
wire _3027_ ;
wire _7280_ ;
wire _8485_ ;
wire _8065_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _6971_ ;
wire _6551_ ;
wire _6131_ ;
wire _7756_ ;
wire _7336_ ;
wire _2891_ ;
wire _2471_ ;
wire _2051_ ;
wire _11754_ ;
wire _11334_ ;
wire _3676_ ;
wire _3256_ ;
wire _9902_ ;
wire _5822_ ;
wire _5402_ ;
wire _8294_ ;
wire _6607_ ;
wire _1742_ ;
wire _1322_ ;
wire _9499_ ;
wire _9079_ ;
wire _10605_ ;
wire _653_ ;
wire _233_ ;
wire _2947_ ;
wire _2527_ ;
wire _2107_ ;
wire _6780_ ;
wire _6360_ ;
wire _7985_ ;
wire _7565_ ;
wire _7145_ ;
wire areg_19_bF$buf0 ;
wire areg_19_bF$buf1 ;
wire _2280_ ;
wire areg_19_bF$buf2 ;
wire areg_19_bF$buf3 ;
wire areg_19_bF$buf4 ;
wire areg_19_bF$buf5 ;
wire _11563_ ;
wire _11143_ ;
wire _3485_ ;
wire _3065_ ;
wire _9711_ ;
wire _5631_ ;
wire _5211_ ;
wire _709_ ;
wire _6836_ ;
wire _6416_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _10834_ ;
wire _10414_ ;
wire _882_ ;
wire _462_ ;
wire _2756_ ;
wire _2336_ ;
wire _11619_ ;
wire _4902_ ;
wire _7794_ ;
wire _7374_ ;
wire _11792_ ;
wire _11372_ ;
wire _8999_ ;
wire _8579_ ;
wire _8159_ ;
wire _3294_ ;
wire _9940_ ;
wire _9520_ ;
wire _9100_ ;
wire _1607_ ;
wire _4499_ ;
wire _4079_ ;
wire _5860_ ;
wire _5440_ ;
wire _5020_ ;
wire _938_ ;
wire _518_ ;
wire _6645_ ;
wire _6225_ ;
wire _1780_ ;
wire _1360_ ;
wire _10643_ ;
wire _10223_ ;
wire _691_ ;
wire _271_ ;
wire _2985_ ;
wire _2565_ ;
wire _2145_ ;
wire _11848_ ;
wire _11428_ ;
wire _11008_ ;
wire _4711_ ;
wire _7183_ ;
wire _11181_ ;
wire _5916_ ;
wire _8388_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _6874_ ;
wire _6454_ ;
wire _6034_ ;
wire _10872_ ;
wire _10452_ ;
wire _10032_ ;
wire _7659_ ;
wire _7239_ ;
wire _2794_ ;
wire _2374_ ;
wire _8600_ ;
wire _11657_ ;
wire _11237_ ;
wire _3999_ ;
wire _3579_ ;
wire _3159_ ;
wire _9805_ ;
wire _4940_ ;
wire _4520_ ;
wire _4100_ ;
wire _5725_ ;
wire _5305_ ;
wire _8197_ ;
wire _1645_ ;
wire _1225_ ;
wire _10928_ ;
wire _10508_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _6683_ ;
wire _6263_ ;
wire _10681_ ;
wire _10261_ ;
wire _7888_ ;
wire _7468_ ;
wire _7048_ ;
wire _2183_ ;
wire _11886_ ;
wire _11466_ ;
wire _11046_ ;
wire _3388_ ;
wire _9614_ ;
wire _5954_ ;
wire _5534_ ;
wire _5114_ ;
wire _6739_ ;
wire _6319_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _10737_ ;
wire _10317_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _3600_ ;
wire _6492_ ;
wire _6072_ ;
wire _10490_ ;
wire _10070_ ;
wire _4805_ ;
wire _7697_ ;
wire _7277_ ;
wire _11695_ ;
wire _11275_ ;
wire _3197_ ;
wire _9843_ ;
wire _9423_ ;
wire _9003_ ;
wire _5763_ ;
wire _5343_ ;
wire _6968_ ;
wire _6548_ ;
wire _6128_ ;
wire _1683_ ;
wire _1263_ ;
wire _10966_ ;
wire _10546_ ;
wire _10126_ ;
wire _594_ ;
wire _174_ ;
wire _2888_ ;
wire _2468_ ;
wire _2048_ ;
wire _4614_ ;
wire _7086_ ;
wire _11084_ ;
wire _5819_ ;
wire _9652_ ;
wire _9232_ ;
wire _1739_ ;
wire _1319_ ;
wire _5992_ ;
wire _5572_ ;
wire _5152_ ;
wire _6777_ ;
wire _6357_ ;
wire _1492_ ;
wire _1072_ ;
wire _7711__bF$buf0 ;
wire _7711__bF$buf1 ;
wire _7711__bF$buf2 ;
wire _7711__bF$buf3 ;
wire _10775_ ;
wire _10355_ ;
wire _2697_ ;
wire _2277_ ;
wire _8923_ ;
wire _8503_ ;
wire _9708_ ;
wire _4843_ ;
wire _4423_ ;
wire _4003_ ;
wire _5628_ ;
wire _5208_ ;
wire _9881_ ;
wire _9461_ ;
wire _9041_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _5381_ ;
wire _879_ ;
wire _459_ ;
wire _6586_ ;
wire _6166_ ;
wire _10584_ ;
wire _10164_ ;
wire _2086_ ;
wire _8732_ ;
wire _8312_ ;
wire _11789_ ;
wire _11369_ ;
wire _9937_ ;
wire _9517_ ;
wire _4652_ ;
wire _4232_ ;
wire _5857_ ;
wire _5437_ ;
wire _5017_ ;
wire _9690_ ;
wire _9270_ ;
wire _1777_ ;
wire _1357_ ;
wire _5190_ ;
wire _688_ ;
wire _268_ ;
wire _3923_ ;
wire _3503_ ;
wire _6395_ ;
wire _10393_ ;
wire _4708_ ;
wire _8961_ ;
wire _8541_ ;
wire _8121_ ;
wire _11598_ ;
wire _11178_ ;
wire _9746_ ;
wire _9326_ ;
wire _4881_ ;
wire _4461_ ;
wire _4041_ ;
wire _900_ ;
wire _5666_ ;
wire _5246_ ;
wire _1586_ ;
wire _1166_ ;
wire _7812_ ;
wire _10869_ ;
wire _10449_ ;
wire _10029_ ;
wire _497_ ;
wire _11810_ ;
wire _3732_ ;
wire _3312_ ;
wire _4937_ ;
wire _4517_ ;
wire _8770_ ;
wire _8350_ ;
wire _9975_ ;
wire _9555_ ;
wire _9135_ ;
wire _4690_ ;
wire _4270_ ;
wire _5895_ ;
wire _5475_ ;
wire _5055_ ;
wire _1395_ ;
wire _7621_ ;
wire _7201_ ;
wire _10678_ ;
wire _10258_ ;
wire _8826_ ;
wire _8406_ ;
wire _3961_ ;
wire _3541_ ;
wire _3121_ ;
wire _2465__bF$buf0 ;
wire _2465__bF$buf1 ;
wire _2465__bF$buf2 ;
wire _2465__bF$buf3 ;
wire _2465__bF$buf4 ;
wire _4746_ ;
wire _4326_ ;
wire _25_ ;
wire _9784_ ;
wire _9364_ ;
wire _2812_ ;
wire _5284_ ;
wire _6489_ ;
wire _6069_ ;
wire _7850_ ;
wire _7430_ ;
wire _7010_ ;
wire _10487_ ;
wire _10067_ ;
wire _8635_ ;
wire _8215_ ;
wire _3770_ ;
wire _3350_ ;
wire _4975_ ;
wire _4555_ ;
wire _4135_ ;
wire _6701_ ;
wire _9593_ ;
wire _9173_ ;
wire _7906_ ;
wire _2621_ ;
wire _2201_ ;
wire _5093_ ;
wire _11904_ ;
wire _3826_ ;
wire _3406_ ;
wire _6298_ ;
wire _10296_ ;
wire _8864_ ;
wire _8444_ ;
wire _8024_ ;
wire _9649_ ;
wire _9229_ ;
wire _4784_ ;
wire _4364_ ;
wire _803_ ;
wire _5989_ ;
wire _5569_ ;
wire _5149_ ;
wire _63_ ;
wire _6930_ ;
wire _6510_ ;
wire _1489_ ;
wire _1069_ ;
wire _7715_ ;
wire _2850_ ;
wire _2430_ ;
wire _2010_ ;
wire _11713_ ;
wire _3635_ ;
wire _3215_ ;
wire _8673_ ;
wire _8253_ ;
wire _1701_ ;
wire _9878_ ;
wire _9458_ ;
wire _9038_ ;
wire _4593_ ;
wire _4173_ ;
wire _612_ ;
wire _2906_ ;
wire _5798_ ;
wire _5378_ ;
wire _1298_ ;
wire _7944_ ;
wire _7524_ ;
wire _7104_ ;
wire _11522_ ;
wire _11102_ ;
wire _10869__bF$buf0 ;
wire _8729_ ;
wire _10869__bF$buf1 ;
wire _8309_ ;
wire _10869__bF$buf2 ;
wire _10869__bF$buf3 ;
wire _3864_ ;
wire _3444_ ;
wire _3024_ ;
wire _4649_ ;
wire _4229_ ;
wire _8482_ ;
wire _8062_ ;
wire _1930_ ;
wire _1510_ ;
wire _9687_ ;
wire _9267_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _5187_ ;
wire breg_12_bF$buf0 ;
wire breg_12_bF$buf1 ;
wire breg_12_bF$buf2 ;
wire breg_12_bF$buf3 ;
wire breg_12_bF$buf4 ;
wire _7753_ ;
wire _7333_ ;
wire _11751_ ;
wire _11331_ ;
wire _8958_ ;
wire _8538_ ;
wire _8118_ ;
wire _3673_ ;
wire _3253_ ;
wire _4878_ ;
wire _4458_ ;
wire _4038_ ;
wire _8291_ ;
wire _6604_ ;
wire _9496_ ;
wire _9076_ ;
wire _10602_ ;
wire _650_ ;
wire _230_ ;
wire _7809_ ;
wire _2944_ ;
wire _2524_ ;
wire _2104_ ;
wire _11807_ ;
wire _3729_ ;
wire _3309_ ;
wire _7982_ ;
wire _7562_ ;
wire _7142_ ;
wire _10199_ ;
wire _11560_ ;
wire _11140_ ;
wire _8767_ ;
wire _8347_ ;
wire _3482_ ;
wire _3062_ ;
wire _4687_ ;
wire _4267_ ;
wire _706_ ;
wire _6833_ ;
wire _6413_ ;
wire _10831_ ;
wire _10411_ ;
wire _7618_ ;
wire _2753_ ;
wire _2333_ ;
wire _11616_ ;
wire _3958_ ;
wire _3538_ ;
wire _3118_ ;
wire _7791_ ;
wire _7371_ ;
wire _8996_ ;
wire _8576_ ;
wire _8156_ ;
wire _3291_ ;
wire _1604_ ;
wire _4496_ ;
wire _4076_ ;
wire _935_ ;
wire _515_ ;
wire _2809_ ;
wire _6642_ ;
wire _6222_ ;
wire _10640_ ;
wire _10220_ ;
wire _7847_ ;
wire _7427_ ;
wire _7007_ ;
wire _2982_ ;
wire _2562_ ;
wire _2142_ ;
wire _11845_ ;
wire _11425_ ;
wire _11005_ ;
wire _3767_ ;
wire _3347_ ;
wire _7180_ ;
wire _5913_ ;
wire _8385_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _6871_ ;
wire _6451_ ;
wire _6031_ ;
wire _7656_ ;
wire _7236_ ;
wire _2791_ ;
wire _2371_ ;
wire _11654_ ;
wire _11234_ ;
wire _3996_ ;
wire _3576_ ;
wire _3156_ ;
wire _9802_ ;
wire _5722_ ;
wire _5302_ ;
wire _8194_ ;
wire _6927_ ;
wire _6507_ ;
wire _1642_ ;
wire _1222_ ;
wire _9399_ ;
wire _10925_ ;
wire _10505_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2847_ ;
wire _2427_ ;
wire _2007_ ;
wire _6680_ ;
wire _6260_ ;
wire _7885_ ;
wire _7465_ ;
wire _7045_ ;
wire _2180_ ;
wire _11883_ ;
wire _11463_ ;
wire _11043_ ;
wire _3385_ ;
wire _9611_ ;
wire _5951_ ;
wire _5531_ ;
wire _5111_ ;
wire _609_ ;
wire _6736_ ;
wire _6316_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire _10734_ ;
wire _10314_ ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _11519_ ;
wire _4802_ ;
wire _7694_ ;
wire _7274_ ;
wire _11692_ ;
wire _11272_ ;
wire _8899_ ;
wire _8479_ ;
wire _8059_ ;
wire _3194_ ;
wire _9840_ ;
wire _9420_ ;
wire _9000_ ;
wire _1927_ ;
wire _1507_ ;
wire _4399_ ;
wire _5760_ ;
wire _5340_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _6965_ ;
wire _6545_ ;
wire _6125_ ;
wire _1680_ ;
wire _1260_ ;
wire _10963_ ;
wire _10543_ ;
wire _10123_ ;
wire _591_ ;
wire _171_ ;
wire _2885_ ;
wire _2465_ ;
wire _2045_ ;
wire _11748_ ;
wire _11328_ ;
wire _4611_ ;
wire _7083_ ;
wire _11081_ ;
wire _5816_ ;
wire _8288_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _6774_ ;
wire _6354_ ;
wire _10772_ ;
wire _10352_ ;
wire _7979_ ;
wire _7559_ ;
wire _7139_ ;
wire _2694_ ;
wire _2274_ ;
wire _8920_ ;
wire _8500_ ;
wire _11557_ ;
wire _11137_ ;
wire _3899_ ;
wire _3479_ ;
wire _3059_ ;
wire _9705_ ;
wire _4840_ ;
wire _4420_ ;
wire _4000_ ;
wire _5625_ ;
wire _5205_ ;
wire _8097_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _10828_ ;
wire _10408_ ;
wire _876_ ;
wire _456_ ;
wire _6583_ ;
wire _6163_ ;
wire _10581_ ;
wire _10161_ ;
wire _7788_ ;
wire _7368_ ;
wire _2083_ ;
wire _11786_ ;
wire _11366_ ;
wire _3288_ ;
wire _9934_ ;
wire _9514_ ;
wire _5854_ ;
wire _5434_ ;
wire _5014_ ;
wire _6639_ ;
wire _6219_ ;
wire _1774_ ;
wire _1354_ ;
wire _10637_ ;
wire _10217_ ;
wire _2551__bF$buf0 ;
wire _2551__bF$buf1 ;
wire _2551__bF$buf2 ;
wire _2551__bF$buf3 ;
wire _685_ ;
wire _265_ ;
wire _2979_ ;
wire _2559_ ;
wire _2139_ ;
wire _3920_ ;
wire _3500_ ;
wire _6392_ ;
wire _10390_ ;
wire _4705_ ;
wire _7597_ ;
wire _7177_ ;
wire _11595_ ;
wire _11175_ ;
wire _3097_ ;
wire _9743_ ;
wire _9323_ ;
wire _5663_ ;
wire _5243_ ;
wire _6868_ ;
wire _6448_ ;
wire _6028_ ;
wire _1583_ ;
wire _1163_ ;
wire _10866_ ;
wire _10446_ ;
wire _10026_ ;
wire _494_ ;
wire _2788_ ;
wire _2368_ ;
wire _4934_ ;
wire _4514_ ;
wire _5719_ ;
wire _9972_ ;
wire _9552_ ;
wire _9132_ ;
wire _1639_ ;
wire _1219_ ;
wire areg_14_bF$buf0 ;
wire areg_14_bF$buf1 ;
wire areg_14_bF$buf2 ;
wire areg_14_bF$buf3 ;
wire areg_14_bF$buf4 ;
wire _5892_ ;
wire _5472_ ;
wire _5052_ ;
wire _6677_ ;
wire _6257_ ;
wire _1392_ ;
wire _10675_ ;
wire _10255_ ;
wire _2597_ ;
wire _2177_ ;
wire _8823_ ;
wire _8403_ ;
wire _9608_ ;
wire _4743_ ;
wire _4323_ ;
wire _5948_ ;
wire _5528_ ;
wire _5108_ ;
wire _22_ ;
wire _9781_ ;
wire _9361_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _5281_ ;
wire _779_ ;
wire _359_ ;
wire _6486_ ;
wire _6066_ ;
wire _10484_ ;
wire _10064_ ;
wire _8632_ ;
wire _8212_ ;

NOR3X1 _21787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_3_),
    .C(_6_),
    .Y(_8_)
);

OAI21X1 _21367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_5921__bF$buf3),
    .C(_11155_),
    .Y(_11457_)
);

NAND2X1 _17915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_29_bF$buf3),
    .Y(_7672_)
);

OAI21X1 _12630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10244_),
    .B(_10178_),
    .C(_10035_),
    .Y(_10255_)
);

OAI21X1 _12210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5409_),
    .B(_5343_),
    .C(_5640_),
    .Y(_5651_)
);

FILL FILL74120x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3199_),
    .B(_3202_),
    .C(_3197_),
    .Y(_3203_)
);

NAND3X1 _13415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .B(_2741_),
    .C(_2742_),
    .Y(_2743_)
);

BUFX2 _23933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[51]),
    .Y(y[51])
);

NOR2X1 _23513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf1),
    .B(_7225__bF$buf2),
    .Y(_1894_)
);

AOI21X1 _18873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8714_),
    .B(_8722_),
    .C(_8701_),
    .Y(_8723_)
);

NOR2X1 _18453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8221_),
    .B(_8217_),
    .Y(_8263_)
);

NAND2X1 _18033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_7802_)
);

NAND3X1 _20638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10341_),
    .B(_10641_),
    .C(_10648_),
    .Y(_10658_)
);

AOI21X1 _20218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9897_),
    .B(_9895_),
    .C(_10196_),
    .Y(_10197_)
);

OAI21X1 _19658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9577_),
    .B(_9583_),
    .C(_9390_),
    .Y(_9584_)
);

AOI21X1 _19238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9122_),
    .B(_9118_),
    .C(_9102_),
    .Y(_9123_)
);

NAND2X1 _14793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf2),
    .B(areg_22_bF$buf1),
    .Y(_4250_)
);

NOR2X1 _14373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3790_),
    .Y(_3791_)
);

DFFPOSX1 _24051_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[9]),
    .CLK(clk_bF$buf1),
    .D(b[9])
);

OAI21X1 _15998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .B(_5569_),
    .C(_5568_),
    .Y(_5571_)
);

NAND2X1 _15578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf4),
    .B(areg_14_bF$buf2),
    .Y(_5110_)
);

AOI21X1 _15158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4613_),
    .B(_4617_),
    .C(_4352_),
    .Y(_4650_)
);

FILL SFILL59320x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10385_),
    .B(_10381_),
    .C(_10351_),
    .Y(_10387_)
);

FILL SFILL3400x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11705_),
    .B(_11704_),
    .C(_11706_),
    .Y(_11707_)
);

OAI21X1 _21176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11245_),
    .B(_11247_),
    .C(_11225_),
    .Y(_11248_)
);

OAI21X1 _17724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7461_),
    .B(_7462_),
    .C(_7457_),
    .Y(_7463_)
);

OAI21X1 _17304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6638_),
    .B(_6644_),
    .C(_6646_),
    .Y(_7003_)
);

NAND3X1 _18929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8766_),
    .B(_8756_),
    .C(_8762_),
    .Y(_8784_)
);

NAND3X1 _18509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8283_),
    .B(_8323_),
    .C(_8318_),
    .Y(_8324_)
);

FILL FILL74200x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_15_bF$buf1),
    .Y(_2993_)
);

OR2X2 _13224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2533_),
    .B(_2532_),
    .Y(_2534_)
);

XNOR2X1 _23742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2143_),
    .Y(_2144_)
);

AND2X2 _23322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(_1684_),
    .Y(_1687_)
);

AOI21X1 _14849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4306_),
    .B(_4307_),
    .C(_4305_),
    .Y(_4312_)
);

NAND3X1 _14429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3850_),
    .B(_3849_),
    .C(_3851_),
    .Y(_3852_)
);

AOI22X1 _14009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_16_bF$buf0),
    .C(breg_4_bF$buf5),
    .D(areg_15_bF$buf3),
    .Y(_3392_)
);

NAND3X1 _18682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8497_),
    .B(_8490_),
    .C(_8502_),
    .Y(_8513_)
);

AOI21X1 _18262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8045_),
    .B(_8053_),
    .C(_7657_),
    .Y(_8054_)
);

NAND2X1 _20867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10904_),
    .B(_10908_),
    .Y(_10909_)
);

OAI21X1 _20447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10201_),
    .B(_10193_),
    .C(_10203_),
    .Y(_10448_)
);

AOI22X1 _20027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9975_),
    .B(_9980_),
    .C(_9623_),
    .D(_9628_),
    .Y(_9987_)
);

NOR2X1 _19887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9833_),
    .B(_9834_),
    .Y(_9835_)
);

NAND3X1 _19467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9371_),
    .B(_9372_),
    .C(_9373_),
    .Y(_9374_)
);

OAI21X1 _19047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_8902_),
    .Y(_8913_)
);

AOI21X1 _14182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3354_),
    .B(_3311_),
    .C(_3349_),
    .Y(_3582_)
);

FILL SFILL8680x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1456_),
    .Y(_1467_)
);

NAND2X1 _15387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4900_),
    .B(_4901_),
    .Y(_4902_)
);

FILL SFILL13640x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert120 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf0)
);

BUFX2 BUFX2_insert121 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .Y(_3646__bF$buf3)
);

BUFX2 BUFX2_insert122 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .Y(_3646__bF$buf2)
);

BUFX2 BUFX2_insert123 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .Y(_3646__bF$buf1)
);

BUFX2 BUFX2_insert124 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646_),
    .Y(_3646__bF$buf0)
);

NOR2X1 _17953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7278_),
    .B(_7713_),
    .Y(_7714_)
);

AOI21X1 _17533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7241_),
    .B(_7240_),
    .C(_7236_),
    .Y(_7253_)
);

BUFX2 BUFX2_insert125 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf5)
);

BUFX2 BUFX2_insert126 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf4)
);

AOI21X1 _17113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6398_),
    .C(_6401_),
    .Y(_6794_)
);

BUFX2 BUFX2_insert127 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf3)
);

BUFX2 BUFX2_insert128 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf2)
);

BUFX2 BUFX2_insert129 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf1)
);

FILL SFILL13560x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8123_),
    .B(_8155_),
    .C(_8573_),
    .Y(_8574_)
);

NOR3X1 _18318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8099_),
    .B(_8085_),
    .C(_8105_),
    .Y(_8114_)
);

AOI21X1 _13873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_3216_),
    .C(_2987_),
    .Y(_3244_)
);

XOR2X1 _13453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .B(_2778_),
    .Y(_2784_)
);

DFFPOSX1 _23971_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[25]),
    .CLK(clk_bF$buf7),
    .D(_0_[25])
);

AOI21X1 _13033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_900_),
    .C(_932_),
    .Y(_2328_)
);

NAND3X1 _23551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1934_),
    .B(_1935_),
    .C(_1931_),
    .Y(_1937_)
);

NAND2X1 _23131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1435_),
    .B(_1431_),
    .Y(_1479_)
);

FILL SFILL64280x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_15_bF$buf5),
    .Y(_4102_)
);

AND2X2 _14238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf5),
    .B(areg_13_bF$buf0),
    .Y(_3643_)
);

FILL SFILL64200x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_24_bF$buf1),
    .Y(_8305_)
);

OAI21X1 _18071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6970_),
    .B(_7825_),
    .C(_7388_),
    .Y(_7844_)
);

NOR2X1 _20676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf0),
    .B(_7225__bF$buf4),
    .Y(_10699_)
);

INVX2 _20256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10211_),
    .Y(_10239_)
);

NAND3X1 _16804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6444_),
    .B(_6452_),
    .C(_6453_),
    .Y(_6454_)
);

NAND3X1 _19696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9269_),
    .B(_9621_),
    .C(_9619_),
    .Y(_9626_)
);

OAI21X1 _19276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9161_),
    .B(_9162_),
    .C(_9164_),
    .Y(_9165_)
);

NAND3X1 _12724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11264_),
    .B(_11275_),
    .C(_11253_),
    .Y(_11286_)
);

AOI21X1 _12304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6549_),
    .B(_6505_),
    .C(_6461_),
    .Y(_6681_)
);

OAI21X1 _22822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf2),
    .B(_5676_),
    .C(_1141_),
    .Y(_1142_)
);

OAI21X1 _22402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_673_),
    .C(_676_),
    .Y(_682_)
);

OAI21X1 _15196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf3),
    .B(_3529__bF$buf3),
    .C(_4688_),
    .Y(_4692_)
);

NAND3X1 _13929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3291_),
    .B(_3302_),
    .C(_3294_),
    .Y(_3305_)
);

NAND2X1 _13509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_11_bF$buf0),
    .Y(_2845_)
);

NAND2X1 _23607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_1896_),
    .Y(_1997_)
);

OAI21X1 _17762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7501_),
    .B(_7502_),
    .C(_7504_),
    .Y(_7505_)
);

INVX2 _17342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7017_),
    .Y(_7045_)
);

OAI21X1 _18967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8690_),
    .B(_8689_),
    .C(_8602_),
    .Y(_8826_)
);

AOI21X1 _18547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_30_bF$buf3),
    .C(_8346_),
    .Y(_8366_)
);

NOR2X1 _18127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7892_),
    .B(_7890_),
    .Y(_7905_)
);

OAI21X1 _13682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2838_),
    .B(_2794_),
    .C(_2828_),
    .Y(_3035_)
);

OAI21X1 _13262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2574_),
    .B(_2378_),
    .C(_2409_),
    .Y(_2575_)
);

XNOR2X1 _23780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2183_),
    .B(_2171_),
    .Y(_2184_)
);

AOI21X1 _23360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1572_),
    .C(_1610_),
    .Y(_1728_)
);

OR2X2 _14887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_4068_),
    .Y(_4353_)
);

AOI21X1 _14467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3886_),
    .B(_3893_),
    .C(_3873_),
    .Y(_3894_)
);

OAI21X1 _14047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3432_),
    .B(_3433_),
    .C(_3431_),
    .Y(_3434_)
);

FILL SFILL8600x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53800x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10481_),
    .B(_10489_),
    .C(_10468_),
    .Y(_10490_)
);

NAND3X1 _20065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10014_),
    .B(_10006_),
    .C(_10018_),
    .Y(_10029_)
);

INVX2 _16613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6222_),
    .Y(_6245_)
);

NOR2X1 _19085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8541_),
    .B(_8605_),
    .Y(_8955_)
);

FILL SFILL74200x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7559_),
    .B(_7485_),
    .C(_7565_),
    .Y(_7566_)
);

FILL SFILL44040x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1870_),
    .Y(_1881_)
);

AOI21X1 _12533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7678_),
    .B(_7722_),
    .C(_7744_),
    .Y(_9192_)
);

AOI22X1 _22631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_929_),
    .C(_928_),
    .D(_10673_),
    .Y(_933_)
);

NAND3X1 _12113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4533_),
    .B(_4577_),
    .C(_4237_),
    .Y(_4588_)
);

NAND3X1 _22211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .B(_469_),
    .C(_470_),
    .Y(_474_)
);

FILL SFILL64280x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2868_),
    .B(_2900_),
    .C(_2917_),
    .Y(_3096_)
);

OAI22X1 _13318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2174_),
    .B(_2635_),
    .C(_2450_),
    .D(_2454_),
    .Y(_2636_)
);

NAND2X1 _23836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2243_),
    .B(_2230_),
    .Y(_2244_)
);

NAND2X1 _23416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_26_bF$buf0),
    .B(breg_27_bF$buf1),
    .Y(_1789_)
);

BUFX2 BUFX2_insert500 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190_),
    .Y(_5190__bF$buf3)
);

FILL SFILL64200x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert501 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190_),
    .Y(_5190__bF$buf2)
);

BUFX2 BUFX2_insert502 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190_),
    .Y(_5190__bF$buf1)
);

BUFX2 BUFX2_insert503 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190_),
    .Y(_5190__bF$buf0)
);

OAI21X1 _17991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7740_),
    .B(_7739_),
    .C(_7737_),
    .Y(_7756_)
);

BUFX2 BUFX2_insert504 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869_),
    .Y(_10869__bF$buf3)
);

NAND3X1 _17571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7275_),
    .B(_7288_),
    .C(_7293_),
    .Y(_7295_)
);

BUFX2 BUFX2_insert505 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869_),
    .Y(_10869__bF$buf2)
);

NAND3X1 _17151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(_6830_),
    .C(_6829_),
    .Y(_6835_)
);

BUFX2 BUFX2_insert506 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869_),
    .Y(_10869__bF$buf1)
);

BUFX2 BUFX2_insert507 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869_),
    .Y(_10869__bF$buf0)
);

BUFX2 BUFX2_insert508 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .Y(_3961__bF$buf4)
);

BUFX2 BUFX2_insert509 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .Y(_3961__bF$buf3)
);

AOI21X1 _18776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8613_),
    .B(_8615_),
    .C(_8611_),
    .Y(_8616_)
);

NAND3X1 _18356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8123_),
    .B(_8151_),
    .C(_8155_),
    .Y(_8156_)
);

NOR2X1 _13491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2634_),
    .Y(_2826_)
);

OAI21X1 _13071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11712_),
    .B(_1511_),
    .C(_2364_),
    .Y(_2366_)
);

FILL SFILL9080x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_134_),
    .C(_130_),
    .Y(_135_)
);

FILL SFILL54200x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3868_),
    .B(_3902_),
    .C(_3911_),
    .Y(_4144_)
);

AND2X2 _14276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf2),
    .B(areg_20_bF$buf3),
    .Y(_3685_)
);

FILL SFILL39000x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10267_),
    .B(_10270_),
    .C(_10208_),
    .Y(_10281_)
);

AOI21X1 _16842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6493_),
    .B(_6495_),
    .C(_6492_),
    .Y(_6496_)
);

NAND3X1 _16422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6029_),
    .B(_6032_),
    .C(_5658_),
    .Y(_6035_)
);

NAND3X1 _16002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5568_),
    .C(_5562_),
    .Y(_5576_)
);

FILL SFILL69320x50 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _21499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11600_),
    .Y(_11601_)
);

AND2X2 _21079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf4),
    .B(areg_23_bF$buf3),
    .Y(_11141_)
);

NOR2X1 _17627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7354_),
    .B(_7355_),
    .Y(_7356_)
);

NOR2X1 _17207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6473_),
    .B(_6895_),
    .Y(_6896_)
);

INVX1 _12762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11690_),
    .Y(_11701_)
);

OAI21X1 _12342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7087_),
    .B(_7065_),
    .C(_5859_),
    .Y(_7098_)
);

NAND3X1 _22860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1104_),
    .B(_1179_),
    .C(_1182_),
    .Y(_1183_)
);

AOI21X1 _22440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_695_),
    .C(_497_),
    .Y(_723_)
);

NAND2X1 _22020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .B(breg_27_bF$buf4),
    .Y(_263_)
);

AOI21X1 _13967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3341_),
    .B(_3342_),
    .C(_3340_),
    .Y(_3346_)
);

NOR2X1 _13547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2881_),
    .B(_2882_),
    .Y(_2887_)
);

NAND2X1 _13127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf1),
    .B(areg_9_bF$buf4),
    .Y(_2427_)
);

XNOR2X1 _23645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .B(_2028_),
    .Y(_2039_)
);

OAI21X1 _23225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1578_),
    .C(_1579_),
    .Y(_1580_)
);

FILL SFILL13720x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6651_),
    .B(_7085_),
    .C(_6660_),
    .Y(_7086_)
);

AOI21X1 _18585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8405_),
    .B(_8406_),
    .C(_8404_),
    .Y(_8407_)
);

AOI21X1 _18165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7516_),
    .B(_7521_),
    .C(_7523_),
    .Y(_7947_)
);

AOI21X1 _21711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11703_),
    .B(_11707_),
    .C(_11604_),
    .Y(_11834_)
);

INVX2 _14085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3246_),
    .Y(_3476_)
);

NOR2X1 _12818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf0),
    .B(_5190__bF$buf1),
    .Y(_407_)
);

NOR3X1 _22916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_948_),
    .B(_1074_),
    .C(_1079_),
    .Y(_1245_)
);

INVX2 _16651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6267_),
    .Y(_6287_)
);

AOI21X1 _16231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5817_),
    .B(_5810_),
    .C(_5779_),
    .Y(_5827_)
);

FILL SFILL28840x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7600_),
    .B(_7601_),
    .C(_7343_),
    .Y(_7608_)
);

NAND3X1 _17436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7145_),
    .B(_7147_),
    .C(_7146_),
    .Y(_7148_)
);

OAI21X1 _17016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_6686__bF$buf1),
    .C(_6683_),
    .Y(_6687_)
);

OR2X2 _12991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_2280_),
    .Y(_2286_)
);

OAI21X1 _12571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9565_),
    .B(_9576_),
    .C(_8544_),
    .Y(_9609_)
);

OAI21X1 _12151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4566_),
    .B(_4544_),
    .C(_4478_),
    .Y(_5003_)
);

FILL SFILL54200x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3111_),
    .B(_3130_),
    .Y(_3137_)
);

OAI21X1 _13356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2676_),
    .C(_2660_),
    .Y(_2678_)
);

INVX1 _23874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2265_),
    .Y(_2284_)
);

NOR2X1 _23454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1826_),
    .Y(_1831_)
);

OAI21X1 _23034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1366_),
    .C(_1363_),
    .Y(_1373_)
);

FILL SFILL18840x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5473_),
    .B(_5482_),
    .C(_5483_),
    .Y(_5488_)
);

INVX2 _15502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5022_),
    .Y(_5027_)
);

AND2X2 _18394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_18_bF$buf1),
    .Y(_8198_)
);

OAI21X1 _20999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11050_),
    .B(_11049_),
    .C(_11048_),
    .Y(_11053_)
);

OAI21X1 _20579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10587_),
    .B(_10588_),
    .C(_10263_),
    .Y(_10593_)
);

NAND3X1 _20159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10126_),
    .B(_10128_),
    .C(_10127_),
    .Y(_10132_)
);

NAND3X1 _16707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6347_),
    .B(_6346_),
    .C(_6345_),
    .Y(_6348_)
);

NOR2X1 _21940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_8773_),
    .Y(_176_)
);

AOI21X1 _21520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11619_),
    .B(_11623_),
    .C(_11610_),
    .Y(_11624_)
);

OAI21X1 _21100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11146_),
    .B(_11150_),
    .C(_11139_),
    .Y(_11164_)
);

AOI21X1 _19599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9502_),
    .B(_9508_),
    .C(_9487_),
    .Y(_9519_)
);

AOI21X1 _19179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9047_),
    .B(_9046_),
    .C(_9044_),
    .Y(_9058_)
);

FILL SFILL48920x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10046_),
    .B(_10200_),
    .C(_10221_),
    .Y(_10232_)
);

NAND2X1 _12207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5497_),
    .B(_5563_),
    .Y(_5618_)
);

NOR2X1 _22725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .B(_1035_),
    .Y(_1036_)
);

AOI21X1 _22305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_566_),
    .C(_544_),
    .Y(_576_)
);

OAI21X1 _15099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4488_),
    .B(_4484_),
    .C(_4491_),
    .Y(_4586_)
);

NAND3X1 _16880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6531_),
    .B(_6532_),
    .C(_6536_),
    .Y(_6537_)
);

AOI21X1 _16460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6065_),
    .B(_6064_),
    .C(_6061_),
    .Y(_6075_)
);

OAI21X1 _16040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5610_),
    .B(_5611_),
    .C(_5463_),
    .Y(_5617_)
);

OAI21X1 _17665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf1),
    .B(_3146__bF$buf1),
    .C(_6606_),
    .Y(_7398_)
);

AND2X2 _17245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_18_bF$buf2),
    .Y(_6938_)
);

NAND2X1 _12380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7470_),
    .B(_7371_),
    .Y(_7514_)
);

FILL SFILL38920x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2833_),
    .B(_2828_),
    .C(_2794_),
    .Y(_2929_)
);

OAI21X1 _13165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2468_),
    .B(_2462_),
    .C(_2459_),
    .Y(_2469_)
);

XNOR2X1 _23683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2079_),
    .B(_2070_),
    .Y(_2080_)
);

AOI21X1 _23263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1614_),
    .B(_1615_),
    .C(_1613_),
    .Y(_1623_)
);

FILL SFILL3560x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9745_),
    .B(_9744_),
    .C(_9742_),
    .Y(_9752_)
);

DFFPOSX1 _24048_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[6]),
    .CLK(clk_bF$buf10),
    .D(b[6])
);

FILL SFILL28920x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4967_),
    .B(_5277_),
    .C(_5270_),
    .Y(_5279_)
);

NOR2X1 _15311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_2669__bF$buf2),
    .Y(_4819_)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf0)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf4)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf3)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf2)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf1)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf0)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[21]),
    .Y(areg_21_bF$buf4)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[21]),
    .Y(areg_21_bF$buf3)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[21]),
    .Y(areg_21_bF$buf2)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[21]),
    .Y(areg_21_bF$buf1)
);

AOI21X1 _20388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10378_),
    .B(_10379_),
    .C(_10354_),
    .Y(_10383_)
);

NAND3X1 _16936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6596_),
    .B(_6598_),
    .C(_6597_),
    .Y(_6599_)
);

NAND2X1 _16516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_20_bF$buf3),
    .Y(_6138_)
);

OAI21X1 _12856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_779_),
    .C(_735_),
    .Y(_823_)
);

NAND3X1 _12436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8084_),
    .B(_8117_),
    .C(_7196_),
    .Y(_8128_)
);

AND2X2 _22954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1270_),
    .B(_1269_),
    .Y(_1286_)
);

NAND2X1 _12016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf4),
    .B(breg_3_bF$buf0),
    .Y(_3525_)
);

NAND3X1 _22534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(_826_),
    .C(_825_),
    .Y(_827_)
);

NAND2X1 _22114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_168_),
    .Y(_366_)
);

FILL SFILL18840x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668__bF$buf0),
    .B(_8773_),
    .C(_2072_),
    .Y(_2140_)
);

XNOR2X1 _23319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1682_),
    .B(_1677_),
    .Y(_1683_)
);

OAI21X1 _17894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7640_),
    .B(_7644_),
    .C(_7648_),
    .Y(_7649_)
);

NAND3X1 _17474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7170_),
    .B(_7176_),
    .C(_7179_),
    .Y(_7189_)
);

NAND3X1 _17054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6652_),
    .B(_6675_),
    .C(_6674_),
    .Y(_6729_)
);

FILL SFILL74360x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10609_),
    .B(_10615_),
    .C(_10461_),
    .Y(_10616_)
);

NOR3X1 _18679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8508_),
    .B(_8504_),
    .C(_8507_),
    .Y(_8509_)
);

AOI21X1 _18259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8036_),
    .B(_8037_),
    .C(_7663_),
    .Y(_8050_)
);

NAND3X1 _13394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2710_),
    .C(_2713_),
    .Y(_2720_)
);

NAND2X1 _23492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1869_),
    .B(_1871_),
    .Y(_1872_)
);

NOR2X1 _23072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf4),
    .B(_6815__bF$buf4),
    .Y(_1414_)
);

NAND3X1 _19620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_29_bF$buf3),
    .C(_9541_),
    .Y(_9542_)
);

OAI21X1 _19200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9064_),
    .B(_9069_),
    .C(_9072_),
    .Y(_9081_)
);

FILL SFILL69080x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11650_),
    .B(_11654_),
    .C(_11658_),
    .Y(_28_)
);

OAI21X1 _14599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4025_),
    .B(_4029_),
    .C(_3778_),
    .Y(_4039_)
);

NAND3X1 _14179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3572_),
    .B(_3577_),
    .C(_3576_),
    .Y(_3578_)
);

AOI21X1 _15960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5522_),
    .B(_5526_),
    .C(_5528_),
    .Y(_5529_)
);

NOR3X1 _15540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5061_),
    .B(_5064_),
    .C(_5060_),
    .Y(_5068_)
);

AOI21X1 _15120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4604_),
    .B(_4603_),
    .C(_4602_),
    .Y(_4609_)
);

FILL SFILL3640x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9818_),
    .B(_9820_),
    .C(_9825_),
    .Y(_10174_)
);

NAND3X1 _16745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6370_),
    .B(_6377_),
    .C(_6380_),
    .Y(_6390_)
);

NAND2X1 _16325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf0),
    .B(areg_25_bF$buf2),
    .Y(_5930_)
);

FILL SFILL59080x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10441_),
    .B(_10573_),
    .C(_10628_),
    .Y(_10639_)
);

OAI21X1 _12245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5705_),
    .B(_4204_),
    .C(_5792_),
    .Y(_6034_)
);

NOR3X1 _22763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .B(_1065_),
    .C(_1068_),
    .Y(_1078_)
);

AOI21X1 _22343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_380_),
    .C(_617_),
    .Y(_618_)
);

DFFPOSX1 _23968_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[22]),
    .CLK(clk_bF$buf2),
    .D(_0_[22])
);

NOR2X1 _23548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1924_),
    .B(_1834_),
    .Y(_1933_)
);

AOI21X1 _23128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1463_),
    .B(_1460_),
    .C(_1440_),
    .Y(_1475_)
);

FILL SFILL49080x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4257_),
    .B(_4253_),
    .C(_4241_),
    .Y(_4271_)
);

AOI21X1 _17283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6968_),
    .B(_6965_),
    .C(_6962_),
    .Y(_6980_)
);

OAI21X1 _18488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8296_),
    .B(_8300_),
    .C(_8289_),
    .Y(_8301_)
);

OAI22X1 _18068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7018_),
    .B(_7838_),
    .C(_7839_),
    .D(_7439_),
    .Y(_7840_)
);

INVX1 _11936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf4),
    .Y(_2650_)
);

OAI21X1 _21614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11453_),
    .B(_11447_),
    .C(_11456_),
    .Y(_11727_)
);

FILL SFILL39320x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315__bF$buf2),
    .B(_6300__bF$buf2),
    .C(_984_),
    .Y(_1138_)
);

FILL SFILL8760x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6267_),
    .B(_6288_),
    .C(_6284_),
    .Y(_6641_)
);

NAND3X1 _16554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6172_),
    .B(_6175_),
    .C(_6179_),
    .Y(_6180_)
);

NOR2X1 _16134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5337_),
    .B(_5719_),
    .Y(_5720_)
);

FILL SFILL53960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7496_),
    .B(_7497_),
    .C(_7488_),
    .Y(_7501_)
);

AOI21X1 _17339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7030_),
    .B(_7029_),
    .C(_7026_),
    .Y(_7041_)
);

AOI21X1 _12894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9850_),
    .B(_9861_),
    .C(_8467_),
    .Y(_1239_)
);

OAI21X1 _12474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8533_),
    .B(_7272_),
    .C(_8008_),
    .Y(_8544_)
);

NOR3X1 _22992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .B(_1320_),
    .C(_1322_),
    .Y(_1327_)
);

NAND3X1 _12054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .B(_3887_),
    .C(_3920_),
    .Y(_3942_)
);

AOI22X1 _22572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_31_bF$buf2),
    .C(breg_17_bF$buf2),
    .D(areg_30_bF$buf1),
    .Y(_869_)
);

OAI21X1 _22152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_408_),
    .C(_404_),
    .Y(_409_)
);

NAND2X1 _18700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_24_bF$buf3),
    .Y(_8532_)
);

OAI21X1 _13679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3021_),
    .B(_3023_),
    .C(_3027_),
    .Y(_3031_)
);

NAND2X1 _13259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2369_),
    .B(_2570_),
    .Y(_2571_)
);

XOR2X1 _23777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2178_),
    .B(_2180_),
    .Y(_2181_)
);

AOI21X1 _23357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1593_),
    .B(_1596_),
    .C(_1720_),
    .Y(_1725_)
);

FILL SFILL3720x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9568_),
    .B(_9528_),
    .C(_9567_),
    .Y(_9855_)
);

OAI21X1 _14620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3798_),
    .B(_3783_),
    .C(_3804_),
    .Y(_4060_)
);

NAND2X1 _14200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_11_bF$buf3),
    .Y(_3601_)
);

NAND3X1 _17092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6764_),
    .B(_6770_),
    .C(_6509_),
    .Y(_6771_)
);

FILL SFILL43880x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48920x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _15825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5380_),
    .Y(_5381_)
);

OAI21X1 _15405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4920_),
    .B(_4921_),
    .C(_4919_),
    .Y(_4922_)
);

NAND2X1 _18297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8089_),
    .B(_8090_),
    .Y(_8091_)
);

NOR3X1 _21843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11680_),
    .B(_11681_),
    .C(_11683_),
    .Y(_70_)
);

NAND2X1 _21423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11197_),
    .B(_11205_),
    .Y(_11519_)
);

OAI21X1 _21003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10782_),
    .B(_10784_),
    .C(_10774_),
    .Y(_11058_)
);

FILL SFILL33880x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10649_),
    .B(_10653_),
    .C(_10656_),
    .Y(_929_)
);

NAND3X1 _22208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_459_),
    .C(_450_),
    .Y(_470_)
);

FILL SFILL49080x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf0),
    .B(_5668__bF$buf2),
    .C(_6049_),
    .Y(_6431_)
);

AOI21X1 _16363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5966_),
    .B(_5965_),
    .C(_5964_),
    .Y(_5972_)
);

FILL SFILL18600x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert470 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[20]),
    .Y(breg_20_bF$buf2)
);

BUFX2 BUFX2_insert471 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[20]),
    .Y(breg_20_bF$buf1)
);

BUFX2 BUFX2_insert472 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[20]),
    .Y(breg_20_bF$buf0)
);

BUFX2 BUFX2_insert473 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[17]),
    .Y(breg_17_bF$buf4)
);

NOR2X1 _17988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7307_),
    .B(_7751_),
    .Y(_7752_)
);

BUFX2 BUFX2_insert474 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[17]),
    .Y(breg_17_bF$buf3)
);

FILL SFILL18840x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf2),
    .B(_3781__bF$buf2),
    .C(_6863_),
    .Y(_7291_)
);

BUFX2 BUFX2_insert475 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[17]),
    .Y(breg_17_bF$buf2)
);

AOI21X1 _17148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6830_),
    .B(_6829_),
    .C(_6828_),
    .Y(_6831_)
);

BUFX2 BUFX2_insert476 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[17]),
    .Y(breg_17_bF$buf1)
);

BUFX2 BUFX2_insert477 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[17]),
    .Y(breg_17_bF$buf0)
);

BUFX2 BUFX2_insert478 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf3)
);

BUFX2 BUFX2_insert479 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf2)
);

AOI21X1 _12283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5135_),
    .B(_5201_),
    .C(_6439_),
    .Y(_6450_)
);

NOR2X1 _22381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_658_),
    .B(_650_),
    .Y(_660_)
);

FILL SFILL54280x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .B(_2818_),
    .C(_2805_),
    .Y(_2822_)
);

INVX8 _13068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf4),
    .Y(_2362_)
);

NAND2X1 _23586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11877_),
    .B(_1973_),
    .Y(_1974_)
);

FILL SFILL23800x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _23166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1513_),
    .C(_1510_),
    .Y(_1517_)
);

NAND2X1 _19714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9360_),
    .B(_9370_),
    .Y(_9645_)
);

FILL SFILL39000x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5167_),
    .B(_5169_),
    .C(_5171_),
    .Y(_5172_)
);

NAND2X1 _15214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_17_bF$buf4),
    .Y(_4712_)
);

INVX1 _16839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6438_),
    .Y(_6492_)
);

OAI21X1 _16419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6030_),
    .B(_6031_),
    .C(_5646_),
    .Y(_6032_)
);

NOR2X1 _11974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_3055_),
    .Y(_3066_)
);

OAI22X1 _21652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11230_),
    .B(_11528_),
    .C(_11526_),
    .D(_11768_),
    .Y(_11769_)
);

OAI21X1 _21232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11296_),
    .B(_11300_),
    .C(_11303_),
    .Y(_11309_)
);

OAI21X1 _12759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10321_),
    .B(_8665_),
    .C(_10397_),
    .Y(_11668_)
);

AOI21X1 _12339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7032_),
    .B(_7031_),
    .C(_5804_),
    .Y(_7065_)
);

AOI21X1 _22857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1176_),
    .B(_1177_),
    .C(_1175_),
    .Y(_1180_)
);

NAND2X1 _22437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11877_),
    .B(_10688_),
    .Y(_720_)
);

AND2X2 _22017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_28_bF$buf1),
    .Y(_260_)
);

FILL SFILL43960x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2796_),
    .B(_3053_),
    .Y(_3054_)
);

NAND2X1 _16592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf1),
    .B(breg_14_bF$buf3),
    .Y(_6222_)
);

NAND2X1 _16172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5757_),
    .B(_5755_),
    .Y(_5762_)
);

AND2X2 _14905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4076_),
    .B(_4371_),
    .Y(_4373_)
);

AOI21X1 _17797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7537_),
    .B(_7539_),
    .C(_7529_),
    .Y(_7543_)
);

OAI21X1 _17377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7080_),
    .B(_7081_),
    .C(_7082_),
    .Y(_7083_)
);

AOI21X1 _12092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3613_),
    .B(_3657_),
    .C(_4346_),
    .Y(_4357_)
);

OAI21X1 _22190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_449_),
    .C(_249_),
    .Y(_450_)
);

FILL SFILL64360x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10969_),
    .B(_10970_),
    .C(_10967_),
    .Y(_10971_)
);

NAND3X1 _20503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10500_),
    .B(_10508_),
    .C(_10509_),
    .Y(_10510_)
);

NAND3X1 _13297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2609_),
    .C(_2611_),
    .Y(_2612_)
);

NAND3X1 _23395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .B(_1766_),
    .C(_1764_),
    .Y(_1767_)
);

NAND3X1 _19943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9891_),
    .B(_9856_),
    .C(_9895_),
    .Y(_9896_)
);

OAI21X1 _19523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf2),
    .B(_3958__bF$buf3),
    .C(_9430_),
    .Y(_9436_)
);

AND2X2 _19103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8552_),
    .B(_8545_),
    .Y(_8975_)
);

FILL SFILL33880x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11541_),
    .B(_11828_),
    .C(_11829_),
    .Y(_11830_)
);

NAND3X1 _15863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5415_),
    .B(_5418_),
    .C(_5422_),
    .Y(_5423_)
);

INVX1 _15443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4648_),
    .Y(_4962_)
);

AND2X2 _15023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_16_bF$buf2),
    .Y(_4503_)
);

FILL SFILL28760x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6272_),
    .B(_6271_),
    .C(_6268_),
    .Y(_6283_)
);

OAI21X1 _16228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5506_),
    .B(_5499_),
    .C(_5509_),
    .Y(_5823_)
);

NAND2X1 _21881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11732_),
    .B(_110_),
    .Y(_112_)
);

FILL SFILL23880x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11555_),
    .B(_11556_),
    .C(_11554_),
    .Y(_11561_)
);

NOR3X1 _21041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11092_),
    .B(_11093_),
    .C(_11095_),
    .Y(_11100_)
);

NAND2X1 _12988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf2),
    .B(areg_12_bF$buf1),
    .Y(_2259_)
);

AOI21X1 _12568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9422_),
    .B(_9466_),
    .C(_8698_),
    .Y(_9576_)
);

FILL SFILL23800x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4862_),
    .B(_4873_),
    .C(_4051_),
    .Y(_4970_)
);

NOR2X1 _22666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(_970_),
    .Y(_971_)
);

NOR2X1 _22246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_510_),
    .Y(_511_)
);

FILL SFILL13880x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_11_bF$buf3),
    .Y(_4164_)
);

OAI21X1 _17186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6868_),
    .B(_6869_),
    .C(_6872_),
    .Y(_6873_)
);

FILL SFILL13800x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .B(_5482_),
    .C(_5473_),
    .Y(_5484_)
);

NOR3X1 _20732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10744_),
    .B(_10747_),
    .C(_10749_),
    .Y(_10761_)
);

AOI21X1 _20312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9950_),
    .B(_9952_),
    .C(_10300_),
    .Y(_10301_)
);

AND2X2 _19752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9682_),
    .B(_9686_),
    .Y(_9687_)
);

OAI21X1 _19332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9219_),
    .B(_9226_),
    .C(_8890_),
    .Y(_9227_)
);

FILL SFILL74440x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_167_),
    .B(_168_),
    .C(_169_),
    .Y(_173_)
);

NOR2X1 _21517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11617_),
    .B(_11620_),
    .Y(_11621_)
);

OAI21X1 _15672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5209_),
    .B(_5208_),
    .C(_5194_),
    .Y(_5214_)
);

AOI21X1 _15252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4751_),
    .B(_4747_),
    .C(_4753_),
    .Y(_4754_)
);

FILL SFILL64040x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6139_),
    .B(_6533_),
    .Y(_6534_)
);

OAI22X1 _16457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5373_),
    .B(_6070_),
    .C(_6071_),
    .D(_5747_),
    .Y(_6072_)
);

NAND3X1 _16037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5368_),
    .B(_5459_),
    .C(_5458_),
    .Y(_5614_)
);

NOR2X1 _21690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11238_),
    .B(_11809_),
    .Y(_11810_)
);

AOI21X1 _21270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11347_),
    .B(_11348_),
    .C(_11334_),
    .Y(_11349_)
);

FILL SFILL64360x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_7_bF$buf1),
    .Y(_177_)
);

NAND2X1 _12377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7470_),
    .B(_7459_),
    .Y(_7481_)
);

AOI21X1 _22895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .B(_1182_),
    .C(_1104_),
    .Y(_1222_)
);

NAND3X1 _22475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_750_),
    .C(_755_),
    .Y(_762_)
);

NAND2X1 _22055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_25_bF$buf2),
    .Y(_302_)
);

NAND3X1 _18603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8408_),
    .B(_8414_),
    .C(_8279_),
    .Y(_8427_)
);

FILL SFILL54040x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9645_),
    .B(_9743_),
    .C(_9747_),
    .Y(_9748_)
);

INVX2 _14943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4391_),
    .Y(_4415_)
);

OAI21X1 _14523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3678_),
    .B(_3682_),
    .C(_3686_),
    .Y(_3956_)
);

AOI22X1 _14103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2983_),
    .B(_3495_),
    .C(_3486_),
    .D(_3480_),
    .Y(_3496_)
);

AOI21X1 _15728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5273_),
    .B(_5274_),
    .C(_5265_),
    .Y(_5275_)
);

INVX1 _15308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4504_),
    .Y(_4815_)
);

INVX2 _20961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11010_),
    .Y(_11012_)
);

NOR3X1 _20541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10544_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10552_)
);

NAND3X1 _20121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10089_),
    .B(_10083_),
    .C(_10041_),
    .Y(_10091_)
);

OAI21X1 _19981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9930_),
    .B(_9936_),
    .C(_9756_),
    .Y(_9938_)
);

AOI21X1 _19561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9472_),
    .B(_9471_),
    .C(_9473_),
    .Y(_9478_)
);

INVX2 _19141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9015_),
    .Y(_9017_)
);

NAND2X1 _21746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11591_),
    .B(_11870_),
    .Y(_11871_)
);

AOI21X1 _21326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11059_),
    .B(_11096_),
    .C(_11100_),
    .Y(_11412_)
);

FILL SFILL8840x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _15481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4998_),
    .B(_5000_),
    .Y(_5004_)
);

NAND2X1 _15061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_23_bF$buf3),
    .Y(_4545_)
);

NAND2X1 _16686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6318_),
    .B(_6311_),
    .Y(_6325_)
);

OAI21X1 _16266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5863_),
    .B(_5864_),
    .C(_5860_),
    .Y(_5865_)
);

FILL SFILL13800x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5376_),
    .B(_5365_),
    .C(_5299_),
    .Y(_5387_)
);

NAND2X1 _22284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf2),
    .B(breg_25_bF$buf1),
    .Y(_553_)
);

OAI21X1 _18832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8661_),
    .B(_8666_),
    .C(_8668_),
    .Y(_8678_)
);

XNOR2X1 _18412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8193_),
    .B(_8189_),
    .Y(_8218_)
);

FILL SFILL38680x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _23489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .Y(_1868_)
);

INVX1 _23069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1409_),
    .Y(_1410_)
);

NAND3X1 _19617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9534_),
    .B(_9538_),
    .C(_9536_),
    .Y(_9539_)
);

INVX2 _14752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4205_),
    .Y(_4206_)
);

OAI21X1 _14332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3735_),
    .B(_3728_),
    .C(_3590_),
    .Y(_3747_)
);

DFFPOSX1 _24010_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[0]),
    .CLK(clk_bF$buf8),
    .D(a[0])
);

NAND3X1 _15957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5526_)
);

OAI21X1 _15537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5060_),
    .B(_5061_),
    .C(_5064_),
    .Y(_5065_)
);

NAND3X1 _15117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4598_),
    .B(_4605_),
    .C(_4361_),
    .Y(_4606_)
);

AOI21X1 _20770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10786_),
    .B(_10793_),
    .C(_10740_),
    .Y(_10802_)
);

INVX1 _20350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10340_),
    .Y(_10341_)
);

NAND3X1 _19790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9688_),
    .B(_9723_),
    .C(_9727_),
    .Y(_9728_)
);

OAI21X1 _19370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9266_),
    .B(_8883_),
    .C(_9245_),
    .Y(_9267_)
);

NAND3X1 _21975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_212_),
    .C(_11888_),
    .Y(_215_)
);

AND2X2 _21555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11135_),
    .B(_11661_),
    .Y(_11662_)
);

AOI21X1 _21135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11184_),
    .B(_11191_),
    .C(_11169_),
    .Y(_11203_)
);

FILL SFILL59480x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _15290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4772_),
    .B(_4794_),
    .Y(_4795_)
);

AOI21X1 _13603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2577_),
    .B(_2717_),
    .C(_2948_),
    .Y(_2949_)
);

OR2X2 _23701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2097_),
    .B(_2060_),
    .Y(_2100_)
);

AOI21X1 _16495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5746_),
    .B(_5832_),
    .C(_5829_),
    .Y(_6115_)
);

NAND2X1 _16075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5653_),
    .B(_5646_),
    .Y(_5656_)
);

NOR3X1 _14808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3968_),
    .B(_3970_),
    .C(_3963_),
    .Y(_4267_)
);

FILL SFILL8520x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_62_),
    .C(_343_),
    .Y(_344_)
);

INVX1 _18641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8466_),
    .Y(_8468_)
);

NAND3X1 _18221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8002_),
    .B(_8003_),
    .C(_8001_),
    .Y(_8009_)
);

OAI21X1 _20826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10863_),
    .B(_10862_),
    .C(_10853_),
    .Y(_10864_)
);

OR2X2 _20406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10396_),
    .B(_10398_),
    .Y(_10403_)
);

NOR2X1 _23298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1658_),
    .B(_1659_),
    .Y(_1660_)
);

NAND2X1 _19846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9783_),
    .B(_9789_),
    .Y(_9790_)
);

INVX1 _19426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9322_),
    .Y(_9329_)
);

OAI21X1 _19006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8865_),
    .B(_8868_),
    .C(_8473_),
    .Y(_8869_)
);

INVX2 _14981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4455_),
    .Y(_4456_)
);

OAI21X1 _14561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3990_),
    .B(_3996_),
    .C(_3915_),
    .Y(_3998_)
);

NOR2X1 _14141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3533_),
    .B(_3535_),
    .Y(_3537_)
);

FILL SFILL69160x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf0),
    .B(_5315__bF$buf1),
    .C(_4973_),
    .Y(_5316_)
);

FILL SFILL74120x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_4857_)
);

OAI21X1 _21784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_11899_),
    .Y(_5_)
);

NOR3X1 _21364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11447_),
    .B(_11449_),
    .C(_11453_),
    .Y(_11454_)
);

NOR2X1 _17912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf1),
    .B(_6815__bF$buf2),
    .Y(_7669_)
);

FILL SFILL23800x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL63960x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28760x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1322_),
    .B(_1321_),
    .C(_1320_),
    .Y(_1323_)
);

OAI21X1 _22569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .B(_643_),
    .C(_645_),
    .Y(_865_)
);

FILL SFILL64120x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_30_bF$buf1),
    .Y(_405_)
);

NOR3X1 _13832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3183_),
    .B(_3181_),
    .C(_3178_),
    .Y(_3200_)
);

NAND3X1 _13412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2549_),
    .C(_2739_),
    .Y(_2740_)
);

BUFX2 _23930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[48]),
    .Y(y[48])
);

XOR2X1 _23510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1890_),
    .B(_1879_),
    .Y(_1891_)
);

NAND2X1 _14617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3535_),
    .B(_3777_),
    .Y(_4057_)
);

FILL SFILL49560x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6762_),
    .B(_6761_),
    .C(_6760_),
    .Y(_6767_)
);

FILL SFILL49160x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8706_),
    .B(_8704_),
    .Y(_8719_)
);

OAI21X1 _18450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8257_),
    .B(_8258_),
    .C(_8225_),
    .Y(_8259_)
);

NAND2X1 _18030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7796_),
    .B(_7797_),
    .Y(_7798_)
);

FILL SFILL54120x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _20635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10314_),
    .B(_10315_),
    .C(_10313_),
    .Y(_10655_)
);

AOI21X1 _20215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10187_),
    .B(_10188_),
    .C(_10186_),
    .Y(_10194_)
);

NAND3X1 _19655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9574_),
    .B(_9573_),
    .C(_9482_),
    .Y(_9581_)
);

NAND3X1 _19235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9113_),
    .B(_9116_),
    .C(_9114_),
    .Y(_9120_)
);

AOI22X1 _14790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_22_bF$buf1),
    .C(breg_1_bF$buf2),
    .D(areg_21_bF$buf1),
    .Y(_4247_)
);

INVX1 _14370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3785_),
    .Y(_3786_)
);

FILL SFILL59240x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5196_),
    .B(_5200_),
    .C(_5204_),
    .Y(_5568_)
);

XOR2X1 _15575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5055_),
    .B(_5106_),
    .Y(_5107_)
);

NAND3X1 _15155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3509_),
    .B(_3515_),
    .C(_4641_),
    .Y(_4647_)
);

FILL SFILL33560x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11699_),
    .B(_11698_),
    .C(_11697_),
    .Y(_11704_)
);

INVX1 _21173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11244_),
    .Y(_11245_)
);

OAI21X1 _17721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_4551__bF$buf1),
    .C(_7446_),
    .Y(_7460_)
);

OAI21X1 _17301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6995_),
    .B(_6994_),
    .C(_6959_),
    .Y(_7000_)
);

OAI21X1 _22798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(_1113_),
    .C(_1114_),
    .Y(_1115_)
);

OR2X2 _22378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_640_),
    .Y(_656_)
);

XNOR2X1 _18926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8776_),
    .B(_8780_),
    .Y(_8781_)
);

AOI21X1 _18506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7938_),
    .B(_7941_),
    .C(_7943_),
    .Y(_8321_)
);

NAND2X1 _13641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_18_bF$buf5),
    .Y(_2990_)
);

NAND3X1 _13221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2528_),
    .C(_2529_),
    .Y(_2531_)
);

FILL SFILL69160x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4301_),
    .B(_4308_),
    .C(_4065_),
    .Y(_4309_)
);

NAND2X1 _14426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3805_),
    .B(_3802_),
    .Y(_3849_)
);

INVX1 _14006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3130_),
    .Y(_3389_)
);

FILL SFILL8920x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10889_),
    .B(_10894_),
    .C(_10901_),
    .Y(_10906_)
);

OAI21X1 _20444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10439_),
    .B(_10440_),
    .C(_10392_),
    .Y(_10445_)
);

NOR3X1 _20024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9971_),
    .B(_9974_),
    .C(_9977_),
    .Y(_9984_)
);

NAND3X1 _19884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9779_),
    .B(_9772_),
    .C(_9777_),
    .Y(_9832_)
);

NAND2X1 _19464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9316_),
    .B(_9313_),
    .Y(_9371_)
);

OAI21X1 _19044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8909_),
    .B(_8908_),
    .C(_8899_),
    .Y(_8910_)
);

FILL SFILL59160x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11754_),
    .B(_11764_),
    .C(_11762_),
    .Y(_11765_)
);

NAND3X1 _21229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11304_),
    .B(_11305_),
    .C(_11303_),
    .Y(_11306_)
);

NAND2X1 _12912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_34_),
    .B(_78_),
    .Y(_1434_)
);

NAND3X1 _15384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4892_),
    .B(_4898_),
    .C(_4812_),
    .Y(_4899_)
);

FILL FILL74120x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5961_),
    .B(_5967_),
    .C(_5886_),
    .Y(_6218_)
);

OAI21X1 _16169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf2),
    .B(_3529__bF$buf1),
    .C(_5757_),
    .Y(_5758_)
);

FILL FILL74040x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18760x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7276_),
    .B(_7277_),
    .C(_7284_),
    .Y(_7710_)
);

OAI21X1 _17530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_6050__bF$buf2),
    .C(_7238_),
    .Y(_7249_)
);

NAND3X1 _17110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6771_),
    .B(_6781_),
    .C(_6777_),
    .Y(_6790_)
);

FILL SFILL54120x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .B(_4270_),
    .Y(_4325_)
);

NAND2X1 _22187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_444_),
    .Y(_447_)
);

OAI21X1 _18735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8569_),
    .B(_8570_),
    .C(_8568_),
    .Y(_8571_)
);

AOI21X1 _18315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8110_),
    .B(_8107_),
    .C(_8082_),
    .Y(_8111_)
);

INVX1 _13870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3239_),
    .Y(_3240_)
);

XNOR2X1 _13450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2779_),
    .B(_2778_),
    .Y(_2780_)
);

NAND3X1 _13030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2312_),
    .B(_2316_),
    .C(_2318_),
    .Y(_2325_)
);

OAI21X1 _14655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3818_),
    .B(_3826_),
    .C(_3814_),
    .Y(_4099_)
);

INVX1 _14235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3365_),
    .Y(_3640_)
);

AOI21X1 _20673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10620_),
    .B(_10619_),
    .C(_10461_),
    .Y(_10696_)
);

AOI21X1 _20253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10223_),
    .B(_10220_),
    .C(_10217_),
    .Y(_10236_)
);

NAND3X1 _16801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6445_),
    .B(_6449_),
    .C(_6448_),
    .Y(_6451_)
);

OAI21X1 _19693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9618_),
    .B(_9622_),
    .C(_9267_),
    .Y(_9623_)
);

AOI21X1 _19273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9150_),
    .B(_9147_),
    .C(_9145_),
    .Y(_9162_)
);

NOR3X1 _21878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_106_),
    .C(_107_),
    .Y(_108_)
);

AOI21X1 _21458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11555_),
    .B(_11556_),
    .C(_11554_),
    .Y(_11557_)
);

OAI21X1 _21038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11092_),
    .B(_11093_),
    .C(_11095_),
    .Y(_11096_)
);

FILL SFILL69240x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10375_),
    .B(_10408_),
    .Y(_11253_)
);

NAND3X1 _12301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6428_),
    .B(_6560_),
    .C(_6637_),
    .Y(_6658_)
);

NAND2X1 _15193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_18_bF$buf4),
    .Y(_4689_)
);

AOI21X1 _13926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3091_),
    .B(_3089_),
    .C(_3301_),
    .Y(_3302_)
);

NAND2X1 _13506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2630_),
    .B(_2640_),
    .Y(_2842_)
);

NAND2X1 _23604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1993_),
    .B(_1986_),
    .Y(_1994_)
);

NAND3X1 _16398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6007_),
    .B(_6006_),
    .C(_6008_),
    .Y(_6009_)
);

FILL SFILL59240x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8822_),
    .B(_8821_),
    .C(_8740_),
    .Y(_8823_)
);

INVX2 _18544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8362_),
    .Y(_8363_)
);

NAND3X1 _18124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7895_),
    .B(_7897_),
    .C(_7896_),
    .Y(_7902_)
);

FILL SFILL24040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10114_),
    .B(_10755_),
    .C(_10756_),
    .D(_10464_),
    .Y(_10757_)
);

NAND3X1 _20309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10296_),
    .B(_10295_),
    .C(_10294_),
    .Y(_10297_)
);

FILL FILL74200x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9680_),
    .B(_9679_),
    .C(_9678_),
    .Y(_9683_)
);

NAND3X1 _19329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9216_),
    .B(_9004_),
    .C(_9217_),
    .Y(_9223_)
);

INVX2 _14884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4349_),
    .Y(_4350_)
);

NOR2X1 _14464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3879_),
    .B(_3877_),
    .Y(_3891_)
);

NAND2X1 _14044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3379_),
    .B(_3384_),
    .Y(_3431_)
);

FILL FILL74120x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5209_),
    .B(_5208_),
    .C(_5207_),
    .Y(_5210_)
);

NAND3X1 _15249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4734_),
    .B(_4738_),
    .C(_4740_),
    .Y(_4750_)
);

NOR2X1 _20482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10473_),
    .B(_10471_),
    .Y(_10487_)
);

NOR3X1 _20062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10025_),
    .B(_10020_),
    .C(_10023_),
    .Y(_10026_)
);

FILL SFILL18760x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6232_),
    .B(_6230_),
    .C(_6228_),
    .Y(_6241_)
);

NAND3X1 _19082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8943_),
    .B(_8947_),
    .C(_8951_),
    .Y(_8952_)
);

FILL SFILL33960x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11794_),
    .B(_11798_),
    .C(_11718_),
    .Y(_11807_)
);

AOI21X1 _21267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11024_),
    .B(_11028_),
    .C(_11031_),
    .Y(_11346_)
);

OAI21X1 _17815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7555_),
    .B(_7556_),
    .C(_7513_),
    .Y(_7563_)
);

NAND3X1 _12950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_),
    .B(_1729_),
    .C(_1805_),
    .Y(_1849_)
);

NOR2X1 _12530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9071_),
    .B(_9092_),
    .Y(_9159_)
);

NOR3X1 _12110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4500_),
    .B(_4357_),
    .C(_4511_),
    .Y(_4555_)
);

FILL SFILL69400x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23560x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3085_),
    .B(_3086_),
    .C(_3083_),
    .Y(_3093_)
);

OAI21X1 _13315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2631_),
    .C(_2632_),
    .Y(_2633_)
);

INVX1 _23833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2192_),
    .Y(_2241_)
);

NAND2X1 _23413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_1683_),
    .Y(_1786_)
);

FILL SFILL23960x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf3),
    .B(_3253__bF$buf1),
    .C(_8612_),
    .Y(_8613_)
);

AOI21X1 _18353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8143_),
    .B(_8140_),
    .C(_8124_),
    .Y(_8153_)
);

FILL SFILL69320x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13560x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10976_),
    .B(_10975_),
    .C(_10697_),
    .Y(_11008_)
);

OAI21X1 _20538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10544_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10548_)
);

AOI21X1 _20118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10086_),
    .B(_10085_),
    .C(_10078_),
    .Y(_10087_)
);

OAI21X1 _19978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9569_),
    .B(_9925_),
    .C(_9928_),
    .Y(_9934_)
);

NAND3X1 _19558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9472_),
    .B(_9473_),
    .C(_9471_),
    .Y(_9474_)
);

XNOR2X1 _19138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9012_),
    .B(_9008_),
    .Y(_9013_)
);

NAND3X1 _14693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4140_),
    .B(_4134_),
    .C(_4139_),
    .Y(_4141_)
);

AOI22X1 _14273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_20_bF$buf3),
    .C(breg_1_bF$buf2),
    .D(areg_19_bF$buf2),
    .Y(_3682_)
);

NAND2X1 _15898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5460_),
    .B(_5456_),
    .Y(_5461_)
);

NAND2X1 _15478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4996_),
    .B(_4991_),
    .Y(_5000_)
);

INVX8 _15058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf4),
    .Y(_4541_)
);

FILL SFILL59320x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10198_),
    .B(_10193_),
    .C(_10201_),
    .Y(_10278_)
);

INVX1 _21496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11597_),
    .Y(_11598_)
);

XNOR2X1 _21076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11137_),
    .B(_11134_),
    .Y(_11138_)
);

NAND2X1 _17624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_20_bF$buf0),
    .Y(_7353_)
);

NAND3X1 _17204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6891_),
    .B(_6892_),
    .C(_6890_),
    .Y(_6893_)
);

AOI21X1 _18829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8667_),
    .B(_8673_),
    .C(_8635_),
    .Y(_8674_)
);

OAI21X1 _18409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8213_),
    .B(_8212_),
    .C(_8197_),
    .Y(_8214_)
);

FILL FILL74200x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3341_),
    .B(_3342_),
    .C(_3340_),
    .Y(_3343_)
);

INVX8 _13544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf5),
    .Y(_2884_)
);

NOR2X1 _13124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_2012_),
    .Y(_2424_)
);

INVX1 _23642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2035_),
    .Y(_2036_)
);

OAI21X1 _23222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1443_),
    .C(_1450_),
    .Y(_1577_)
);

OAI21X1 _14749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3946_),
    .B(_4201_),
    .C(_3994_),
    .Y(_4202_)
);

OAI21X1 _14329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3736_),
    .B(_3742_),
    .C(_3522_),
    .Y(_3743_)
);

DFFPOSX1 _24007_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[61]),
    .CLK(clk_bF$buf9),
    .D(_0_[61])
);

NAND2X1 _18582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8403_),
    .B(_8401_),
    .Y(_8404_)
);

NAND3X1 _18162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7938_),
    .B(_7941_),
    .C(_7943_),
    .Y(_7944_)
);

OAI21X1 _20767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10553_),
    .B(_10550_),
    .C(_10543_),
    .Y(_10799_)
);

AOI21X1 _20347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10305_),
    .B(_10309_),
    .C(_9995_),
    .Y(_10338_)
);

NOR3X1 _19787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9720_),
    .B(_9719_),
    .C(_9721_),
    .Y(_9725_)
);

NAND2X1 _19367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9256_),
    .B(_8470_),
    .Y(_9264_)
);

AOI21X1 _14082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3457_),
    .B(_3451_),
    .C(_3309_),
    .Y(_3473_)
);

NAND3X1 _12815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_373_),
    .C(_352_),
    .Y(_374_)
);

OAI21X1 _22913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1233_),
    .C(_1235_),
    .Y(_1242_)
);

OAI21X1 _15287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4790_),
    .B(_4791_),
    .C(_4789_),
    .Y(_4792_)
);

FILL SFILL74280x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7336_),
    .B(_7329_),
    .C(_7334_),
    .Y(_7605_)
);

NAND2X1 _17433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7143_),
    .B(_7144_),
    .Y(_7145_)
);

NAND2X1 _17013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_26_bF$buf1),
    .Y(_6684_)
);

NAND3X1 _18638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7654_),
    .B(_8061_),
    .C(_8065_),
    .Y(_8464_)
);

OAI21X1 _18218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7998_),
    .B(_8004_),
    .C(_7880_),
    .Y(_8005_)
);

NAND3X1 _13773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3129_),
    .B(_3133_),
    .C(_3132_),
    .Y(_3134_)
);

NAND3X1 _13353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2674_),
    .B(_2671_),
    .C(_2662_),
    .Y(_2675_)
);

INVX1 _23871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2277_),
    .Y(_2281_)
);

NAND2X1 _23451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1826_),
    .Y(_1828_)
);

NAND3X1 _23031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1364_),
    .C(_1368_),
    .Y(_1370_)
);

FILL SFILL64280x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _14978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4452_),
    .B(_4449_),
    .Y(_4453_)
);

NAND3X1 _14558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3987_),
    .B(_3988_),
    .C(_3948_),
    .Y(_3994_)
);

NOR2X1 _14138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .B(_3532_),
    .Y(_3533_)
);

FILL SFILL64200x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _18391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8193_),
    .B(_8190_),
    .Y(_8195_)
);

NOR3X1 _20996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11034_),
    .B(_11020_),
    .C(_11040_),
    .Y(_11050_)
);

NAND3X1 _20576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10556_),
    .B(_10586_),
    .C(_10589_),
    .Y(_10590_)
);

AOI21X1 _20156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10128_),
    .B(_10127_),
    .C(_10126_),
    .Y(_10129_)
);

NAND2X1 _16704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6343_),
    .B(_6344_),
    .Y(_6345_)
);

OAI21X1 _19596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9179_),
    .B(_9143_),
    .C(_9169_),
    .Y(_9516_)
);

AOI21X1 _19176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8697_),
    .B(_9054_),
    .C(_9053_),
    .Y(_9055_)
);

NOR2X1 _17909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_7225__bF$buf1),
    .Y(_7665_)
);

NOR2X1 _12624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10090_),
    .B(_10156_),
    .Y(_10189_)
);

NAND2X1 _12204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5574_),
    .B(_5563_),
    .Y(_5585_)
);

INVX1 _22722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .Y(_1033_)
);

OAI21X1 _22302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_372_),
    .C(_395_),
    .Y(_573_)
);

OAI21X1 _15096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4581_),
    .B(_4582_),
    .C(_4580_),
    .Y(_4583_)
);

NOR3X1 _13829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2921_),
    .C(_2920_),
    .Y(_3196_)
);

AOI21X1 _13409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2730_),
    .B(_2731_),
    .C(_2553_),
    .Y(_2736_)
);

BUFX2 _23927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[45]),
    .Y(y[45])
);

OAI21X1 _23507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(_1886_),
    .C(_1887_),
    .Y(_1888_)
);

NAND3X1 _17662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7388_),
    .B(_7391_),
    .C(_7394_),
    .Y(_7395_)
);

NAND2X1 _17242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_18_bF$buf2),
    .Y(_6935_)
);

NAND3X1 _18867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8710_),
    .B(_8712_),
    .C(_8711_),
    .Y(_8716_)
);

NAND3X1 _18447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8250_),
    .B(_8251_),
    .C(_8252_),
    .Y(_8256_)
);

INVX2 _18027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7794_),
    .Y(_7795_)
);

NAND3X1 _13582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2820_),
    .B(_2824_),
    .C(_2832_),
    .Y(_2926_)
);

OAI21X1 _13162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_2465__bF$buf2),
    .C(_2294_),
    .Y(_2466_)
);

NOR2X1 _23680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .B(_2073_),
    .Y(_2076_)
);

XOR2X1 _23260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1618_),
    .Y(_1619_)
);

FILL SFILL44120x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4243_),
    .Y(_4244_)
);

INVX2 _14367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3782_),
    .Y(_3783_)
);

DFFPOSX1 _24045_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[3]),
    .CLK(clk_bF$buf8),
    .D(b[3])
);

FILL SFILL74280x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10354_),
    .B(_10378_),
    .C(_10379_),
    .Y(_10380_)
);

AND2X2 _16933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6200_),
    .B(_6192_),
    .Y(_6596_)
);

XOR2X1 _16513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6070_),
    .B(_6134_),
    .Y(_6135_)
);

FILL SFILL74200x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7451_),
    .B(_7443_),
    .C(_7455_),
    .Y(_7456_)
);

FILL SFILL44040x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_735_),
    .C(_779_),
    .Y(_790_)
);

OAI21X1 _12433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8052_),
    .B(_8063_),
    .C(_7294_),
    .Y(_8095_)
);

XOR2X1 _22951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1274_),
    .Y(_1283_)
);

OAI21X1 _12013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2946_),
    .B(_2901_),
    .C(_3482_),
    .Y(_3493_)
);

NAND2X1 _22531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_765_),
    .Y(_824_)
);

OAI21X1 _22111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_357_),
    .C(_354_),
    .Y(_363_)
);

FILL SFILL64280x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2933_),
    .B(_2925_),
    .C(_2793_),
    .Y(_2986_)
);

NAND3X1 _13218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2358_),
    .B(_2523_),
    .C(_2526_),
    .Y(_2527_)
);

NAND2X1 _23736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_29_bF$buf0),
    .B(breg_29_bF$buf3),
    .Y(_2137_)
);

OAI21X1 _23316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686__bF$buf0),
    .B(_5668__bF$buf1),
    .C(_1564_),
    .Y(_1680_)
);

NOR2X1 _17891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7214_),
    .B(_7638_),
    .Y(_7646_)
);

NAND3X1 _17471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6814_),
    .B(_6916_),
    .C(_6917_),
    .Y(_7186_)
);

AOI21X1 _17051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6708_),
    .B(_6715_),
    .C(_6693_),
    .Y(_6726_)
);

OAI21X1 _18676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf1),
    .B(_5668__bF$buf3),
    .C(_8493_),
    .Y(_8506_)
);

AOI21X1 _18256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7221_),
    .B(_7616_),
    .C(_8046_),
    .Y(_8047_)
);

OAI21X1 _13391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_2715_),
    .C(_2713_),
    .Y(_2717_)
);

AOI21X1 _21802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11671_),
    .B(_11675_),
    .C(_11677_),
    .Y(_25_)
);

FILL SFILL54200x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4031_),
    .B(_4035_),
    .C(_3775_),
    .Y(_4036_)
);

NAND3X1 _14176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3560_),
    .B(_3565_),
    .C(_3567_),
    .Y(_3575_)
);

FILL SFILL39000x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1282_),
    .B(_1228_),
    .C(_1391_),
    .Y(_1401_)
);

AOI21X1 _20194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10152_),
    .B(_10155_),
    .C(_10159_),
    .Y(_10171_)
);

NAND3X1 _16742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6116_),
    .B(_6048_),
    .C(_6120_),
    .Y(_6387_)
);

OAI21X1 _16322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5926_),
    .B(_5924_),
    .C(_5916_),
    .Y(_5927_)
);

AND2X2 _21399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11181_),
    .B(_11230_),
    .Y(_11492_)
);

AOI21X1 _17947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7295_),
    .B(_7299_),
    .C(_7301_),
    .Y(_7707_)
);

OAI21X1 _17527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7245_),
    .B(_7244_),
    .C(_7235_),
    .Y(_7246_)
);

NAND3X1 _17107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6786_),
    .B(_6421_),
    .C(_6778_),
    .Y(_6787_)
);

INVX1 _12662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9005_),
    .Y(_10606_)
);

NAND3X1 _12242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5815_),
    .B(_5793_),
    .C(_5760_),
    .Y(_6001_)
);

AOI21X1 _22760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1073_),
    .B(_1069_),
    .C(_949_),
    .Y(_1074_)
);

NAND2X1 _22340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_612_),
    .Y(_614_)
);

NAND2X1 _13867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3234_),
    .B(_3237_),
    .Y(_3238_)
);

DFFPOSX1 _23965_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[19]),
    .CLK(clk_bF$buf0),
    .D(_0_[19])
);

INVX1 _13447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2776_),
    .Y(_2777_)
);

NAND3X1 _13027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1881_),
    .B(_2317_),
    .C(_2321_),
    .Y(_2322_)
);

OAI21X1 _23545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1928_),
    .B(_1929_),
    .C(_1873_),
    .Y(_1930_)
);

NAND2X1 _23125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1462_),
    .B(_1455_),
    .Y(_1472_)
);

FILL SFILL8600x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _17280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6223_),
    .B(_6606_),
    .C(_6631_),
    .D(_6975_),
    .Y(_6976_)
);

FILL SFILL13640x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8294_),
    .B(_8291_),
    .Y(_8298_)
);

AOI21X1 _18065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7826_),
    .B(_7824_),
    .C(_7822_),
    .Y(_7837_)
);

NAND2X1 _11933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2616_),
    .B(_2497_),
    .Y(_2617_)
);

AND2X2 _21611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11442_),
    .B(_11721_),
    .Y(_11724_)
);

FILL SFILL38840x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10693_),
    .B(_11055_),
    .C(_11121_),
    .Y(_11220_)
);

OAI21X1 _22816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_791_),
    .C(_994_),
    .Y(_1135_)
);

AOI21X1 _16971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6635_),
    .B(_6630_),
    .C(_6636_),
    .Y(_6638_)
);

NAND2X1 _16551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_15_bF$buf2),
    .Y(_6177_)
);

NAND3X1 _16131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5714_),
    .B(_5713_),
    .C(_5715_),
    .Y(_5717_)
);

FILL SFILL28840x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7488_),
    .B(_7496_),
    .C(_7497_),
    .Y(_7498_)
);

NAND3X1 _17336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7033_),
    .B(_7024_),
    .C(_7037_),
    .Y(_7038_)
);

NAND2X1 _12891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1151_),
    .B(_1195_),
    .Y(_1206_)
);

NAND2X1 _12471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7250_),
    .B(_7261_),
    .Y(_8511_)
);

OAI21X1 _12051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3854_),
    .C(_3383_),
    .Y(_3909_)
);

NOR3X1 _13676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3021_),
    .B(_3023_),
    .C(_3027_),
    .Y(_3028_)
);

NOR2X1 _13256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2565_),
    .Y(_2568_)
);

OAI22X1 _23774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2139_),
    .C(_2141_),
    .D(_2137_),
    .Y(_2178_)
);

NAND2X1 _23354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1693_),
    .B(_1721_),
    .Y(_1722_)
);

NOR3X1 _19902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9830_),
    .B(_9838_),
    .C(_9841_),
    .Y(_9852_)
);

XNOR2X1 _15822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5377_),
    .B(_5371_),
    .Y(_5378_)
);

NAND2X1 _15402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4916_),
    .B(_4918_),
    .Y(_4919_)
);

INVX2 _18294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8087_),
    .Y(_8088_)
);

FILL SFILL44200x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10910_),
    .B(_10939_),
    .C(_10943_),
    .Y(_10944_)
);

NAND3X1 _20479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10477_),
    .B(_10479_),
    .C(_10478_),
    .Y(_10483_)
);

OAI21X1 _20059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf0),
    .B(_5668__bF$buf4),
    .C(_10009_),
    .Y(_10022_)
);

NAND3X1 _16607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6233_),
    .B(_6237_),
    .C(_6226_),
    .Y(_6238_)
);

OAI21X1 _21840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_59_),
    .C(_55_),
    .Y(_66_)
);

NAND3X1 _21420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11501_),
    .B(_11506_),
    .C(_11471_),
    .Y(_11515_)
);

NAND3X1 _21000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11018_),
    .B(_11046_),
    .C(_11041_),
    .Y(_11054_)
);

NOR2X1 _19499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9023_),
    .B(_9408_),
    .Y(_9409_)
);

NAND2X1 _19079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_22_bF$buf0),
    .Y(_8948_)
);

FILL SFILL48920x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1772_),
    .B(_1783_),
    .C(_1805_),
    .Y(_1816_)
);

NAND3X1 _12527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9060_),
    .B(_9115_),
    .C(_9103_),
    .Y(_9126_)
);

OAI21X1 _22625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9976_),
    .B(_9618_),
    .C(_925_),
    .Y(_926_)
);

OAI21X1 _12107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4511_),
    .B(_4500_),
    .C(_4357_),
    .Y(_4522_)
);

NOR2X1 _22205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_466_),
    .Y(_467_)
);

INVX4 _16780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_29_bF$buf1),
    .Y(_6427_)
);

NAND3X1 _16360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5961_),
    .B(_5967_),
    .C(_5886_),
    .Y(_5968_)
);

BUFX2 BUFX2_insert440 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf4)
);

BUFX2 BUFX2_insert441 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf3)
);

BUFX2 BUFX2_insert442 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf2)
);

BUFX2 BUFX2_insert443 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf1)
);

OAI21X1 _17985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7747_),
    .B(_7748_),
    .C(_7746_),
    .Y(_7749_)
);

BUFX2 BUFX2_insert444 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf0)
);

NAND3X1 _17565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7280_),
    .B(_7285_),
    .C(_7287_),
    .Y(_7288_)
);

BUFX2 BUFX2_insert445 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[26]),
    .Y(breg_26_bF$buf4)
);

INVX2 _17145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6820_),
    .Y(_6828_)
);

BUFX2 BUFX2_insert446 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[26]),
    .Y(breg_26_bF$buf3)
);

BUFX2 BUFX2_insert447 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[26]),
    .Y(breg_26_bF$buf2)
);

BUFX2 BUFX2_insert448 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[26]),
    .Y(breg_26_bF$buf1)
);

BUFX2 BUFX2_insert449 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[26]),
    .Y(breg_26_bF$buf0)
);

NOR2X1 _12280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6396_),
    .B(_6407_),
    .Y(_6417_)
);

FILL SFILL38920x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2813_),
    .B(_2818_),
    .C(_2804_),
    .Y(_2819_)
);

NAND2X1 _13065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11723_),
    .B(_1445_),
    .Y(_2359_)
);

OAI21X1 _23583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1966_),
    .B(_1970_),
    .C(_7650_),
    .Y(_1971_)
);

NAND3X1 _23163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1513_),
    .C(_1510_),
    .Y(_1514_)
);

FILL SFILL3560x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _19711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9640_),
    .Y(_9642_)
);

AOI21X1 _15631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5159_),
    .B(_5158_),
    .C(_5154_),
    .Y(_5169_)
);

AND2X2 _15211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4703_),
    .B(_4707_),
    .Y(_4709_)
);

FILL SFILL28840x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10273_),
    .B(_10272_),
    .Y(_10274_)
);

FILL SFILL18920x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6441_),
    .B(_6479_),
    .C(_6474_),
    .Y(_6489_)
);

NAND3X1 _16416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6021_),
    .B(_6028_),
    .C(_5664_),
    .Y(_6029_)
);

OAI21X1 _11971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3022_),
    .B(_3011_),
    .C(_2420_),
    .Y(_3033_)
);

NAND2X1 _12756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11582_),
    .B(_11625_),
    .Y(_11636_)
);

NAND3X1 _12336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6911_),
    .B(_6944_),
    .C(_6966_),
    .Y(_7032_)
);

NAND3X1 _22854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1167_),
    .B(_1160_),
    .C(_1165_),
    .Y(_1177_)
);

INVX1 _22434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .Y(_717_)
);

OAI21X1 _22014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11907_),
    .B(_11896_),
    .C(_11901_),
    .Y(_257_)
);

FILL SFILL63880x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18840x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _23639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .B(areg_31_bF$buf4),
    .C(breg_26_bF$buf1),
    .D(areg_30_bF$buf4),
    .Y(_2032_)
);

NAND3X1 _23219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1446_),
    .B(_1450_),
    .C(_1453_),
    .Y(_1574_)
);

NAND2X1 _14902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_20_bF$buf2),
    .Y(_4370_)
);

NAND3X1 _17794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7529_),
    .B(_7537_),
    .C(_7539_),
    .Y(_7540_)
);

AOI21X1 _17374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7074_),
    .B(_7075_),
    .C(_7067_),
    .Y(_7080_)
);

FILL SFILL74360x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10966_),
    .B(_10965_),
    .Y(_10967_)
);

FILL SFILL53880x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10501_),
    .B(_10505_),
    .C(_10504_),
    .Y(_10506_)
);

NAND3X1 _18999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8479_),
    .B(_8855_),
    .C(_8856_),
    .Y(_8861_)
);

AOI21X1 _18579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8392_),
    .B(_8399_),
    .C(_8330_),
    .Y(_8400_)
);

OAI21X1 _18159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_7934_),
    .Y(_7940_)
);

NAND3X1 _13294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2606_),
    .B(_2607_),
    .C(_2608_),
    .Y(_2609_)
);

OAI21X1 _23392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1649_),
    .B(_1550_),
    .C(_1641_),
    .Y(_1764_)
);

AOI21X1 _19940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9876_),
    .B(_9882_),
    .C(_9860_),
    .Y(_9893_)
);

NAND2X1 _19520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_20_bF$buf0),
    .Y(_9432_)
);

AOI21X1 _19100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8633_),
    .B(_8630_),
    .C(_8970_),
    .Y(_8971_)
);

AOI21X1 _21705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11826_),
    .B(_11821_),
    .C(_11716_),
    .Y(_11827_)
);

INVX1 _14499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3670_),
    .Y(_3929_)
);

OAI21X1 _14079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3455_),
    .B(_3456_),
    .C(_3310_),
    .Y(_3469_)
);

NAND2X1 _15860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_13_bF$buf2),
    .Y(_5419_)
);

NAND3X1 _15440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4629_),
    .B(_4958_),
    .C(_4959_),
    .Y(_4960_)
);

OAI21X1 _15020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4203_),
    .B(_4498_),
    .C(_4213_),
    .Y(_4499_)
);

FILL SFILL3640x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10061_),
    .B(_10060_),
    .C(_10063_),
    .Y(_10064_)
);

INVX1 _16645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6279_),
    .Y(_6280_)
);

OAI21X1 _16225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5814_),
    .B(_5816_),
    .C(_5780_),
    .Y(_5820_)
);

FILL SFILL59080x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69320x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_527_),
    .Y(_2228_)
);

NOR3X1 _12565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8052_),
    .B(_8063_),
    .C(_8029_),
    .Y(_9543_)
);

NAND2X1 _12145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4917_),
    .B(_4906_),
    .Y(_4939_)
);

NAND2X1 _22663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_967_),
    .B(_962_),
    .Y(_968_)
);

OAI21X1 _22243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_258_),
    .C(_262_),
    .Y(_508_)
);

XNOR2X1 _23868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2277_),
    .Y(_0_[62])
);

NAND2X1 _23448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1823_),
    .Y(_1824_)
);

AOI21X1 _23028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1339_),
    .C(_1268_),
    .Y(_1366_)
);

XOR2X1 _14711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4158_),
    .B(_4159_),
    .Y(_4161_)
);

NOR2X1 _17183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6455_),
    .B(_6514_),
    .Y(_6870_)
);

NAND2X1 _15916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_17_bF$buf4),
    .Y(_5481_)
);

NAND2X1 _18388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_22_bF$buf0),
    .Y(_8191_)
);

AOI21X1 _21934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_168_),
    .B(_169_),
    .C(_167_),
    .Y(_170_)
);

OAI21X1 _21514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_11617_),
    .Y(_11618_)
);

NAND3X1 _22719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_1022_),
    .C(_1017_),
    .Y(_1029_)
);

AOI21X1 _16874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6146_),
    .B(_6148_),
    .C(_6140_),
    .Y(_6531_)
);

NAND3X1 _16454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6060_),
    .B(_6067_),
    .C(_6068_),
    .Y(_6069_)
);

AOI21X1 _16034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5592_),
    .B(_5598_),
    .C(_5511_),
    .Y(_5611_)
);

FILL SFILL53960x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7381_),
    .B(_7389_),
    .C(_7390_),
    .Y(_7391_)
);

XNOR2X1 _17239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6930_),
    .B(_6926_),
    .Y(_6931_)
);

OAI21X1 _12794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10693_),
    .B(_11055_),
    .C(_11165_),
    .Y(_144_)
);

NAND3X1 _12374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7327_),
    .B(_7349_),
    .C(_7437_),
    .Y(_7448_)
);

NAND2X1 _22892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_1218_),
    .Y(_1219_)
);

NAND3X1 _22472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_749_),
    .C(_751_),
    .Y(_759_)
);

NAND2X1 _22052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf3),
    .B(breg_26_bF$buf0),
    .Y(_299_)
);

NOR3X1 _18600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7998_),
    .B(_8004_),
    .C(_8007_),
    .Y(_8423_)
);

NOR3X1 _13999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3376_),
    .B(_3377_),
    .C(_3375_),
    .Y(_3381_)
);

NOR3X1 _13579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2868_),
    .B(_2900_),
    .C(_2908_),
    .Y(_2922_)
);

NOR2X1 _13159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2294_),
    .B(_2461_),
    .Y(_2462_)
);

NOR2X1 _23677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2013_),
    .B(_2072_),
    .Y(_2073_)
);

NAND3X1 _23257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1613_),
    .B(_1614_),
    .C(_1615_),
    .Y(_1616_)
);

FILL SFILL3720x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9735_),
    .B(_9728_),
    .C(_9687_),
    .Y(_9745_)
);

AOI21X1 _14940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4398_),
    .B(_4396_),
    .C(_4393_),
    .Y(_4411_)
);

AOI22X1 _14520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_18_bF$buf4),
    .C(breg_4_bF$buf4),
    .D(areg_17_bF$buf1),
    .Y(_3952_)
);

NAND3X1 _14100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3232_),
    .C(_2981_),
    .Y(_3492_)
);

FILL SFILL3640x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4673_),
    .B(_4931_),
    .C(_5271_),
    .Y(_5272_)
);

NAND2X1 _15305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4811_),
    .B(_4806_),
    .Y(_4812_)
);

FILL SFILL59080x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7974_),
    .B(_7976_),
    .C(_7977_),
    .Y(_7982_)
);

NAND2X1 _21743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11590_),
    .B(_11865_),
    .Y(_11868_)
);

AOI21X1 _21323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11393_),
    .B(_11398_),
    .C(_11399_),
    .Y(_11409_)
);

NAND2X1 _22948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_29_bF$buf1),
    .Y(_1279_)
);

AOI21X1 _22528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_802_),
    .C(_773_),
    .Y(_820_)
);

NAND3X1 _22108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_355_),
    .C(_359_),
    .Y(_360_)
);

NAND3X1 _16683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6307_),
    .B(_6321_),
    .C(_6316_),
    .Y(_6322_)
);

OAI21X1 _16263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_3146__bF$buf2),
    .C(_5476_),
    .Y(_5862_)
);

FILL SFILL49000x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7629_),
    .B(_7632_),
    .C(_7218_),
    .Y(_7642_)
);

FILL SFILL18840x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7180_),
    .B(_7181_),
    .C(_7179_),
    .Y(_7182_)
);

NOR3X1 _17048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6326_),
    .B(_6323_),
    .C(_6327_),
    .Y(_6722_)
);

FILL SFILL18760x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .B(_4522_),
    .C(_4555_),
    .Y(_5354_)
);

NAND2X1 _22281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_548_),
    .Y(_550_)
);

FILL SFILL23880x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2422_),
    .B(_2500_),
    .C(_2712_),
    .Y(_2713_)
);

NOR2X1 _23486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1775_),
    .B(_1861_),
    .Y(_1865_)
);

NAND2X1 _23066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1340_),
    .Y(_1407_)
);

NAND2X1 _19614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9146_),
    .B(_9535_),
    .Y(_9536_)
);

FILL SFILL39000x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5516_),
    .Y(_5523_)
);

NOR2X1 _15534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4723_),
    .B(_4771_),
    .Y(_5062_)
);

OAI21X1 _15114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4595_),
    .B(_4596_),
    .C(_4447_),
    .Y(_4603_)
);

FILL SFILL53960x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6381_),
    .B(_6382_),
    .C(_6380_),
    .Y(_6383_)
);

NAND3X1 _16319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5917_),
    .B(_5922_),
    .C(_5920_),
    .Y(_5923_)
);

OAI22X1 _21972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_207_),
    .B(_208_),
    .C(_211_),
    .D(_209_),
    .Y(_212_)
);

INVX1 _21552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11654_),
    .Y(_11659_)
);

NAND3X1 _21132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11190_),
    .B(_11177_),
    .C(_11180_),
    .Y(_11200_)
);

NAND3X1 _12659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10562_),
    .B(_10496_),
    .C(_10540_),
    .Y(_10573_)
);

AOI21X1 _12239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .B(_5936_),
    .C(_4928_),
    .Y(_5969_)
);

OAI21X1 _22757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(_1067_),
    .C(_1062_),
    .Y(_1071_)
);

FILL SFILL3720x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_25_bF$buf2),
    .Y(_611_)
);

FILL SFILL43960x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2942_),
    .B(_2943_),
    .C(_2944_),
    .Y(_2945_)
);

OAI21X1 _16492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6107_),
    .B(_6108_),
    .C(_6057_),
    .Y(_6112_)
);

OAI21X1 _16072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5652_),
    .B(_5650_),
    .C(_5647_),
    .Y(_5653_)
);

NAND3X1 _14805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4254_),
    .B(_4252_),
    .C(_4249_),
    .Y(_4264_)
);

NAND3X1 _17697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7430_),
    .B(_7432_),
    .C(_7431_),
    .Y(_7433_)
);

OAI21X1 _17277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6972_),
    .B(_6971_),
    .C(_6961_),
    .Y(_6973_)
);

NAND3X1 _22090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_295_),
    .C(_339_),
    .Y(_340_)
);

NAND2X1 _20823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf3),
    .B(areg_25_bF$buf3),
    .Y(_10861_)
);

AND2X2 _20403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10396_),
    .B(_10398_),
    .Y(_10400_)
);

NAND3X1 _13197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2494_),
    .B(_2488_),
    .C(_2496_),
    .Y(_2504_)
);

AOI21X1 _23295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1643_),
    .C(_1648_),
    .Y(_1657_)
);

NOR3X1 _19843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9779_),
    .B(_9781_),
    .C(_9780_),
    .Y(_9787_)
);

NOR2X1 _19423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9324_),
    .B(_9325_),
    .Y(_9326_)
);

NAND3X1 _19003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8861_),
    .B(_8477_),
    .C(_8862_),
    .Y(_8866_)
);

INVX2 _21608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11719_),
    .Y(_11720_)
);

AND2X2 _15763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_24_bF$buf1),
    .Y(_5313_)
);

OAI21X1 _15343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4547_),
    .B(_4537_),
    .C(_4540_),
    .Y(_4854_)
);

NAND3X1 _16968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6623_),
    .B(_6617_),
    .C(_6621_),
    .Y(_6634_)
);

OAI21X1 _16548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf0),
    .B(_2560__bF$buf3),
    .C(_6169_),
    .Y(_6173_)
);

INVX2 _16128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5673_),
    .Y(_5713_)
);

AOI21X1 _21781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11904_),
    .B(_11908_),
    .C(_11895_),
    .Y(_2_)
);

FILL SFILL23880x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_23_bF$buf3),
    .Y(_11451_)
);

NOR3X1 _12888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1118_),
    .B(_1129_),
    .C(_1107_),
    .Y(_1173_)
);

AOI21X1 _12468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8435_),
    .B(_8446_),
    .C(_7020_),
    .Y(_8478_)
);

INVX2 _22986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1298_),
    .Y(_1320_)
);

FILL SFILL23800x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3799_),
    .B(_3832_),
    .C(_3493_),
    .Y(_3876_)
);

NAND2X1 _22566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_861_),
    .B(_860_),
    .Y(_862_)
);

OAI21X1 _22146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_132_),
    .B(_130_),
    .C(_138_),
    .Y(_402_)
);

FILL SFILL13880x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4045_),
    .B(_4049_),
    .C(_3770_),
    .Y(_4054_)
);

FILL SFILL29000x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6756_),
    .B(_6763_),
    .C(_6511_),
    .Y(_6764_)
);

FILL SFILL13800x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5372_),
    .B(_5373_),
    .Y(_5374_)
);

OAI21X1 _20632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10636_),
    .B(_10640_),
    .C(_10643_),
    .Y(_10652_)
);

AOI21X1 _20212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9884_),
    .B(_9889_),
    .C(_9890_),
    .Y(_10191_)
);

OAI21X1 _19652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9479_),
    .B(_9478_),
    .C(_9391_),
    .Y(_9578_)
);

AOI21X1 _19232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9116_),
    .B(_9114_),
    .C(_9113_),
    .Y(_9117_)
);

NAND3X1 _21837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_62_),
    .C(_57_),
    .Y(_63_)
);

NOR3X1 _21417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11251_),
    .B(_11511_),
    .C(_11507_),
    .Y(_11512_)
);

FILL SFILL43960x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5203_),
    .B(_5564_),
    .Y(_5565_)
);

NAND2X1 _15572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4788_),
    .B(_4793_),
    .Y(_5104_)
);

NOR2X1 _15152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4342_),
    .B(_4640_),
    .Y(_4644_)
);

FILL SFILL64040x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6102_),
    .B(_6111_),
    .Y(_6424_)
);

OAI21X1 _16357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5957_),
    .B(_5959_),
    .C(_5915_),
    .Y(_5965_)
);

NAND3X1 _21590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11699_),
    .B(_11698_),
    .C(_11697_),
    .Y(_11700_)
);

NOR2X1 _21170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11240_),
    .B(_11236_),
    .Y(_11241_)
);

OAI21X1 _12697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10968_),
    .B(_10979_),
    .C(_10957_),
    .Y(_10990_)
);

FILL SFILL54440x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .B(areg_6_bF$buf4),
    .Y(_6385_)
);

OAI21X1 _22795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_959_),
    .C(_967_),
    .Y(_1112_)
);

XNOR2X1 _22375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_642_),
    .Y(_653_)
);

OAI21X1 _18923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8770_),
    .B(_7968_),
    .C(_8777_),
    .Y(_8778_)
);

OAI21X1 _18503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8310_),
    .B(_8314_),
    .C(_8317_),
    .Y(_8318_)
);

INVX2 _19708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9637_),
    .Y(_9638_)
);

OAI21X1 _14843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4298_),
    .B(_4299_),
    .C(_4154_),
    .Y(_4306_)
);

AOI21X1 _14423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3831_),
    .B(_3825_),
    .C(_3809_),
    .Y(_3846_)
);

OAI21X1 _14003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3174_),
    .B(_3139_),
    .C(_3167_),
    .Y(_3386_)
);

OAI21X1 _15628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4848_),
    .B(_4850_),
    .C(_5164_),
    .Y(_5165_)
);

OAI21X1 _15208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4700_),
    .B(_4701_),
    .C(_4685_),
    .Y(_4705_)
);

OAI21X1 _20861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10898_),
    .B(_10899_),
    .C(_10901_),
    .Y(_10903_)
);

OAI21X1 _20441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10439_),
    .B(_10440_),
    .C(_10436_),
    .Y(_10442_)
);

NAND2X1 _20021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9975_),
    .B(_9980_),
    .Y(_9982_)
);

NAND3X1 _19881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9823_),
    .B(_9824_),
    .C(_9827_),
    .Y(_9829_)
);

AOI21X1 _19461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9353_),
    .B(_9349_),
    .C(_9320_),
    .Y(_9368_)
);

NAND2X1 _19041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_8907_)
);

FILL SFILL8920x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _11968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2989_),
    .C(_2978_),
    .Y(_3000_)
);

FILL SFILL23800x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf3),
    .B(_7100__bF$buf0),
    .C(_11761_),
    .Y(_11762_)
);

AOI21X1 _21226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10690_),
    .B(_10991_),
    .C(_11302_),
    .Y(_11303_)
);

FILL FILL73960x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4890_),
    .B(_4889_),
    .C(_4888_),
    .Y(_4896_)
);

NAND3X1 _16586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6200_),
    .B(_6205_),
    .C(_6204_),
    .Y(_6215_)
);

AND2X2 _16166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_18_bF$buf0),
    .Y(_5755_)
);

NOR2X1 _12086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4160_),
    .B(_4281_),
    .Y(_4292_)
);

NAND2X1 _22184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_443_),
    .Y(_444_)
);

AND2X2 _18732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8144_),
    .B(_8140_),
    .Y(_8568_)
);

OAI21X1 _18312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8103_),
    .B(_8104_),
    .C(_8100_),
    .Y(_8108_)
);

AOI21X1 _20917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10963_),
    .B(_10958_),
    .C(_10811_),
    .Y(_10964_)
);

NOR3X1 _23389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1747_),
    .B(_1752_),
    .C(_1662_),
    .Y(_1760_)
);

OAI21X1 _19937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9559_),
    .B(_9529_),
    .C(_9551_),
    .Y(_9890_)
);

INVX1 _19517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9428_),
    .Y(_9429_)
);

NAND3X1 _14652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4092_),
    .B(_4093_),
    .C(_4095_),
    .Y(_4096_)
);

OAI21X1 _14232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3636_),
    .B(_3634_),
    .C(_3633_),
    .Y(_3637_)
);

FILL SFILL64040x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf0),
    .B(_2560__bF$buf1),
    .C(_5412_),
    .Y(_5416_)
);

NAND3X1 _15437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4956_),
    .B(_4948_),
    .C(_4649_),
    .Y(_4957_)
);

AOI21X1 _15017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(_4265_),
    .C(_4235_),
    .Y(_4496_)
);

OAI21X1 _20670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10646_),
    .B(_10346_),
    .C(_10637_),
    .Y(_10692_)
);

OAI21X1 _20250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf3),
    .B(_7520__bF$buf3),
    .C(_10219_),
    .Y(_10231_)
);

NAND3X1 _19690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9272_),
    .B(_9613_),
    .C(_9616_),
    .Y(_9619_)
);

AOI21X1 _19270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8780_),
    .B(_8774_),
    .C(_9157_),
    .Y(_9158_)
);

NAND2X1 _21875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_26_bF$buf2),
    .Y(_105_)
);

NAND2X1 _21455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11553_),
    .B(_11552_),
    .Y(_11554_)
);

AOI21X1 _21035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11075_),
    .B(_11082_),
    .C(_11060_),
    .Y(_11093_)
);

INVX2 _15190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4684_),
    .Y(_4685_)
);

AOI21X1 _13923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3292_),
    .B(_3293_),
    .C(_3256_),
    .Y(_3299_)
);

OAI21X1 _13503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2837_),
    .B(_2838_),
    .C(_2835_),
    .Y(_2839_)
);

AND2X2 _23601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1989_),
    .B(_1948_),
    .Y(_1991_)
);

NAND2X1 _16395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6004_),
    .B(_6005_),
    .Y(_6006_)
);

INVX1 _14708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4156_),
    .Y(_4157_)
);

FILL SFILL8520x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8813_),
    .B(_8818_),
    .Y(_8820_)
);

NAND2X1 _18541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8354_),
    .B(_8358_),
    .Y(_8360_)
);

AOI21X1 _18121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7897_),
    .B(_7896_),
    .C(_7895_),
    .Y(_7899_)
);

NAND3X1 _20726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10751_),
    .B(_10753_),
    .C(_10752_),
    .Y(_10754_)
);

NAND2X1 _20306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10292_),
    .B(_10293_),
    .Y(_10294_)
);

OAI21X1 _23198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(_1516_),
    .C(_1514_),
    .Y(_1551_)
);

NOR3X1 _19746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9665_),
    .B(_9650_),
    .C(_9671_),
    .Y(_9680_)
);

AOI21X1 _19326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8999_),
    .B(_9000_),
    .C(_8998_),
    .Y(_9220_)
);

AOI21X1 _14881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4320_),
    .C(_4059_),
    .Y(_4347_)
);

AOI21X1 _14461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3607_),
    .B(_3609_),
    .C(_3615_),
    .Y(_3888_)
);

AOI21X1 _14041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3418_),
    .B(_3411_),
    .C(_3395_),
    .Y(_3428_)
);

AOI21X1 _15666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4856_),
    .B(_4860_),
    .C(_4864_),
    .Y(_5207_)
);

NAND3X1 _15246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4739_),
    .B(_4746_),
    .C(_4709_),
    .Y(_4747_)
);

AOI21X1 _21684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11799_),
    .B(_11803_),
    .C(_11717_),
    .Y(_11804_)
);

NOR2X1 _21264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11336_),
    .B(_11337_),
    .Y(_11343_)
);

NAND3X1 _17812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7507_),
    .B(_7500_),
    .C(_7505_),
    .Y(_7560_)
);

FILL SFILL23800x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64280x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_1190_),
    .Y(_1215_)
);

OAI21X1 _22469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_754_),
    .C(_751_),
    .Y(_755_)
);

FILL SFILL64120x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_64_),
    .B(_294_),
    .C(_57_),
    .Y(_295_)
);

NAND3X1 _13732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3050_),
    .B(_3084_),
    .C(_3089_),
    .Y(_3090_)
);

NOR2X1 _13312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf1),
    .B(_5420__bF$buf0),
    .Y(_2630_)
);

NOR2X1 _23830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .B(_2236_),
    .Y(_2237_)
);

NOR2X1 _23410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf3),
    .B(_7225__bF$buf2),
    .Y(_1782_)
);

INVX2 _14937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4407_),
    .Y(_4408_)
);

NOR2X1 _14517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf1),
    .B(_2669__bF$buf0),
    .Y(_3949_)
);

NOR2X1 _18770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf3),
    .B(_3526_),
    .Y(_8609_)
);

OAI21X1 _18350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7812_),
    .B(_7814_),
    .C(_7806_),
    .Y(_8149_)
);

FILL SFILL54120x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11004_),
    .B(_10691_),
    .C(_10989_),
    .Y(_11005_)
);

AOI21X1 _20535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10534_),
    .B(_10527_),
    .C(_10495_),
    .Y(_10545_)
);

AOI21X1 _20115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9689_),
    .B(_9722_),
    .C(_9725_),
    .Y(_10084_)
);

OAI21X1 _19975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9852_),
    .B(_9851_),
    .C(_9757_),
    .Y(_9931_)
);

NAND3X1 _19555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9465_),
    .B(_9467_),
    .C(_9464_),
    .Y(_9471_)
);

NOR2X1 _19135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8948_),
    .B(_9009_),
    .Y(_9010_)
);

NAND3X1 _14690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4128_),
    .B(_4121_),
    .C(_4125_),
    .Y(_4137_)
);

NAND2X1 _14270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf1),
    .B(areg_18_bF$buf3),
    .Y(_3678_)
);

FILL SFILL59240x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33880x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .B(_5451_),
    .C(_5454_),
    .Y(_5458_)
);

AND2X2 _15475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4991_),
    .B(_4996_),
    .Y(_4997_)
);

INVX2 _15055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4537_),
    .Y(_4538_)
);

AOI21X1 _21493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11574_),
    .B(_11577_),
    .C(_11322_),
    .Y(_11595_)
);

NAND2X1 _21073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_22_bF$buf3),
    .Y(_11135_)
);

NOR2X1 _17621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7347_),
    .B(_7348_),
    .Y(_7350_)
);

INVX2 _17201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .Y(_6890_)
);

NOR2X1 _22698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_999_),
    .Y(_1006_)
);

INVX1 _22278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_300_),
    .Y(_546_)
);

AOI21X1 _18826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8646_),
    .B(_8649_),
    .C(_8659_),
    .Y(_8671_)
);

NAND2X1 _18406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_18_bF$buf1),
    .Y(_8211_)
);

XNOR2X1 _13961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_3312_),
    .Y(_3340_)
);

NAND2X1 _13541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_16_bF$buf0),
    .Y(_2881_)
);

NAND3X1 _13121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2416_),
    .B(_2418_),
    .C(_2417_),
    .Y(_2421_)
);

FILL SFILL38760x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4196_),
    .B(_4197_),
    .C(_4198_),
    .Y(_4199_)
);

NAND3X1 _14326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3730_),
    .B(_3733_),
    .C(_3729_),
    .Y(_3740_)
);

DFFPOSX1 _24004_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[58]),
    .CLK(clk_bF$buf9),
    .D(_0_[58])
);

FILL SFILL69080x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10790_),
    .B(_10791_),
    .C(_10741_),
    .Y(_10796_)
);

NOR2X1 _20344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10335_),
    .B(_10330_),
    .Y(_0_[38])
);

OAI21X1 _19784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9720_),
    .B(_9719_),
    .C(_9721_),
    .Y(_9722_)
);

NAND2X1 _19364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9260_),
    .B(_8878_),
    .Y(_9261_)
);

FILL SFILL28760x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_86_),
    .C(_11889_),
    .Y(_208_)
);

FILL SFILL64120x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11653_),
    .B(_11654_),
    .C(_11650_),
    .Y(_11655_)
);

OAI21X1 _21129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11194_),
    .B(_11195_),
    .C(_11193_),
    .Y(_11196_)
);

NOR2X1 _12812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_330_),
    .B(_10595_),
    .Y(_341_)
);

NAND3X1 _22910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .B(_1237_),
    .C(_1235_),
    .Y(_1238_)
);

AOI21X1 _15284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4456_),
    .B(_4461_),
    .C(_4464_),
    .Y(_4789_)
);

AOI21X1 _16489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6095_),
    .B(_6090_),
    .C(_6058_),
    .Y(_6108_)
);

NAND3X1 _16069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5635_),
    .B(_5626_),
    .C(_5633_),
    .Y(_5649_)
);

FILL SFILL49160x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7583_),
    .B(_7588_),
    .C(_7434_),
    .Y(_7601_)
);

NAND3X1 _17430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7135_),
    .B(_7091_),
    .C(_7140_),
    .Y(_7141_)
);

NAND2X1 _17010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_24_bF$buf3),
    .Y(_6680_)
);

FILL SFILL54120x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38760x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .C(_333_),
    .Y(_337_)
);

NAND3X1 _18635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8460_),
    .B(_8461_),
    .C(_8459_),
    .Y(_8462_)
);

NAND3X1 _18215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7994_),
    .B(_7995_),
    .C(_7928_),
    .Y(_8002_)
);

NAND2X1 _13770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_15_bF$buf3),
    .Y(_3130_)
);

NAND3X1 _13350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2664_),
    .B(_2670_),
    .C(_2668_),
    .Y(_2671_)
);

NAND2X1 _14975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_13_bF$buf3),
    .Y(_4450_)
);

NAND3X1 _14555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3934_),
    .B(_3939_),
    .C(_3941_),
    .Y(_3991_)
);

OAI21X1 _14135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf2),
    .B(_3529__bF$buf0),
    .C(_3251_),
    .Y(_3530_)
);

AOI21X1 _20993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11046_),
    .B(_11041_),
    .C(_11018_),
    .Y(_11047_)
);

AOI21X1 _20573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10582_),
    .B(_10583_),
    .C(_10581_),
    .Y(_10587_)
);

INVX2 _20153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10118_),
    .Y(_10126_)
);

NAND3X1 _16701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6335_),
    .B(_6340_),
    .C(_6291_),
    .Y(_6342_)
);

OAI21X1 _19593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9506_),
    .B(_9507_),
    .C(_9489_),
    .Y(_9513_)
);

NAND3X1 _19173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9043_),
    .B(_9050_),
    .C(_9051_),
    .Y(_9052_)
);

NOR2X1 _21778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11902_),
    .B(_11905_),
    .Y(_11906_)
);

NAND2X1 _21358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf4),
    .B(areg_22_bF$buf2),
    .Y(_11447_)
);

AOI21X1 _17906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7589_),
    .B(_7596_),
    .C(_7343_),
    .Y(_7662_)
);

FILL SFILL69240x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10134_),
    .B(_10123_),
    .Y(_10156_)
);

NAND3X1 _12201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5431_),
    .B(_5464_),
    .C(_5541_),
    .Y(_5552_)
);

AOI21X1 _15093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4233_),
    .B(_4272_),
    .C(_4579_),
    .Y(_4580_)
);

OAI21X1 _13826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3178_),
    .B(_3181_),
    .C(_3183_),
    .Y(_3193_)
);

NAND3X1 _13406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2729_),
    .B(_2552_),
    .C(_2732_),
    .Y(_2733_)
);

BUFX2 _23924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[42]),
    .Y(y[42])
);

NAND2X1 _23504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_26_bF$buf1),
    .B(breg_29_bF$buf2),
    .Y(_1885_)
);

OAI21X1 _16298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5551_),
    .B(_5543_),
    .C(_5547_),
    .Y(_5900_)
);

FILL SFILL23320x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8712_),
    .B(_8711_),
    .C(_8710_),
    .Y(_8713_)
);

AOI21X1 _18444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8251_),
    .B(_8252_),
    .C(_8250_),
    .Y(_8253_)
);

AOI21X1 _18024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7362_),
    .B(_7364_),
    .C(_7356_),
    .Y(_7792_)
);

NAND3X1 _20629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10644_),
    .B(_10643_),
    .C(_10647_),
    .Y(_10648_)
);

OAI21X1 _20209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10177_),
    .B(_10179_),
    .C(_10142_),
    .Y(_10187_)
);

NAND2X1 _19649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9528_),
    .B(_9568_),
    .Y(_9574_)
);

INVX2 _19229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9106_),
    .Y(_9113_)
);

XNOR2X1 _14784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4240_),
    .B(_4236_),
    .Y(_4241_)
);

NAND2X1 _14364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3566_),
    .B(_3572_),
    .Y(_3780_)
);

DFFPOSX1 _24042_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[0]),
    .CLK(clk_bF$buf9),
    .D(b[0])
);

INVX2 _15989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5560_),
    .Y(_5561_)
);

NAND3X1 _15569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5098_),
    .B(_5099_),
    .C(_5097_),
    .Y(_5100_)
);

XNOR2X1 _15149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4345_),
    .B(_4640_),
    .Y(_0_[23])
);

OAI21X1 _20382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10376_),
    .B(_10369_),
    .C(_10355_),
    .Y(_10377_)
);

FILL SFILL49160x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6221_),
    .B(_6259_),
    .C(_6256_),
    .Y(_6592_)
);

NAND2X1 _16510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_23_bF$buf0),
    .Y(_6131_)
);

FILL SFILL33960x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11645_),
    .B(_11642_),
    .Y(_11697_)
);

NOR2X1 _21167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10570_),
    .B(_11237_),
    .Y(_11238_)
);

NOR2X1 _17715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7034_),
    .B(_7452_),
    .Y(_7453_)
);

NAND3X1 _12850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .B(_571_),
    .C(_604_),
    .Y(_757_)
);

AOI21X1 _12430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7876_),
    .B(_7920_),
    .C(_7547_),
    .Y(_8063_)
);

INVX2 _12010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3449_),
    .Y(_3460_)
);

OAI21X1 _13635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2982_),
    .B(_2756_),
    .C(_2947_),
    .Y(_2983_)
);

OAI21X1 _13215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_2521_),
    .C(_2361_),
    .Y(_2524_)
);

NAND2X1 _23733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2132_),
    .B(_2133_),
    .Y(_2134_)
);

AOI21X1 _23313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1566_),
    .C(_1676_),
    .Y(_1677_)
);

FILL SFILL23960x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8497_),
    .B(_8502_),
    .C(_8490_),
    .Y(_8503_)
);

AOI21X1 _18253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8042_),
    .B(_8043_),
    .C(_7660_),
    .Y(_8044_)
);

FILL SFILL13560x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10888_),
    .B(_10882_),
    .C(_10849_),
    .Y(_10899_)
);

OAI21X1 _20438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10425_),
    .B(_10426_),
    .C(_10423_),
    .Y(_10438_)
);

NAND3X1 _20018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9637_),
    .B(_9972_),
    .C(_9973_),
    .Y(_9978_)
);

NOR3X1 _19878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9810_),
    .B(_9807_),
    .C(_9809_),
    .Y(_9825_)
);

NAND3X1 _19458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9342_),
    .B(_9347_),
    .C(_9352_),
    .Y(_9364_)
);

NAND2X1 _19038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8901_),
    .B(_8902_),
    .Y(_8903_)
);

NAND3X1 _14593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_4028_),
    .C(_4026_),
    .Y(_4033_)
);

NAND3X1 _14173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3537_),
    .B(_3566_),
    .C(_3571_),
    .Y(_3572_)
);

NOR2X1 _12906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1206_),
    .B(_1217_),
    .Y(_1369_)
);

NAND3X1 _15798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4979_),
    .B(_5342_),
    .C(_5338_),
    .Y(_5351_)
);

NAND3X1 _15378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4885_),
    .B(_4814_),
    .C(_4891_),
    .Y(_4892_)
);

NAND3X1 _20191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10144_),
    .B(_10160_),
    .C(_10166_),
    .Y(_10168_)
);

FILL SFILL59240x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11488_),
    .B(_11482_),
    .C(_11486_),
    .Y(_11489_)
);

NAND3X1 _17944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7668_),
    .B(_7695_),
    .C(_7692_),
    .Y(_7704_)
);

NAND2X1 _17524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_28_bF$buf0),
    .Y(_7243_)
);

AOI21X1 _17104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6783_),
    .B(_6782_),
    .C(_6774_),
    .Y(_6784_)
);

AOI21X1 _18729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8220_),
    .B(_8218_),
    .C(_8563_),
    .Y(_8564_)
);

AOI21X1 _18309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8092_),
    .B(_8091_),
    .C(_8088_),
    .Y(_8104_)
);

FILL FILL74200x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3223_),
    .B(_3228_),
    .C(_2958_),
    .Y(_3235_)
);

DFFPOSX1 _23962_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[16]),
    .CLK(clk_bF$buf10),
    .D(_0_[16])
);

INVX1 _13444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2773_),
    .Y(_2774_)
);

AOI21X1 _13024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2315_),
    .C(_2313_),
    .Y(_2319_)
);

OR2X2 _23542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1924_),
    .Y(_1927_)
);

OAI21X1 _23122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1468_),
    .B(_1466_),
    .C(_1465_),
    .Y(_1469_)
);

INVX1 _14649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4071_),
    .Y(_4092_)
);

AND2X2 _14229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3339_),
    .B(_3335_),
    .Y(_3633_)
);

OAI21X1 _18482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_5921__bF$buf2),
    .C(_8294_),
    .Y(_8295_)
);

AOI21X1 _18062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7465_),
    .B(_7833_),
    .C(_7831_),
    .Y(_7834_)
);

NOR3X1 _20667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10640_),
    .B(_10636_),
    .C(_10643_),
    .Y(_10689_)
);

OAI21X1 _20247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10227_),
    .B(_10226_),
    .C(_10216_),
    .Y(_10228_)
);

OAI21X1 _11930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_2562__bF$buf0),
    .C(_2573_),
    .Y(_2584_)
);

OAI21X1 _19687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9614_),
    .B(_9615_),
    .C(_9274_),
    .Y(_9616_)
);

NAND3X1 _19267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9144_),
    .B(_9152_),
    .C(_9154_),
    .Y(_9155_)
);

AOI21X1 _12715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11132_),
    .B(_11176_),
    .C(_10430_),
    .Y(_11187_)
);

AND2X2 _22813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1131_),
    .B(_1127_),
    .Y(_1132_)
);

NOR2X1 _15187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4681_),
    .B(_4680_),
    .Y(_4682_)
);

FILL SFILL69000x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7489_),
    .B(_7494_),
    .C(_7491_),
    .Y(_7495_)
);

NOR2X1 _17333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6618_),
    .B(_7034_),
    .Y(_7035_)
);

FILL SFILL74200x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8779_),
    .B(_8374_),
    .C(_8777_),
    .Y(_8816_)
);

NOR3X1 _18538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8351_),
    .B(_8352_),
    .C(_8350_),
    .Y(_8356_)
);

INVX2 _18118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7889_),
    .Y(_7895_)
);

FILL SFILL54040x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .B(_2766_),
    .Y(_3025_)
);

OAI21X1 _13253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(_2381_),
    .C(_2385_),
    .Y(_2565_)
);

NAND2X1 _23771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2135_),
    .B(_2144_),
    .Y(_2175_)
);

NAND2X1 _23351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .B(_1717_),
    .Y(_1719_)
);

FILL SFILL64280x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4341_),
    .B(_4335_),
    .Y(_4343_)
);

OAI22X1 _14458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_10869__bF$buf2),
    .C(_7217__bF$buf2),
    .D(_9104__bF$buf2),
    .Y(_3884_)
);

NAND3X1 _14038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3423_),
    .B(_3419_),
    .C(_3386_),
    .Y(_3424_)
);

INVX2 _18291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8083_),
    .Y(_8085_)
);

AOI21X1 _20896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10936_),
    .B(_10937_),
    .C(_10934_),
    .Y(_10941_)
);

AOI21X1 _20476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10479_),
    .B(_10478_),
    .C(_10477_),
    .Y(_10480_)
);

AOI21X1 _20056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10014_),
    .B(_10018_),
    .C(_10006_),
    .Y(_10019_)
);

NOR2X1 _16604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5854_),
    .B(_6234_),
    .Y(_6235_)
);

OAI22X1 _19496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf3),
    .B(_3253__bF$buf2),
    .C(_3146__bF$buf3),
    .D(_3529__bF$buf0),
    .Y(_9406_)
);

OR2X2 _19076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8938_),
    .B(_8940_),
    .Y(_8945_)
);

AOI21X1 _17809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7541_),
    .B(_7545_),
    .C(_7527_),
    .Y(_7556_)
);

AOI21X1 _12944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1674_),
    .C(_1533_),
    .Y(_1783_)
);

NAND2X1 _12524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9071_),
    .B(_9092_),
    .Y(_9103_)
);

INVX1 _12104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .Y(_4489_)
);

NOR2X1 _22622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11875_),
    .B(_922_),
    .Y(_923_)
);

AOI21X1 _22202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_461_),
    .B(_463_),
    .C(_247_),
    .Y(_464_)
);

AOI21X1 _13729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3070_),
    .B(_3076_),
    .C(_3058_),
    .Y(_3086_)
);

OAI21X1 _13309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .B(_2447_),
    .C(_2493_),
    .Y(_2626_)
);

XNOR2X1 _23827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2215_),
    .B(_2234_),
    .Y(_2235_)
);

INVX1 _23407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1733_),
    .Y(_1779_)
);

BUFX2 BUFX2_insert410 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .Y(_2551__bF$buf3)
);

BUFX2 BUFX2_insert411 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .Y(_2551__bF$buf2)
);

BUFX2 BUFX2_insert412 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .Y(_2551__bF$buf1)
);

BUFX2 BUFX2_insert413 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .Y(_2551__bF$buf0)
);

INVX2 _17982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7709_),
    .Y(_7746_)
);

BUFX2 BUFX2_insert414 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .Y(_7225__bF$buf4)
);

BUFX2 BUFX2_insert415 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .Y(_7225__bF$buf3)
);

NAND3X1 _17562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7281_),
    .B(_7282_),
    .C(_7284_),
    .Y(_7285_)
);

AND2X2 _17142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_27_bF$buf0),
    .Y(_6825_)
);

BUFX2 BUFX2_insert416 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .Y(_7225__bF$buf2)
);

BUFX2 BUFX2_insert417 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .Y(_7225__bF$buf1)
);

BUFX2 BUFX2_insert418 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7225_),
    .Y(_7225__bF$buf0)
);

BUFX2 BUFX2_insert419 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf4)
);

XOR2X1 _18767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8541_),
    .B(_8605_),
    .Y(_8606_)
);

NAND3X1 _18347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8137_),
    .B(_8131_),
    .C(_8135_),
    .Y(_8146_)
);

NOR2X1 _13482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2596_),
    .B(_2815_),
    .Y(_2816_)
);

NOR2X1 _23580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2750_),
    .B(_2974_),
    .Y(_1967_)
);

AOI21X1 _13062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2353_),
    .B(_1412_),
    .C(_2355_),
    .Y(_2356_)
);

NOR3X1 _23160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1367_),
    .C(_1366_),
    .Y(_1510_)
);

FILL SFILL8680x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4097_),
    .B(_4126_),
    .C(_4133_),
    .Y(_4134_)
);

AOI21X1 _14267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3671_),
    .B(_3673_),
    .C(_3674_),
    .Y(_3675_)
);

FILL SFILL8600x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10267_),
    .B(_10270_),
    .C(_10208_),
    .Y(_10271_)
);

OAI21X1 _16833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6480_),
    .B(_6485_),
    .C(_6440_),
    .Y(_6486_)
);

AOI21X1 _16413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6024_),
    .B(_6025_),
    .C(_6017_),
    .Y(_6026_)
);

FILL SFILL74200x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_21_bF$buf0),
    .Y(_7346_)
);

NAND3X1 _12753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9707_),
    .B(_11527_),
    .C(_11494_),
    .Y(_11603_)
);

OAI21X1 _12333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6977_),
    .B(_6988_),
    .C(_6966_),
    .Y(_6999_)
);

NAND3X1 _22851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1172_),
    .C(_1132_),
    .Y(_1174_)
);

NOR2X1 _22431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_700_),
    .B(_697_),
    .Y(_714_)
);

OAI21X1 _22011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_11894_),
    .C(_11_),
    .Y(_254_)
);

FILL SFILL3880x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3328_),
    .B(_3327_),
    .C(_3324_),
    .Y(_3337_)
);

INVX2 _13538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .Y(_2877_)
);

OAI21X1 _13118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1663_),
    .C(_1685_),
    .Y(_2416_)
);

INVX1 _23636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .Y(_2029_)
);

XNOR2X1 _23216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1559_),
    .B(_1570_),
    .Y(_1571_)
);

FILL SFILL33800x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_31_bF$buf4),
    .C(_7116_),
    .Y(_7537_)
);

NAND3X1 _17371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7067_),
    .B(_7074_),
    .C(_7075_),
    .Y(_7077_)
);

OAI21X1 _18996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8854_),
    .B(_8857_),
    .C(_8477_),
    .Y(_8858_)
);

AND2X2 _18576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8381_),
    .B(_8379_),
    .Y(_8397_)
);

OAI22X1 _18156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_4116__bF$buf2),
    .D(_6300__bF$buf0),
    .Y(_7937_)
);

XNOR2X1 _13291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2589_),
    .B(_2581_),
    .Y(_2606_)
);

NAND3X1 _21702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11717_),
    .B(_11799_),
    .C(_11803_),
    .Y(_11824_)
);

OAI21X1 _14496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf4),
    .B(_2287__bF$buf2),
    .C(_3921_),
    .Y(_3926_)
);

NAND3X1 _14076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3458_),
    .B(_3465_),
    .C(_3248_),
    .Y(_3466_)
);

OAI21X1 _12809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_275_),
    .C(_297_),
    .Y(_308_)
);

AOI21X1 _22907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .B(_949_),
    .C(_1078_),
    .Y(_1235_)
);

NOR3X1 _20094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10045_),
    .B(_10049_),
    .C(_10050_),
    .Y(_10061_)
);

OAI21X1 _16642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_4551__bF$buf2),
    .C(_6269_),
    .Y(_6277_)
);

OAI21X1 _16222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5814_),
    .B(_5816_),
    .C(_5811_),
    .Y(_5817_)
);

FILL SFILL23720x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44200x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11379_),
    .B(_11381_),
    .C(_11380_),
    .Y(_11382_)
);

NOR3X1 _17847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7167_),
    .B(_7168_),
    .C(_7166_),
    .Y(_7598_)
);

AOI21X1 _17427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7133_),
    .B(_7132_),
    .C(_7130_),
    .Y(_7138_)
);

NAND2X1 _17007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6676_),
    .B(_6672_),
    .Y(_6677_)
);

AND2X2 _12982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1979_),
    .B(_2174_),
    .Y(_2196_)
);

NAND3X1 _12562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9411_),
    .B(_9367_),
    .C(_9433_),
    .Y(_9510_)
);

OAI21X1 _12142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3372_),
    .B(_3986_),
    .C(_4895_),
    .Y(_4906_)
);

NAND2X1 _22660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_27_bF$buf1),
    .Y(_964_)
);

OAI21X1 _22240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_256_),
    .C(_281_),
    .Y(_504_)
);

FILL SFILL8680x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3126_),
    .Y(_3127_)
);

NOR2X1 _23865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2274_),
    .B(_2265_),
    .Y(_2275_)
);

INVX1 _13347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2667_),
    .Y(_2668_)
);

XOR2X1 _23445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1818_),
    .B(_1806_),
    .Y(_1821_)
);

AND2X2 _23025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1360_),
    .Y(_1363_)
);

FILL SFILL8600x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6859_),
    .B(_6862_),
    .C(_6865_),
    .Y(_6866_)
);

NAND2X1 _15913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_16_bF$buf4),
    .Y(_5478_)
);

NAND2X1 _18385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7862_),
    .B(_7868_),
    .Y(_8188_)
);

NOR2X1 _21931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11817_),
    .B(_11810_),
    .Y(_167_)
);

AND2X2 _21511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_27_bF$buf4),
    .Y(_11615_)
);

NOR2X1 _12618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8588_),
    .B(_10112_),
    .Y(_10123_)
);

OAI21X1 _22716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1025_),
    .C(_879_),
    .Y(_1026_)
);

FILL SFILL64200x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _16871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf0),
    .B(_3253__bF$buf3),
    .C(_9104__bF$buf3),
    .D(_3529__bF$buf1),
    .Y(_6528_)
);

NAND3X1 _16451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6061_),
    .B(_6065_),
    .C(_6064_),
    .Y(_6066_)
);

NOR3X1 _16031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5231_),
    .B(_5232_),
    .C(_5230_),
    .Y(_5608_)
);

FILL SFILL28840x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7383_),
    .B(_7387_),
    .C(_7386_),
    .Y(_7388_)
);

NOR2X1 _17236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6863_),
    .B(_6927_),
    .Y(_6928_)
);

OAI21X1 _12791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_45_),
    .B(_56_),
    .C(_23_),
    .Y(_111_)
);

OAI21X1 _12371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf3),
    .B(_5420__bF$buf2),
    .C(_7360_),
    .Y(_7415_)
);

OAI21X1 _13996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3375_),
    .B(_3376_),
    .C(_3377_),
    .Y(_3378_)
);

NAND3X1 _13576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2918_),
    .B(_2909_),
    .C(_2841_),
    .Y(_2919_)
);

NAND2X1 _13156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf2),
    .B(areg_13_bF$buf1),
    .Y(_2459_)
);

OAI21X1 _23674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2015_),
    .B(_2011_),
    .C(_2069_),
    .Y(_2070_)
);

AOI21X1 _23254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_1436_),
    .C(_1480_),
    .Y(_1613_)
);

OAI21X1 _19802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9476_),
    .B(_9478_),
    .C(_9474_),
    .Y(_9742_)
);

DFFPOSX1 _24039_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[29]),
    .CLK(clk_bF$buf1),
    .D(a[29])
);

OAI21X1 _15722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5266_),
    .B(_5268_),
    .C(_5265_),
    .Y(_5269_)
);

OAI21X1 _15302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4802_),
    .B(_4803_),
    .C(_4804_),
    .Y(_4809_)
);

OAI21X1 _18194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7978_),
    .C(_7957_),
    .Y(_7979_)
);

FILL SFILL8760x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44200x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10828_),
    .B(_10833_),
    .C(_10821_),
    .Y(_10834_)
);

AOI21X1 _20379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10371_),
    .B(_10372_),
    .C(_10357_),
    .Y(_10373_)
);

AOI21X1 _16927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6583_),
    .B(_6587_),
    .C(_6588_),
    .Y(_6589_)
);

AOI21X1 _16507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5975_),
    .B(_5981_),
    .C(_5838_),
    .Y(_6128_)
);

NAND2X1 _21740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11864_),
    .B(_11859_),
    .Y(_11865_)
);

NAND3X1 _21320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11370_),
    .B(_11400_),
    .C(_11404_),
    .Y(_11405_)
);

NOR3X1 _19399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9285_),
    .B(_9294_),
    .C(_9295_),
    .Y(_9299_)
);

FILL SFILL48920x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_680_),
    .B(_713_),
    .C(_396_),
    .Y(_724_)
);

OAI21X1 _12427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7898_),
    .B(_7909_),
    .C(_7558_),
    .Y(_8040_)
);

OAI21X1 _22945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf2),
    .B(_5668__bF$buf1),
    .C(_1113_),
    .Y(_1276_)
);

OAI21X1 _12007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .B(_2727_),
    .C(_3416_),
    .Y(_3427_)
);

NOR3X1 _22525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_576_),
    .C(_577_),
    .Y(_817_)
);

AOI21X1 _22105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_347_),
    .C(_293_),
    .Y(_357_)
);

NAND2X1 _16680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_28_bF$buf4),
    .Y(_6318_)
);

NAND3X1 _16260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5846_),
    .B(_5853_),
    .C(_5857_),
    .Y(_5858_)
);

OAI21X1 _17885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5660_),
    .B(_6033_),
    .C(_6029_),
    .Y(_7639_)
);

AOI21X1 _17465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6600_),
    .B(_6755_),
    .C(_7178_),
    .Y(_7179_)
);

NAND3X1 _17045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6707_),
    .B(_6709_),
    .C(_6702_),
    .Y(_6719_)
);

AOI21X1 _12180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5233_),
    .B(_5168_),
    .C(_5124_),
    .Y(_5321_)
);

FILL SFILL38920x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2709_),
    .B(_2708_),
    .C(_2707_),
    .Y(_2710_)
);

NAND3X1 _23483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .B(_1859_),
    .C(_1775_),
    .Y(_1863_)
);

AOI21X1 _23063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .B(_1389_),
    .C(_1403_),
    .Y(_1404_)
);

FILL SFILL28920x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_28_bF$buf1),
    .Y(_9533_)
);

NAND2X1 _15951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5517_),
    .B(_5518_),
    .Y(_5520_)
);

NAND3X1 _15531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5051_),
    .B(_5054_),
    .C(_5057_),
    .Y(_5059_)
);

NAND3X1 _15111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4440_),
    .B(_4433_),
    .C(_4438_),
    .Y(_4600_)
);

FILL SFILL28840x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf0),
    .B(_6300__bF$buf1),
    .C(_9811_),
    .Y(_10164_)
);

AOI21X1 _16736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5835_),
    .B(_5987_),
    .C(_6379_),
    .Y(_6380_)
);

OR2X2 _16316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5918_),
    .B(_5919_),
    .Y(_5920_)
);

NAND2X1 _12656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10507_),
    .B(_10529_),
    .Y(_10540_)
);

OAI21X1 _12236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5914_),
    .B(_5925_),
    .C(_5870_),
    .Y(_5936_)
);

NOR3X1 _22754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(_1062_),
    .C(_1067_),
    .Y(_1068_)
);

OAI21X1 _22334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_428_),
    .B(_430_),
    .C(_426_),
    .Y(_608_)
);

DFFPOSX1 _23959_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[13]),
    .CLK(clk_bF$buf2),
    .D(_0_[13])
);

NAND3X1 _23539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1921_),
    .B(_1920_),
    .C(_1922_),
    .Y(_1923_)
);

INVX2 _23119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .Y(_1465_)
);

INVX2 _14802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4236_),
    .Y(_4261_)
);

NAND2X1 _17694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6990_),
    .B(_6997_),
    .Y(_7430_)
);

NAND2X1 _17274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf2),
    .B(breg_15_bF$buf2),
    .Y(_6970_)
);

NAND2X1 _20820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10855_),
    .B(_10856_),
    .Y(_10857_)
);

NAND2X1 _20400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_25_bF$buf0),
    .Y(_10396_)
);

OAI21X1 _18899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf2),
    .B(_7100__bF$buf2),
    .C(_8747_),
    .Y(_8751_)
);

AND2X2 _18479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_24_bF$buf1),
    .Y(_8291_)
);

NAND3X1 _18059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7820_),
    .B(_7828_),
    .C(_7829_),
    .Y(_7830_)
);

NAND3X1 _13194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2422_),
    .B(_2495_),
    .C(_2500_),
    .Y(_2501_)
);

NAND3X1 _23292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(_1548_),
    .C(_1650_),
    .Y(_1654_)
);

NAND3X1 _19840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9778_),
    .B(_9782_),
    .C(_9764_),
    .Y(_9783_)
);

NAND2X1 _19420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_26_bF$buf3),
    .Y(_9322_)
);

NAND3X1 _19000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8480_),
    .B(_8853_),
    .C(_8846_),
    .Y(_8862_)
);

INVX8 _11927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .Y(_2551_)
);

NAND2X1 _21605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11509_),
    .B(_11514_),
    .Y(_11717_)
);

OAI21X1 _14399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf0),
    .B(_2763_),
    .C(_3818_),
    .Y(_3819_)
);

NAND2X1 _15760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_26_bF$buf4),
    .Y(_5309_)
);

AOI22X1 _15340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_21_bF$buf1),
    .C(breg_4_bF$buf3),
    .D(areg_20_bF$buf3),
    .Y(_4850_)
);

INVX2 _16965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6605_),
    .Y(_6631_)
);

NAND2X1 _16545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6168_),
    .B(_6169_),
    .Y(_6170_)
);

AOI21X1 _16125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5397_),
    .B(_5378_),
    .C(_5401_),
    .Y(_5710_)
);

FILL SFILL59080x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69320x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1118_),
    .B(_1129_),
    .C(_1107_),
    .Y(_1140_)
);

NAND3X1 _12465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8249_),
    .B(_8183_),
    .C(_8227_),
    .Y(_8446_)
);

XNOR2X1 _22983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1310_),
    .B(_1299_),
    .Y(_1317_)
);

NAND3X1 _12045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3788_),
    .B(_3799_),
    .C(_3832_),
    .Y(_3843_)
);

NAND2X1 _22563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_857_),
    .Y(_859_)
);

NOR2X1 _22143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_392_),
    .Y(_399_)
);

FILL SFILL28920x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520__bF$buf2),
    .B(_7225__bF$buf1),
    .Y(_2171_)
);

NOR2X1 _23348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1713_),
    .B(_1714_),
    .Y(_1715_)
);

XNOR2X1 _14611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3773_),
    .B(_4050_),
    .Y(_0_[21])
);

OAI21X1 _17083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6753_),
    .B(_6754_),
    .C(_6602_),
    .Y(_6761_)
);

FILL SFILL18920x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _15816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5370_),
    .Y(_5371_)
);

INVX1 _18288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8080_),
    .Y(_8081_)
);

NOR3X1 _21834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11741_),
    .B(_11739_),
    .C(_11735_),
    .Y(_60_)
);

NAND3X1 _21414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11503_),
    .B(_11504_),
    .C(_11473_),
    .Y(_11509_)
);

NAND2X1 _22619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_919_),
    .Y(_0_[47])
);

NAND2X1 _16774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6124_),
    .B(_6386_),
    .Y(_6421_)
);

NAND3X1 _16354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_5910_),
    .C(_5909_),
    .Y(_5962_)
);

BUFX2 BUFX2_insert380 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .Y(_2519__bF$buf3)
);

BUFX2 BUFX2_insert381 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .Y(_2519__bF$buf2)
);

BUFX2 BUFX2_insert382 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .Y(_2519__bF$buf1)
);

BUFX2 BUFX2_insert383 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .Y(_2519__bF$buf0)
);

BUFX2 BUFX2_insert384 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf4)
);

AOI21X1 _17979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7376_),
    .B(_7374_),
    .C(_7741_),
    .Y(_7742_)
);

INVX1 _17559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7276_),
    .Y(_7281_)
);

BUFX2 BUFX2_insert385 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf3)
);

BUFX2 BUFX2_insert386 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf2)
);

NAND2X1 _17139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_27_bF$buf0),
    .Y(_6821_)
);

BUFX2 BUFX2_insert387 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf1)
);

BUFX2 BUFX2_insert388 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[8]),
    .Y(areg_8_bF$buf0)
);

AOI21X1 _12694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9060_),
    .B(_9115_),
    .C(_9148_),
    .Y(_10957_)
);

BUFX2 BUFX2_insert389 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[25]),
    .Y(areg_25_bF$buf4)
);

OAI21X1 _12274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5321_),
    .B(_5299_),
    .C(_5244_),
    .Y(_6352_)
);

NAND2X1 _22792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_957_),
    .B(_969_),
    .Y(_1109_)
);

XOR2X1 _22372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_642_),
    .Y(_650_)
);

OAI21X1 _18920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_8773_),
    .C(_8369_),
    .Y(_8774_)
);

AOI21X1 _18500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8312_),
    .B(_8313_),
    .C(_8311_),
    .Y(_8314_)
);

INVX1 _13899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3271_),
    .Y(_3272_)
);

INVX1 _13479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2806_),
    .Y(_2812_)
);

DFFPOSX1 _23997_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[51]),
    .CLK(clk_bF$buf6),
    .D(_0_[51])
);

XOR2X1 _13059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1412_),
    .B(_2353_),
    .Y(_0_[14])
);

AND2X2 _23577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4639_),
    .B(_4636_),
    .Y(_1964_)
);

INVX1 _23157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1503_),
    .Y(_1507_)
);

FILL SFILL3720x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9613_),
    .B(_9616_),
    .C(_9272_),
    .Y(_9635_)
);

NAND3X1 _14840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4147_),
    .B(_4141_),
    .C(_4145_),
    .Y(_4302_)
);

NAND3X1 _14420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3816_),
    .B(_3823_),
    .C(_3819_),
    .Y(_3842_)
);

AOI21X1 _14000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3368_),
    .B(_3371_),
    .C(_3373_),
    .Y(_3382_)
);

FILL SFILL3640x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48760x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3402__bF$buf2),
    .C(_5155_),
    .Y(_5162_)
);

OAI21X1 _15205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4700_),
    .B(_4701_),
    .C(_4684_),
    .Y(_4702_)
);

FILL SFILL59080x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7783_),
    .B(_7867_),
    .C(_7871_),
    .Y(_7872_)
);

NAND2X1 _11965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2957_),
    .B(_2880_),
    .Y(_2968_)
);

AND2X2 _21643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_11759_)
);

AOI21X1 _21223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11298_),
    .B(_11299_),
    .C(_11006_),
    .Y(_11300_)
);

AOI21X1 _22848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1169_),
    .C(_1161_),
    .Y(_1170_)
);

NAND2X1 _22428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_707_),
    .Y(_711_)
);

NAND2X1 _22008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_75_),
    .Y(_250_)
);

FILL SFILL49080x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6211_),
    .B(_6206_),
    .C(_6130_),
    .Y(_6212_)
);

XNOR2X1 _16163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5751_),
    .B(_5748_),
    .Y(_5752_)
);

AOI22X1 _17788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_31_bF$buf1),
    .C(breg_1_bF$buf5),
    .D(areg_30_bF$buf5),
    .Y(_7533_)
);

FILL SFILL18840x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7068_),
    .B(_7072_),
    .C(_7071_),
    .Y(_7073_)
);

NOR2X1 _12083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf2),
    .B(_4258__bF$buf3),
    .Y(_4259_)
);

AOI21X1 _22181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_436_),
    .C(_435_),
    .Y(_441_)
);

FILL SFILL23880x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL63960x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _20914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10605_),
    .B(_10950_),
    .Y(_10961_)
);

XNOR2X1 _13288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .B(_2601_),
    .Y(_2602_)
);

NAND3X1 _23386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1755_),
    .B(_1756_),
    .C(_1754_),
    .Y(_1757_)
);

OAI21X1 _19934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9880_),
    .B(_9881_),
    .C(_9862_),
    .Y(_9887_)
);

AND2X2 _19514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_20_bF$buf0),
    .Y(_9426_)
);

NAND2X1 _15854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5411_),
    .B(_5412_),
    .Y(_5413_)
);

AOI21X1 _15434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4953_),
    .B(_4952_),
    .C(_4652_),
    .Y(_4954_)
);

NAND3X1 _15014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4475_),
    .B(_4482_),
    .C(_4483_),
    .Y(_4493_)
);

FILL SFILL29000x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6268_),
    .B(_6272_),
    .C(_6271_),
    .Y(_6273_)
);

OAI21X1 _16219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5799_),
    .B(_5800_),
    .C(_5797_),
    .Y(_5813_)
);

XNOR2X1 _21872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_96_),
    .Y(_102_)
);

AOI21X1 _21452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11545_),
    .B(_11550_),
    .C(_11438_),
    .Y(_11551_)
);

OAI21X1 _21032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10820_),
    .B(_11089_),
    .C(_10845_),
    .Y(_11090_)
);

INVX2 _12979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2153_),
    .Y(_2163_)
);

NAND3X1 _12559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8698_),
    .B(_9422_),
    .C(_9466_),
    .Y(_9477_)
);

OAI21X1 _12139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4807_),
    .B(_4818_),
    .C(_3460_),
    .Y(_4873_)
);

OAI21X1 _22657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_747_),
    .B(_959_),
    .C(_960_),
    .Y(_961_)
);

FILL SFILL3720x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _22237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_340_),
    .Y(_501_)
);

FILL SFILL74360x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3078_),
    .B(_3082_),
    .C(_3083_),
    .Y(_3295_)
);

OAI21X1 _13500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .B(_2602_),
    .C(_2604_),
    .Y(_2835_)
);

NAND3X1 _16392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5996_),
    .B(_5743_),
    .C(_6002_),
    .Y(_6003_)
);

OAI21X1 _14705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3913_),
    .B(_4153_),
    .C(_4009_),
    .Y(_4154_)
);

OAI21X1 _17597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7318_),
    .B(_7319_),
    .C(_7273_),
    .Y(_7323_)
);

NAND2X1 _17177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_22_bF$buf1),
    .Y(_6863_)
);

INVX1 _20723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10744_),
    .Y(_10751_)
);

NAND3X1 _20303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10283_),
    .B(_10290_),
    .C(_10108_),
    .Y(_10291_)
);

OAI21X1 _13097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf2),
    .B(_6044__bF$buf2),
    .C(_1598_),
    .Y(_2394_)
);

OAI21X1 _23195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1527_),
    .C(_1525_),
    .Y(_1548_)
);

AOI21X1 _19743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9676_),
    .B(_9672_),
    .C(_9648_),
    .Y(_9677_)
);

NAND3X1 _19323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9204_),
    .B(_9197_),
    .C(_9095_),
    .Y(_9217_)
);

FILL SFILL33880x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_150_),
    .C(_156_),
    .Y(_163_)
);

NAND2X1 _21508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_29_bF$buf4),
    .Y(_11611_)
);

NOR2X1 _15663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4863_),
    .B(_5203_),
    .Y(_5204_)
);

AOI21X1 _15243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4742_),
    .B(_4743_),
    .C(_4735_),
    .Y(_4744_)
);

OAI21X1 _16868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf3),
    .B(_3529__bF$buf1),
    .C(_6523_),
    .Y(_6524_)
);

AND2X2 _16448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_24_bF$buf5),
    .Y(_6063_)
);

NAND3X1 _16028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5584_),
    .B(_5591_),
    .C(_5594_),
    .Y(_5604_)
);

AOI21X1 _21681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11796_),
    .B(_11797_),
    .C(_11795_),
    .Y(_11801_)
);

FILL SFILL23880x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11335_),
    .B(_11339_),
    .C(_11338_),
    .Y(_11340_)
);

FILL SFILL54280x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_45_),
    .B(_56_),
    .C(_67_),
    .Y(_78_)
);

NAND2X1 _12368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf5),
    .B(areg_6_bF$buf4),
    .Y(_7382_)
);

XOR2X1 _22886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1211_),
    .B(_1202_),
    .Y(_1212_)
);

FILL SFILL23800x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_748_),
    .Y(_752_)
);

NAND3X1 _22046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .B(_291_),
    .C(_290_),
    .Y(_292_)
);

FILL SFILL8760x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4158_),
    .B(_4159_),
    .Y(_4405_)
);

NAND2X1 _14514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3940_),
    .B(_3945_),
    .Y(_3946_)
);

FILL SFILL29000x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5006_),
    .B(_5002_),
    .Y(_5265_)
);

NOR2X1 _20952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10994_),
    .B(_11001_),
    .Y(_11002_)
);

OAI21X1 _20532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10541_),
    .B(_10209_),
    .C(_10252_),
    .Y(_10542_)
);

AOI21X1 _20112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10065_),
    .B(_10070_),
    .C(_10071_),
    .Y(_10081_)
);

NOR2X1 _19972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9922_),
    .B(_9917_),
    .Y(_9928_)
);

AOI21X1 _19552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9465_),
    .B(_9467_),
    .C(_9464_),
    .Y(_9468_)
);

NOR2X1 _19132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf1),
    .B(_5369_),
    .Y(_9007_)
);

NAND3X1 _21737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11597_),
    .B(_11856_),
    .C(_11857_),
    .Y(_11862_)
);

AOI21X1 _21317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11387_),
    .B(_11392_),
    .C(_11371_),
    .Y(_11402_)
);

FILL SFILL43960x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5452_),
    .B(_5451_),
    .C(_5454_),
    .Y(_5455_)
);

NAND3X1 _15472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4662_),
    .B(_4988_),
    .C(_4989_),
    .Y(_4994_)
);

XOR2X1 _15052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4534_),
    .B(_4529_),
    .Y(_4535_)
);

INVX2 _16677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6314_),
    .Y(_6315_)
);

NOR2X1 _16257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5481_),
    .B(_5854_),
    .Y(_5855_)
);

NAND3X1 _21490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11317_),
    .B(_11587_),
    .C(_11588_),
    .Y(_11591_)
);

NOR2X1 _21070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10950_),
    .B(_10605_),
    .Y(_11131_)
);

FILL SFILL64360x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8413_),
    .B(_9883_),
    .Y(_0_[11])
);

NAND3X1 _12177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5091_),
    .B(_5244_),
    .C(_5278_),
    .Y(_5289_)
);

NAND2X1 _22695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_999_),
    .Y(_1003_)
);

NAND2X1 _22275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_320_),
    .Y(_543_)
);

AOI21X1 _18823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8250_),
    .B(_8252_),
    .C(_8257_),
    .Y(_8668_)
);

OAI21X1 _18403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8202_),
    .B(_8207_),
    .C(_8196_),
    .Y(_8208_)
);

AOI21X1 _19608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .B(_9146_),
    .C(_9161_),
    .Y(_9529_)
);

AND2X2 _14743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3903_),
    .B(_3897_),
    .Y(_4196_)
);

NAND3X1 _14323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3586_),
    .B(_3578_),
    .C(_3583_),
    .Y(_3737_)
);

DFFPOSX1 _24001_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[55]),
    .CLK(clk_bF$buf9),
    .D(_0_[55])
);

NOR2X1 _15948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_3146__bF$buf3),
    .Y(_5516_)
);

NAND2X1 _15528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_13_bF$buf3),
    .Y(_5055_)
);

AOI21X1 _15108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4578_),
    .B(_4583_),
    .C(_4495_),
    .Y(_4596_)
);

OAI21X1 _20761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10790_),
    .B(_10791_),
    .C(_10787_),
    .Y(_10793_)
);

NAND3X1 _20341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10317_),
    .B(_10322_),
    .C(_9992_),
    .Y(_10333_)
);

AOI21X1 _19781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9713_),
    .B(_9714_),
    .C(_9712_),
    .Y(_9719_)
);

NAND2X1 _19361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9252_),
    .B(_9253_),
    .Y(_9258_)
);

AOI21X1 _21966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_204_),
    .C(_11826_),
    .Y(_205_)
);

NAND2X1 _21546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf1),
    .B(breg_24_bF$buf0),
    .Y(_11652_)
);

INVX2 _21126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11169_),
    .Y(_11193_)
);

FILL SFILL74200x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4778_),
    .B(_4779_),
    .Y(_4786_)
);

FILL SFILL13880x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6081_),
    .B(_6085_),
    .C(_6094_),
    .Y(_6105_)
);

NAND3X1 _16066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5642_),
    .B(_5303_),
    .C(_5645_),
    .Y(_5646_)
);

FILL SFILL74120x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .C(_333_),
    .Y(_334_)
);

AOI21X1 _18632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7655_),
    .B(_8056_),
    .C(_8062_),
    .Y(_8459_)
);

OAI21X1 _18212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7924_),
    .B(_7923_),
    .C(_7881_),
    .Y(_7999_)
);

INVX1 _20817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10853_),
    .Y(_10854_)
);

NAND3X1 _23289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1647_),
    .B(_1650_),
    .C(_1646_),
    .Y(_1651_)
);

NOR3X1 _19837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9766_),
    .B(_9775_),
    .C(_9776_),
    .Y(_9780_)
);

OAI21X1 _19417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9318_),
    .B(_8975_),
    .C(_8967_),
    .Y(_9319_)
);

OAI21X1 _14972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4290_),
    .B(_4446_),
    .C(_4280_),
    .Y(_4447_)
);

NAND3X1 _14552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3969_),
    .B(_3977_),
    .C(_3955_),
    .Y(_3988_)
);

NOR2X1 _14132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_3526_),
    .Y(_3527_)
);

INVX2 _15757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5305_),
    .Y(_5306_)
);

OAI21X1 _15337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4846_),
    .B(_4559_),
    .C(_4549_),
    .Y(_4847_)
);

OAI21X1 _20990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11038_),
    .B(_11039_),
    .C(_11035_),
    .Y(_11042_)
);

NAND3X1 _20570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10575_),
    .B(_10572_),
    .C(_10569_),
    .Y(_10583_)
);

AND2X2 _20150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf5),
    .B(areg_20_bF$buf1),
    .Y(_10122_)
);

NAND3X1 _19590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9502_),
    .B(_9508_),
    .C(_9487_),
    .Y(_9509_)
);

NAND3X1 _19170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9044_),
    .B(_9047_),
    .C(_9046_),
    .Y(_9048_)
);

OAI21X1 _21775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_11902_),
    .Y(_11903_)
);

OAI21X1 _21355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11383_),
    .B(_11442_),
    .C(_11443_),
    .Y(_11444_)
);

OAI21X1 _17903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7658_),
    .B(_7618_),
    .C(_7611_),
    .Y(_7659_)
);

NAND3X1 _15090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4575_),
    .B(_4573_),
    .C(_4574_),
    .Y(_4576_)
);

AOI21X1 _13823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3182_),
    .B(_3189_),
    .C(_3095_),
    .Y(_3190_)
);

BUFX2 _23921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[39]),
    .Y(y[39])
);

OAI21X1 _13403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .B(_2726_),
    .C(_2556_),
    .Y(_2730_)
);

NOR2X1 _23501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1679_),
    .B(_1880_),
    .Y(_1882_)
);

OAI21X1 _16295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf0),
    .B(_3958__bF$buf1),
    .C(_5893_),
    .Y(_5897_)
);

AOI22X1 _14608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3774_),
    .B(_3519_),
    .C(_4043_),
    .D(_4042_),
    .Y(_4048_)
);

FILL SFILL44040x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8703_),
    .Y(_8710_)
);

OAI21X1 _18441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7825_),
    .B(_8248_),
    .C(_7827_),
    .Y(_8250_)
);

AND2X2 _18021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7721_),
    .B(_7786_),
    .Y(_7789_)
);

NOR3X1 _20626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10622_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10645_)
);

AOI21X1 _20206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10132_),
    .B(_10133_),
    .C(_10117_),
    .Y(_10184_)
);

OAI21X1 _23098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315__bF$buf0),
    .B(_7100__bF$buf1),
    .C(_1301_),
    .Y(_1442_)
);

OAI21X1 _19646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9570_),
    .B(_9569_),
    .C(_9482_),
    .Y(_9571_)
);

AND2X2 _19226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_26_bF$buf3),
    .Y(_9110_)
);

AND2X2 _14781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_19_bF$buf0),
    .Y(_4238_)
);

NAND2X1 _14361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3578_),
    .B(_3584_),
    .Y(_3777_)
);

FILL SFILL43880x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf1),
    .B(areg_26_bF$buf2),
    .Y(_5558_)
);

AND2X2 _15566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4747_),
    .B(_4739_),
    .Y(_5097_)
);

NAND3X1 _15146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4625_),
    .B(_4628_),
    .C(_4631_),
    .Y(_4638_)
);

AOI21X1 _21584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11678_),
    .B(_11684_),
    .C(_11648_),
    .Y(_11694_)
);

INVX2 _21164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11234_),
    .Y(_11235_)
);

OAI22X1 _17712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_4551__bF$buf1),
    .C(_7217__bF$buf1),
    .D(_3961__bF$buf2),
    .Y(_7450_)
);

FILL SFILL59160x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf2),
    .B(_7225__bF$buf0),
    .Y(_1105_)
);

OAI21X1 _22369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_8773_),
    .C(_405_),
    .Y(_646_)
);

NAND2X1 _18917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_29_bF$buf0),
    .Y(_8771_)
);

OAI21X1 _13632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .B(_2979_),
    .C(_2977_),
    .Y(_2980_)
);

AOI21X1 _13212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2506_),
    .B(_2512_),
    .C(_2374_),
    .Y(_2521_)
);

NOR2X1 _23730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100__bF$buf3),
    .B(_7225__bF$buf1),
    .Y(_2130_)
);

INVX1 _23310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .Y(_1673_)
);

AOI21X1 _14837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4280_),
    .B(_4286_),
    .C(_4200_),
    .Y(_4299_)
);

NAND2X1 _14417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3549_),
    .B(_3545_),
    .Y(_3839_)
);

FILL SFILL28680x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74040x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8094_),
    .B(_8498_),
    .Y(_8499_)
);

AOI21X1 _18250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8033_),
    .B(_8038_),
    .C(_7661_),
    .Y(_8039_)
);

FILL SFILL54120x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10895_),
    .B(_10591_),
    .C(_10586_),
    .Y(_10896_)
);

NAND3X1 _20435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10429_),
    .B(_10392_),
    .C(_10434_),
    .Y(_10435_)
);

OAI21X1 _20015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9971_),
    .B(_9974_),
    .C(_9636_),
    .Y(_9975_)
);

FILL SFILL54040x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9815_),
    .B(_9821_),
    .C(_9791_),
    .Y(_9822_)
);

NAND2X1 _19455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8959_),
    .B(_8964_),
    .Y(_9361_)
);

INVX2 _19035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8899_),
    .Y(_8900_)
);

AOI21X1 _14590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4027_),
    .B(_4028_),
    .C(_4026_),
    .Y(_4029_)
);

AOI21X1 _14170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3563_),
    .B(_3564_),
    .C(_3562_),
    .Y(_3568_)
);

FILL SFILL59240x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1195_),
    .B(_1151_),
    .Y(_1336_)
);

OAI21X1 _15795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5344_),
    .B(_5347_),
    .C(_5308_),
    .Y(_5348_)
);

OAI21X1 _15375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4882_),
    .B(_4881_),
    .C(_4847_),
    .Y(_4889_)
);

FILL SFILL48760x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11476_),
    .B(_11484_),
    .C(_11485_),
    .Y(_11486_)
);

NOR3X1 _17941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7697_),
    .B(_7698_),
    .C(_7699_),
    .Y(_7701_)
);

NAND2X1 _17521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7237_),
    .B(_7238_),
    .Y(_7240_)
);

AOI21X1 _17101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6383_),
    .B(_6127_),
    .C(_6779_),
    .Y(_6781_)
);

AOI21X1 _22598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_896_),
    .C(_729_),
    .Y(_897_)
);

NAND3X1 _22178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(_428_),
    .C(_422_),
    .Y(_437_)
);

AOI21X1 _18726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8554_),
    .B(_8556_),
    .C(_8553_),
    .Y(_8561_)
);

OAI21X1 _18306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf4),
    .B(_6050__bF$buf0),
    .C(_8090_),
    .Y(_8101_)
);

OAI21X1 _13861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3218_),
    .B(_3222_),
    .C(_3225_),
    .Y(_3232_)
);

FILL SFILL69240x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2561_),
    .B(_2768_),
    .C(_2769_),
    .Y(_2771_)
);

NAND3X1 _13021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2315_),
    .C(_2313_),
    .Y(_2316_)
);

FILL SFILL69160x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4075_),
    .B(_4077_),
    .C(_4080_),
    .Y(_4089_)
);

OAI21X1 _14226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3380_),
    .B(_3382_),
    .C(_3374_),
    .Y(_3630_)
);

FILL SFILL69080x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9264_),
    .B(_10685_),
    .Y(_10686_)
);

NAND2X1 _20244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_29_bF$buf3),
    .Y(_10225_)
);

NAND3X1 _19684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9273_),
    .B(_9606_),
    .C(_9607_),
    .Y(_9613_)
);

OAI21X1 _19264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf1),
    .B(_7520__bF$buf0),
    .C(_9146_),
    .Y(_9152_)
);

FILL SFILL28760x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_97_),
    .Y(_98_)
);

NAND3X1 _21449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11522_),
    .B(_11539_),
    .C(_11518_),
    .Y(_11547_)
);

OAI21X1 _21029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11078_),
    .B(_11076_),
    .C(_11074_),
    .Y(_11086_)
);

OAI21X1 _12712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11099_),
    .B(_11110_),
    .C(_11066_),
    .Y(_11154_)
);

NAND2X1 _22810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1110_),
    .Y(_1128_)
);

NAND2X1 _15184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_22_bF$buf2),
    .Y(_4679_)
);

FILL FILL74120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3288_),
    .B(_3289_),
    .C(_3259_),
    .Y(_3292_)
);

AOI21X1 _16389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .B(_5994_),
    .C(_5992_),
    .Y(_5999_)
);

FILL FILL74040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7486_),
    .B(_7490_),
    .Y(_7491_)
);

OAI21X1 _17330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_3961__bF$buf2),
    .C(_6618_),
    .Y(_7030_)
);

FILL SFILL39080x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _18955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8809_),
    .B(_8810_),
    .C(_8812_),
    .D(_8811_),
    .Y(_8813_)
);

OAI21X1 _18535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8350_),
    .B(_8351_),
    .C(_8352_),
    .Y(_8353_)
);

AND2X2 _18115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_22_bF$buf4),
    .Y(_7892_)
);

AOI21X1 _13670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3016_),
    .B(_3017_),
    .C(_3015_),
    .Y(_3021_)
);

NAND2X1 _13250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg_15_bF$buf1),
    .Y(_2561_)
);

OAI21X1 _14875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4339_),
    .B(_4340_),
    .C(_4338_),
    .Y(_4341_)
);

AOI21X1 _14455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3878_),
    .B(_3880_),
    .C(_3875_),
    .Y(_3881_)
);

OAI21X1 _14035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3415_),
    .B(_3417_),
    .C(_3396_),
    .Y(_3421_)
);

NAND3X1 _20893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10936_),
    .B(_10937_),
    .C(_10934_),
    .Y(_10938_)
);

INVX2 _20473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10470_),
    .Y(_10477_)
);

NOR2X1 _20053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9660_),
    .B(_10015_),
    .Y(_10016_)
);

OAI21X1 _16601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_3402__bF$buf0),
    .C(_5854_),
    .Y(_6232_)
);

AND2X2 _19493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_9403_)
);

AND2X2 _19073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8938_),
    .B(_8940_),
    .Y(_8942_)
);

NAND3X1 _21678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11780_),
    .B(_11784_),
    .C(_11787_),
    .Y(_11797_)
);

AND2X2 _21258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_27_bF$buf5),
    .Y(_11337_)
);

NOR3X1 _17806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7121_),
    .B(_7126_),
    .C(_7127_),
    .Y(_7553_)
);

FILL SFILL69240x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1740_),
    .B(_341_),
    .C(_242_),
    .Y(_1751_)
);

INVX2 _12521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9049_),
    .Y(_9060_)
);

OAI21X1 _12101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4336_),
    .B(_4423_),
    .C(_4445_),
    .Y(_4466_)
);

OAI21X1 _13726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2864_),
    .B(_2866_),
    .C(_2856_),
    .Y(_3083_)
);

AOI21X1 _13306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2604_),
    .B(_2609_),
    .C(_2611_),
    .Y(_2623_)
);

OAI21X1 _23824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2191_),
    .B(_2189_),
    .C(_2187_),
    .Y(_2232_)
);

INVX1 _23404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1775_),
    .Y(_1776_)
);

NAND3X1 _16198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5784_),
    .B(_5788_),
    .C(_5787_),
    .Y(_5789_)
);

FILL SFILL3800x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_8603_)
);

OAI21X1 _18344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8142_),
    .B(_8141_),
    .C(_8137_),
    .Y(_8143_)
);

INVX1 _20949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10998_),
    .Y(_10999_)
);

NAND3X1 _20529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10528_),
    .B(_10522_),
    .C(_10526_),
    .Y(_10538_)
);

NAND3X1 _20109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10043_),
    .B(_10076_),
    .C(_10072_),
    .Y(_10077_)
);

AND2X2 _19969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9527_),
    .B(_9523_),
    .Y(_9924_)
);

AND2X2 _19549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9423_),
    .B(_9418_),
    .Y(_9464_)
);

AOI21X1 _19129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8805_),
    .B(_8823_),
    .C(_8694_),
    .Y(_9003_)
);

AOI21X1 _14684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4130_),
    .B(_4129_),
    .C(_4122_),
    .Y(_4131_)
);

NAND2X1 _14264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf4),
    .B(areg_17_bF$buf1),
    .Y(_3672_)
);

FILL FILL74120x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .B(_5447_),
    .C(_5445_),
    .Y(_5451_)
);

AOI21X1 _15469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4988_),
    .B(_4989_),
    .C(_4662_),
    .Y(_4990_)
);

AND2X2 _15049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_20_bF$buf3),
    .Y(_4531_)
);

NAND3X1 _20282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10251_),
    .B(_10252_),
    .C(_10253_),
    .Y(_10268_)
);

FILL SFILL18760x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6466_),
    .B(_6470_),
    .C(_6478_),
    .Y(_6482_)
);

AOI21X1 _16410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5306_),
    .B(_5641_),
    .C(_5643_),
    .Y(_6022_)
);

NAND3X1 _21487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11587_),
    .B(_11588_),
    .C(_11586_),
    .Y(_11589_)
);

OAI21X1 _21067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11120_),
    .B(_11119_),
    .C(_11117_),
    .Y(_11128_)
);

OAI21X1 _17615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7173_),
    .B(_7342_),
    .C(_7163_),
    .Y(_7343_)
);

OAI21X1 _12750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11549_),
    .B(_11560_),
    .C(_9707_),
    .Y(_11571_)
);

AOI21X1 _12330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4215_),
    .B(_5771_),
    .C(_5749_),
    .Y(_6966_)
);

FILL SFILL69400x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39160x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3333_),
    .B(_3332_),
    .C(_3323_),
    .Y(_3334_)
);

XOR2X1 _13535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2872_),
    .B(_2873_),
    .Y(_2874_)
);

AOI21X1 _13115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1914_),
    .B(_2066_),
    .C(_2412_),
    .Y(_2413_)
);

XOR2X1 _23633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2025_),
    .B(_2002_),
    .Y(_2026_)
);

XNOR2X1 _23213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1562_),
    .Y(_1568_)
);

NAND3X1 _18993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8849_),
    .B(_8850_),
    .C(_8482_),
    .Y(_8855_)
);

AOI21X1 _18573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7987_),
    .B(_7989_),
    .C(_8393_),
    .Y(_8394_)
);

AND2X2 _18153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_25_bF$buf0),
    .Y(_7934_)
);

FILL SFILL69320x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10775_),
    .B(_10776_),
    .C(_10773_),
    .Y(_10789_)
);

OAI21X1 _20338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10323_),
    .B(_10328_),
    .C(_9989_),
    .Y(_10329_)
);

NAND3X1 _19778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9712_),
    .B(_9713_),
    .C(_9714_),
    .Y(_9715_)
);

NAND2X1 _19358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9254_),
    .B(_9249_),
    .Y(_9255_)
);

OAI21X1 _14493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf1),
    .B(_2465__bF$buf2),
    .C(_3916_),
    .Y(_3923_)
);

NOR3X1 _14073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3456_),
    .B(_3455_),
    .C(_3452_),
    .Y(_3463_)
);

NOR2X1 _12806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_166_),
    .B(_264_),
    .Y(_275_)
);

NAND3X1 _22904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .B(_1220_),
    .C(_1224_),
    .Y(_1232_)
);

NAND3X1 _15698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5240_),
    .B(_5239_),
    .C(_5238_),
    .Y(_5241_)
);

NAND3X1 _15278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4777_),
    .B(_4781_),
    .C(_4780_),
    .Y(_4782_)
);

FILL SFILL59320x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9394_),
    .B(_10056_),
    .C(_9761_),
    .D(_9758_),
    .Y(_10058_)
);

FILL SFILL59240x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11372_),
    .Y(_11379_)
);

NAND3X1 _17844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7573_),
    .B(_7582_),
    .C(_7585_),
    .Y(_7595_)
);

NAND3X1 _17424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7093_),
    .B(_7134_),
    .C(_7129_),
    .Y(_7135_)
);

OAI21X1 _17004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6667_),
    .B(_6668_),
    .C(_6669_),
    .Y(_6674_)
);

OAI21X1 _18629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8443_),
    .B(_8447_),
    .C(_8449_),
    .Y(_8455_)
);

NAND3X1 _18209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7955_),
    .B(_7979_),
    .C(_7984_),
    .Y(_7995_)
);

FILL FILL74200x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3106_),
    .B(_3109_),
    .C(_3113_),
    .Y(_3124_)
);

INVX1 _23862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .Y(_2272_)
);

NAND2X1 _13344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_15_bF$buf3),
    .Y(_2665_)
);

XOR2X1 _23442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .B(_1808_),
    .Y(_1818_)
);

NAND2X1 _23022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1345_),
    .Y(_1360_)
);

NAND3X1 _14969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4440_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4443_)
);

NOR3X1 _14549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3683_),
    .B(_3691_),
    .C(_3688_),
    .Y(_3984_)
);

NAND2X1 _14129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3286_),
    .B(_3291_),
    .Y(_3523_)
);

INVX2 _15910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5473_),
    .Y(_5474_)
);

NAND2X1 _18382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8179_),
    .B(_8184_),
    .Y(_8185_)
);

AOI21X1 _20987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11028_),
    .B(_11027_),
    .C(_11024_),
    .Y(_11039_)
);

INVX2 _20567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10557_),
    .Y(_10580_)
);

NAND2X1 _20147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf3),
    .B(areg_20_bF$buf1),
    .Y(_10119_)
);

AOI21X1 _19587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9504_),
    .B(_9505_),
    .C(_9490_),
    .Y(_9506_)
);

AND2X2 _19167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf4),
    .B(areg_20_bF$buf0),
    .Y(_9045_)
);

FILL SFILL69400x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_8555_),
    .Y(_10090_)
);

NAND3X1 _22713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .B(_1022_),
    .C(_1017_),
    .Y(_1023_)
);

NAND2X1 _15087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4571_),
    .B(_4572_),
    .Y(_4573_)
);

FILL SFILL69000x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _23918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[36]),
    .Y(y[36])
);

FILL SFILL74280x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf2),
    .B(areg_16_bF$buf1),
    .Y(_7385_)
);

FILL SFILL13960x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_6925_)
);

FILL SFILL74200x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_24_bF$buf1),
    .Y(_8706_)
);

OAI21X1 _18438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8241_),
    .B(_8242_),
    .C(_8245_),
    .Y(_8246_)
);

INVX1 _18018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7784_),
    .Y(_7785_)
);

AOI21X1 _13993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3369_),
    .B(_3370_),
    .C(_3362_),
    .Y(_3375_)
);

OAI21X1 _13573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2907_),
    .B(_2906_),
    .C(_2903_),
    .Y(_2916_)
);

XNOR2X1 _13153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2450_),
    .Y(_2456_)
);

AOI21X1 _23671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2017_),
    .C(_2020_),
    .Y(_2067_)
);

NOR2X1 _23251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1602_),
    .Y(_1610_)
);

AOI21X1 _14778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3971_),
    .B(_3976_),
    .C(_3956_),
    .Y(_4234_)
);

OAI21X1 _14358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3516_),
    .B(_3772_),
    .C(_3771_),
    .Y(_3773_)
);

DFFPOSX1 _24036_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[26]),
    .CLK(clk_bF$buf6),
    .D(a[26])
);

FILL SFILL64200x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7970_),
    .B(_7966_),
    .Y(_7976_)
);

NAND2X1 _20796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_21_bF$buf0),
    .Y(_10831_)
);

AOI21X1 _20376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10008_),
    .B(_10012_),
    .C(_10016_),
    .Y(_10370_)
);

NAND3X1 _16924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6572_),
    .B(_6576_),
    .C(_6578_),
    .Y(_6586_)
);

OAI21X1 _16504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6117_),
    .B(_6118_),
    .C(_6115_),
    .Y(_6125_)
);

OAI21X1 _19396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9295_),
    .B(_9294_),
    .C(_9285_),
    .Y(_9296_)
);

AND2X2 _17709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_21_bF$buf2),
    .Y(_7446_)
);

NOR3X1 _12844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_648_),
    .B(_484_),
    .C(_637_),
    .Y(_692_)
);

OAI21X1 _12424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7975_),
    .B(_7986_),
    .C(_7964_),
    .Y(_7997_)
);

NOR2X1 _22942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf0),
    .B(_6815__bF$buf4),
    .Y(_1273_)
);

NAND2X1 _12004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_6_bF$buf2),
    .Y(_3394_)
);

OAI21X1 _22522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_806_),
    .C(_800_),
    .Y(_814_)
);

OAI21X1 _22102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_94_),
    .C(_173_),
    .Y(_354_)
);

NAND2X1 _13629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_),
    .B(_2969_),
    .Y(_2976_)
);

NAND3X1 _13209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .B(_2361_),
    .C(_2513_),
    .Y(_2517_)
);

AOI21X1 _23727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2041_),
    .B(_2062_),
    .C(_2095_),
    .Y(_2127_)
);

NAND2X1 _23307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .B(_1569_),
    .Y(_1670_)
);

NAND3X1 _17882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7202_),
    .B(_7634_),
    .C(_7636_),
    .Y(_7637_)
);

NAND3X1 _17462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7174_),
    .B(_7175_),
    .C(_7173_),
    .Y(_7176_)
);

NAND3X1 _17042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6708_),
    .B(_6715_),
    .C(_6693_),
    .Y(_6716_)
);

OAI21X1 _18667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf1),
    .B(_5668__bF$buf3),
    .C(_8094_),
    .Y(_8496_)
);

NAND3X1 _18247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8030_),
    .B(_8031_),
    .C(_8028_),
    .Y(_8036_)
);

NAND2X1 _13382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_2706_),
    .Y(_2707_)
);

OAI21X1 _23480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1857_),
    .B(_1858_),
    .C(_1856_),
    .Y(_1859_)
);

NAND2X1 _23060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .B(_1399_),
    .Y(_1400_)
);

FILL SFILL44120x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3735_),
    .B(_3590_),
    .C(_3740_),
    .Y(_4026_)
);

NAND3X1 _14167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3562_),
    .B(_3563_),
    .C(_3564_),
    .Y(_3565_)
);

FILL SFILL74280x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10153_),
    .B(_10154_),
    .C(_10146_),
    .Y(_10161_)
);

NAND3X1 _16733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6375_),
    .B(_6376_),
    .C(_6373_),
    .Y(_6377_)
);

INVX1 _16313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5916_),
    .Y(_5917_)
);

FILL SFILL13560x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7232_),
    .B(_7256_),
    .C(_7254_),
    .Y(_7697_)
);

INVX2 _17518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7235_),
    .Y(_7236_)
);

NOR2X1 _12653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf2),
    .B(_5420__bF$buf2),
    .Y(_10507_)
);

NAND2X1 _12233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5804_),
    .B(_5848_),
    .Y(_5903_)
);

AOI21X1 _22751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1027_),
    .B(_1032_),
    .C(_1063_),
    .Y(_1065_)
);

NAND3X1 _22331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_597_),
    .C(_592_),
    .Y(_605_)
);

NAND3X1 _13858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3226_),
    .B(_3227_),
    .C(_3225_),
    .Y(_3228_)
);

NAND2X1 _13438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .B(_2766_),
    .Y(_2767_)
);

DFFPOSX1 _23956_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[10]),
    .CLK(clk_bF$buf2),
    .D(_0_[10])
);

AND2X2 _13018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2120_),
    .Y(_2313_)
);

OAI21X1 _23536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(_1825_),
    .C(_1822_),
    .Y(_1920_)
);

INVX1 _23116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .Y(_1462_)
);

FILL SFILL33800x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7058_),
    .B(_7056_),
    .C(_7425_),
    .Y(_7427_)
);

NAND2X1 _17271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_6967_)
);

NAND2X1 _18896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8743_),
    .B(_8747_),
    .Y(_8748_)
);

XNOR2X1 _18476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8287_),
    .B(_8285_),
    .Y(_8288_)
);

NAND3X1 _18056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7822_),
    .B(_7826_),
    .C(_7824_),
    .Y(_7827_)
);

AOI21X1 _13191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2493_),
    .C(_2491_),
    .Y(_2498_)
);

INVX8 _11924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .Y(_2519_)
);

NAND3X1 _21602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11710_),
    .B(_11711_),
    .C(_11713_),
    .Y(_11714_)
);

NAND3X1 _14396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3811_),
    .B(_3815_),
    .C(_3814_),
    .Y(_3816_)
);

NOR3X1 _12709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11099_),
    .B(_11110_),
    .C(_11066_),
    .Y(_11121_)
);

AND2X2 _22807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1110_),
    .B(_1124_),
    .Y(_1125_)
);

AOI21X1 _16962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6616_),
    .B(_6614_),
    .C(_6612_),
    .Y(_6628_)
);

INVX1 _16542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6166_),
    .Y(_6167_)
);

NAND3X1 _16122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5704_),
    .C(_5706_),
    .Y(_5707_)
);

NAND2X1 _21199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11259_),
    .B(_11262_),
    .Y(_11273_)
);

NAND2X1 _17747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_23_bF$buf2),
    .Y(_7488_)
);

AND2X2 _17327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_20_bF$buf2),
    .Y(_7027_)
);

AOI21X1 _12882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11373_),
    .B(_11384_),
    .C(_11361_),
    .Y(_1107_)
);

NOR2X1 _12462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8391_),
    .B(_8402_),
    .Y(_8413_)
);

AOI21X1 _22980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1199_),
    .B(_1212_),
    .C(_1312_),
    .Y(_1313_)
);

NOR2X1 _12042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3591_),
    .B(_3679_),
    .Y(_3810_)
);

OAI21X1 _22560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_627_),
    .B(_852_),
    .C(_854_),
    .Y(_855_)
);

NAND3X1 _22140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_395_)
);

FILL SFILL8680x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3015_),
    .B(_3016_),
    .C(_3017_),
    .Y(_3018_)
);

NAND2X1 _13247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg_16_bF$buf1),
    .Y(_2558_)
);

OAI21X1 _23765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2166_),
    .B(_2145_),
    .C(_2167_),
    .Y(_2168_)
);

NOR2X1 _23345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .B(_1711_),
    .Y(_1712_)
);

FILL SFILL8600x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6512_),
    .B(_6598_),
    .C(_6597_),
    .Y(_6757_)
);

NAND2X1 _15813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5072_),
    .B(_5079_),
    .Y(_5368_)
);

OAI21X1 _18285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7780_),
    .B(_8077_),
    .C(_8030_),
    .Y(_8078_)
);

FILL SFILL43800x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .C(_55_),
    .Y(_57_)
);

NAND3X1 _21411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11503_),
    .B(_11504_),
    .C(_11502_),
    .Y(_11506_)
);

FILL SFILL38840x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1631_),
    .Y(_1718_)
);

XNOR2X1 _12518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9016_),
    .B(_8972_),
    .Y(_9027_)
);

AND2X2 _22616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_714_),
    .B(_492_),
    .Y(_917_)
);

FILL SFILL33800x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6042_),
    .B(_6416_),
    .C(_6412_),
    .Y(_6418_)
);

AOI21X1 _16351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5941_),
    .B(_5948_),
    .C(_5928_),
    .Y(_5959_)
);

BUFX2 BUFX2_insert350 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104_),
    .Y(_9104__bF$buf1)
);

BUFX2 BUFX2_insert351 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104_),
    .Y(_9104__bF$buf0)
);

BUFX2 BUFX2_insert352 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf4)
);

BUFX2 BUFX2_insert353 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf3)
);

AOI21X1 _17976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7732_),
    .B(_7734_),
    .C(_7731_),
    .Y(_7739_)
);

BUFX2 BUFX2_insert354 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf2)
);

NAND2X1 _17556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_25_bF$buf5),
    .Y(_7278_)
);

BUFX2 BUFX2_insert355 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf1)
);

BUFX2 BUFX2_insert356 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(breg_12_bF$buf0)
);

NOR2X1 _17136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6051_),
    .B(_6430_),
    .Y(_6818_)
);

BUFX2 BUFX2_insert357 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf6)
);

BUFX2 BUFX2_insert358 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf5)
);

NOR2X1 _12691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10836_),
    .B(_10847_),
    .Y(_10924_)
);

BUFX2 BUFX2_insert359 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf4)
);

OAI21X1 _12271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6253_),
    .B(_6242_),
    .C(_6198_),
    .Y(_6319_)
);

FILL SFILL54200x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf1),
    .B(_2763_),
    .C(_3268_),
    .Y(_3269_)
);

OAI21X1 _13476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2801_),
    .B(_2807_),
    .C(_2808_),
    .Y(_2809_)
);

DFFPOSX1 _23994_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[48]),
    .CLK(clk_bF$buf6),
    .D(_0_[48])
);

AOI21X1 _23574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3234_),
    .B(_3237_),
    .C(_3498_),
    .Y(_1961_)
);

AOI21X1 _13056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2340_),
    .C(_1173_),
    .Y(_2351_)
);

AOI21X1 _23154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1494_),
    .C(_1503_),
    .Y(_1504_)
);

INVX1 _19702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9265_),
    .Y(_9632_)
);

OAI21X1 _15622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3402__bF$buf2),
    .C(_5151_),
    .Y(_5159_)
);

INVX1 _15202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .Y(_4699_)
);

NAND3X1 _18094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7848_),
    .B(_7816_),
    .C(_7855_),
    .Y(_7869_)
);

NOR3X1 _20699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10723_),
    .B(_10719_),
    .C(_10722_),
    .Y(_10724_)
);

NOR2X1 _20279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10261_),
    .B(_10263_),
    .Y(_10264_)
);

OAI21X1 _16827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6475_),
    .B(_6476_),
    .C(_6478_),
    .Y(_6479_)
);

AOI21X1 _16407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6003_),
    .B(_6009_),
    .C(_5667_),
    .Y(_6019_)
);

INVX1 _11962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2781_),
    .Y(_2935_)
);

OAI21X1 _21640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11480_),
    .B(_11754_),
    .C(_11482_),
    .Y(_11755_)
);

AOI21X1 _21220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11295_),
    .B(_11290_),
    .C(_11007_),
    .Y(_11296_)
);

NAND3X1 _19299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9134_),
    .B(_9136_),
    .C(_9130_),
    .Y(_9190_)
);

NAND3X1 _12747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9948_),
    .B(_11527_),
    .C(_11494_),
    .Y(_11538_)
);

AOI21X1 _12327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6780_),
    .B(_6823_),
    .C(_6110_),
    .Y(_6933_)
);

AOI21X1 _22845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_981_),
    .B(_1003_),
    .C(_1006_),
    .Y(_1167_)
);

AOI22X1 _22425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_707_),
    .C(_490_),
    .D(_488_),
    .Y(_708_)
);

NAND2X1 _22005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_87_),
    .Y(_247_)
);

AOI21X1 _16580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6199_),
    .B(_6192_),
    .C(_6161_),
    .Y(_6208_)
);

INVX2 _16160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5747_),
    .Y(_5748_)
);

INVX1 _17785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7529_),
    .Y(_7530_)
);

AND2X2 _17365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .B(areg_24_bF$buf3),
    .Y(_7070_)
);

NOR2X1 _12080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4193_),
    .B(_4215_),
    .Y(_4226_)
);

OAI21X1 _20911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10956_),
    .B(_10952_),
    .C(_10813_),
    .Y(_10958_)
);

FILL SFILL38840x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _13285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2598_),
    .B(_2595_),
    .Y(_2599_)
);

OAI21X1 _23383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1629_),
    .B(_1553_),
    .C(_1632_),
    .Y(_1754_)
);

FILL SFILL28920x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9876_),
    .B(_9882_),
    .C(_9860_),
    .Y(_9884_)
);

OAI21X1 _19511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9420_),
    .B(_9421_),
    .C(_9419_),
    .Y(_9423_)
);

INVX1 _15851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5408_),
    .Y(_5410_)
);

AOI21X1 _15431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4350_),
    .B(_4624_),
    .C(_4949_),
    .Y(_4951_)
);

OAI21X1 _15011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4488_),
    .B(_4484_),
    .C(_4448_),
    .Y(_4490_)
);

FILL SFILL28840x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf3),
    .B(_5315__bF$buf4),
    .C(_10047_),
    .Y(_10054_)
);

AND2X2 _16636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .B(areg_22_bF$buf0),
    .Y(_6270_)
);

NAND3X1 _16216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5805_),
    .B(_5780_),
    .C(_5809_),
    .Y(_5810_)
);

NAND2X1 _12976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2120_),
    .Y(_2131_)
);

AOI21X1 _12556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9389_),
    .B(_9400_),
    .C(_9378_),
    .Y(_9444_)
);

NAND3X1 _12136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .B(_4796_),
    .C(_4829_),
    .Y(_4840_)
);

OAI21X1 _22654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_747_),
    .C(_749_),
    .Y(_958_)
);

NAND2X1 _22234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_360_),
    .Y(_498_)
);

OAI21X1 _23859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2267_),
    .B(_2246_),
    .C(_2266_),
    .Y(_2268_)
);

OAI21X1 _23439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1703_),
    .B(_1811_),
    .C(_1813_),
    .Y(_1814_)
);

XOR2X1 _23019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1351_),
    .B(_1355_),
    .Y(_1356_)
);

NAND3X1 _14702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4147_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4151_)
);

OAI21X1 _17594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7318_),
    .B(_7319_),
    .C(_7317_),
    .Y(_7320_)
);

NOR2X1 _17174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6849_),
    .B(_6857_),
    .Y(_6860_)
);

FILL SFILL44200x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _15907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .B(_5467_),
    .Y(_5471_)
);

NOR2X1 _20720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10745_),
    .B(_10746_),
    .Y(_10747_)
);

AOI21X1 _20300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10285_),
    .B(_10286_),
    .C(_10279_),
    .Y(_10287_)
);

AND2X2 _18799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf2),
    .B(areg_19_bF$buf5),
    .Y(_8641_)
);

NAND3X1 _18379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8177_),
    .B(_8171_),
    .C(_8167_),
    .Y(_8181_)
);

INVX2 _13094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .Y(_2391_)
);

OAI21X1 _23192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .B(_1540_),
    .C(_1544_),
    .Y(_1545_)
);

OAI21X1 _19740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9669_),
    .B(_9670_),
    .C(_9666_),
    .Y(_9673_)
);

NOR3X1 _19320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8794_),
    .B(_8801_),
    .C(_8804_),
    .Y(_9213_)
);

FILL SFILL69080x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_154_),
    .C(_126_),
    .Y(_160_)
);

NOR2X1 _21505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf1),
    .B(_6815__bF$buf0),
    .Y(_11608_)
);

NAND2X1 _14299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3708_),
    .B(_3709_),
    .Y(_3710_)
);

INVX2 _15660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5199_),
    .Y(_5200_)
);

AOI21X1 _15240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4391_),
    .B(_4413_),
    .C(_4416_),
    .Y(_4740_)
);

FILL SFILL38920x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_18_bF$buf0),
    .Y(_6521_)
);

NAND2X1 _16445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_26_bF$buf0),
    .Y(_6060_)
);

OAI21X1 _16025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .B(_5499_),
    .C(_5506_),
    .Y(_5601_)
);

FILL SFILL69320x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11898_),
    .B(_11887_),
    .C(_11876_),
    .Y(_45_)
);

OAI21X1 _12365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf2),
    .B(_5453__bF$buf5),
    .C(_6143_),
    .Y(_7349_)
);

NAND2X1 _22883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1207_),
    .B(_1205_),
    .Y(_1209_)
);

NAND2X1 _22463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .B(_748_),
    .Y(_749_)
);

OAI21X1 _22043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_288_),
    .B(_283_),
    .C(_252_),
    .Y(_289_)
);

FILL SFILL28920x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2041_),
    .B(_2062_),
    .Y(_2063_)
);

NAND3X1 _23248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1605_),
    .C(_1572_),
    .Y(_1606_)
);

NOR2X1 _14931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4397_),
    .B(_4400_),
    .Y(_4402_)
);

NOR3X1 _14511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3936_),
    .B(_3938_),
    .C(_3935_),
    .Y(_3943_)
);

AOI21X1 _15716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5242_),
    .B(_5248_),
    .C(_5101_),
    .Y(_5262_)
);

NOR2X1 _18188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7970_),
    .B(_7966_),
    .Y(_7972_)
);

OAI21X1 _21734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11854_),
    .B(_11858_),
    .C(_11596_),
    .Y(_11859_)
);

OAI21X1 _21314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11138_),
    .B(_11159_),
    .C(_11163_),
    .Y(_11399_)
);

NAND3X1 _22939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1116_),
    .B(_1121_),
    .C(_1112_),
    .Y(_1269_)
);

NAND3X1 _22519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_809_),
    .C(_802_),
    .Y(_810_)
);

FILL SFILL18600x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_28_bF$buf4),
    .Y(_6312_)
);

OAI22X1 _16254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_3146__bF$buf1),
    .C(_7217__bF$buf3),
    .D(_2884__bF$buf1),
    .Y(_5852_)
);

NAND3X1 _17879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7218_),
    .B(_7629_),
    .C(_7632_),
    .Y(_7633_)
);

NAND2X1 _17459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7171_),
    .B(_7172_),
    .Y(_7173_)
);

AOI21X1 _17039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6710_),
    .B(_6711_),
    .C(_6695_),
    .Y(_6712_)
);

NAND3X1 _12594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8478_),
    .B(_9795_),
    .C(_9806_),
    .Y(_9861_)
);

NOR2X1 _12174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5245_),
    .B(_5212_),
    .Y(_5256_)
);

INVX1 _22692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_848_),
    .Y(_1000_)
);

AND2X2 _22272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .B(_539_),
    .Y(_540_)
);

OAI21X1 _18820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8655_),
    .B(_8656_),
    .C(_8652_),
    .Y(_8664_)
);

NAND2X1 _18400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8200_),
    .B(_8198_),
    .Y(_8204_)
);

FILL SFILL69080x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3157_),
    .B(_3158_),
    .C(_3162_),
    .Y(_3163_)
);

NAND3X1 _13379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .B(_2702_),
    .C(_2625_),
    .Y(_2703_)
);

BUFX2 _23897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[15]),
    .Y(y[15])
);

INVX1 _23477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .Y(_1856_)
);

XNOR2X1 _23057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1261_),
    .B(_1397_),
    .Y(_0_[50])
);

OAI21X1 _19605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9518_),
    .B(_9519_),
    .C(_9516_),
    .Y(_9526_)
);

AOI21X1 _14740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .B(_3939_),
    .C(_3943_),
    .Y(_4192_)
);

OAI21X1 _14320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3731_),
    .B(_3732_),
    .C(_3638_),
    .Y(_3733_)
);

OAI21X1 _15945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5512_),
    .B(_5224_),
    .C(_5217_),
    .Y(_5513_)
);

OAI21X1 _15525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf0),
    .B(_2560__bF$buf4),
    .C(_5048_),
    .Y(_5052_)
);

NOR3X1 _15105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4284_),
    .B(_4285_),
    .C(_4283_),
    .Y(_4593_)
);

AOI21X1 _21963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_185_),
    .C(_11829_),
    .Y(_202_)
);

OAI21X1 _21543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11372_),
    .B(_11377_),
    .C(_11380_),
    .Y(_11649_)
);

AOI21X1 _21123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10933_),
    .B(_11189_),
    .C(_11188_),
    .Y(_11190_)
);

NAND2X1 _22748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1058_),
    .Y(_1061_)
);

OAI21X1 _22328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_600_),
    .C(_433_),
    .Y(_601_)
);

FILL SFILL49080x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6096_),
    .B(_6057_),
    .C(_6101_),
    .Y(_6102_)
);

NOR3X1 _16063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5638_),
    .B(_5639_),
    .C(_5635_),
    .Y(_5643_)
);

FILL SFILL49000x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7417_),
    .B(_7418_),
    .C(_7416_),
    .Y(_7423_)
);

AND2X2 _17268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_6963_)
);

NAND2X1 _22081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_118_),
    .Y(_331_)
);

FILL SFILL39000x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_10851_)
);

NAND3X1 _13188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2493_),
    .C(_2491_),
    .Y(_2494_)
);

NOR3X1 _23286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1634_),
    .C(_1636_),
    .Y(_1648_)
);

OAI21X1 _19834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9776_),
    .B(_9775_),
    .C(_9766_),
    .Y(_9777_)
);

NAND3X1 _19414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9278_),
    .B(_9315_),
    .C(_9314_),
    .Y(_9316_)
);

FILL SFILL8760x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5282_),
    .B(_5280_),
    .C(_5270_),
    .Y(_5303_)
);

OAI21X1 _15334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4842_),
    .B(_4843_),
    .C(_4816_),
    .Y(_4844_)
);

OAI21X1 _16959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf1),
    .B(_3402__bF$buf0),
    .C(_6613_),
    .Y(_6624_)
);

INVX1 _16539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5786_),
    .Y(_6163_)
);

OAI21X1 _16119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5695_),
    .B(_5696_),
    .C(_5689_),
    .Y(_5703_)
);

AND2X2 _21772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_27_bF$buf4),
    .Y(_11900_)
);

NAND2X1 _21352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf1),
    .B(breg_23_bF$buf0),
    .Y(_11441_)
);

OAI21X1 _17900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7259_),
    .B(_7227_),
    .C(_7268_),
    .Y(_7655_)
);

FILL SFILL19080x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL4040x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_911_),
    .B(_954_),
    .C(_976_),
    .Y(_1075_)
);

XNOR2X1 _12459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8370_),
    .B(_8359_),
    .Y(_0_[10])
);

XNOR2X1 _22977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1309_),
    .B(_1308_),
    .Y(_1310_)
);

NAND2X1 _12039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2781_),
    .B(_2913_),
    .Y(_3787_)
);

NAND2X1 _22557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_29_bF$buf1),
    .Y(_852_)
);

FILL SFILL3720x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _22137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_372_),
    .C(_387_),
    .Y(_392_)
);

FILL SFILL43960x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(_3175_),
    .C(_3128_),
    .Y(_3186_)
);

AOI21X1 _13400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2711_),
    .B(_2717_),
    .C(_2577_),
    .Y(_2726_)
);

NAND2X1 _16292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5891_),
    .B(_5893_),
    .Y(_5894_)
);

OAI21X1 _14605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4041_),
    .B(_4044_),
    .C(_3767_),
    .Y(_4045_)
);

XNOR2X1 _17497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6808_),
    .B(_7213_),
    .Y(_0_[30])
);

AOI21X1 _17077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6735_),
    .B(_6741_),
    .C(_6648_),
    .Y(_6754_)
);

NOR3X1 _20623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10302_),
    .B(_10303_),
    .C(_10301_),
    .Y(_10642_)
);

NAND3X1 _20203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10180_),
    .B(_10141_),
    .C(_10173_),
    .Y(_10181_)
);

NAND2X1 _23095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1299_),
    .B(_1310_),
    .Y(_1439_)
);

NAND2X1 _19643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9567_),
    .B(_9562_),
    .Y(_9568_)
);

NAND2X1 _19223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_26_bF$buf3),
    .Y(_9107_)
);

NAND3X1 _21828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_51_),
    .C(_52_),
    .Y(_53_)
);

AOI21X1 _21408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11169_),
    .B(_11191_),
    .C(_11194_),
    .Y(_11502_)
);

OAI21X1 _15983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5195_),
    .B(_5199_),
    .C(_5198_),
    .Y(_5555_)
);

AOI21X1 _15563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4769_),
    .B(_4809_),
    .C(_4805_),
    .Y(_5094_)
);

OAI21X1 _15143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4633_),
    .B(_4634_),
    .C(_4631_),
    .Y(_4635_)
);

NAND3X1 _16768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6413_),
    .B(_6021_),
    .C(_6414_),
    .Y(_6415_)
);

NOR3X1 _16348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5569_),
    .B(_5568_),
    .C(_5570_),
    .Y(_5955_)
);

NAND3X1 _21581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11685_),
    .B(_11647_),
    .C(_11689_),
    .Y(_11691_)
);

OAI21X1 _21161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11229_),
    .B(_7520__bF$buf3),
    .C(_11230_),
    .Y(_11232_)
);

FILL SFILL39000x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10825_),
    .B(_10880_),
    .C(_10858_),
    .Y(_10891_)
);

NAND3X1 _12268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6121_),
    .B(_6275_),
    .C(_6209_),
    .Y(_6286_)
);

NAND2X1 _22786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .B(_1027_),
    .Y(_1102_)
);

NAND2X1 _22366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf2),
    .B(areg_29_bF$buf1),
    .Y(_643_)
);

AOI21X1 _18914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8750_),
    .B(_8754_),
    .C(_8755_),
    .Y(_8768_)
);

FILL FILL73960x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3990_),
    .B(_3996_),
    .C(_4000_),
    .Y(_4296_)
);

AOI21X1 _14414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3816_),
    .B(_3819_),
    .C(_3824_),
    .Y(_3836_)
);

FILL SFILL53960x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_18_bF$buf4),
    .Y(_5155_)
);

FILL SFILL74040x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10883_),
    .B(_10876_),
    .C(_10881_),
    .Y(_10893_)
);

NOR3X1 _20432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10425_),
    .B(_10426_),
    .C(_10427_),
    .Y(_10432_)
);

NAND3X1 _20012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9967_),
    .B(_9968_),
    .C(_9639_),
    .Y(_9972_)
);

NAND3X1 _19872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9800_),
    .B(_9803_),
    .C(_9813_),
    .Y(_9819_)
);

AOI21X1 _19452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9342_),
    .B(_9347_),
    .C(_9348_),
    .Y(_9358_)
);

INVX2 _19032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8896_),
    .Y(_8897_)
);

INVX1 _11959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2803_),
    .Y(_2902_)
);

FILL SFILL3720x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11482_),
    .B(_11486_),
    .C(_11493_),
    .Y(_11752_)
);

NAND3X1 _21217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11010_),
    .B(_11287_),
    .C(_11288_),
    .Y(_11293_)
);

XNOR2X1 _12900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1228_),
    .Y(_0_[13])
);

NAND3X1 _15792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(_5336_),
    .C(_5341_),
    .Y(_5345_)
);

NAND3X1 _15372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4816_),
    .B(_4839_),
    .C(_4834_),
    .Y(_4886_)
);

AOI21X1 _16997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6660_),
    .B(_6664_),
    .C(_6665_),
    .Y(_6666_)
);

OAI21X1 _16577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5873_),
    .B(_5879_),
    .C(_5882_),
    .Y(_6205_)
);

OAI21X1 _16157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5616_),
    .B(_5744_),
    .C(_5606_),
    .Y(_5745_)
);

NAND3X1 _21390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11477_),
    .B(_11481_),
    .C(_11479_),
    .Y(_11482_)
);

FILL SFILL64360x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8742_),
    .Y(_8797_)
);

NOR2X1 _12077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4149_),
    .B(_4182_),
    .Y(_4193_)
);

NAND2X1 _22595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_893_),
    .B(_688_),
    .Y(_894_)
);

INVX1 _22175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .Y(_434_)
);

AOI21X1 _18723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8210_),
    .B(_8214_),
    .C(_8196_),
    .Y(_8558_)
);

OAI21X1 _18303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8097_),
    .B(_8096_),
    .C(_8087_),
    .Y(_8098_)
);

AOI21X1 _20908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10897_),
    .B(_10903_),
    .C(_10815_),
    .Y(_10954_)
);

AOI21X1 _19928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9878_),
    .B(_9879_),
    .C(_9863_),
    .Y(_9880_)
);

XNOR2X1 _19508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9397_),
    .B(_9392_),
    .Y(_9419_)
);

NAND3X1 _14643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4082_),
    .B(_4085_),
    .C(_4084_),
    .Y(_4086_)
);

OAI21X1 _14223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3625_),
    .B(_3619_),
    .C(_3626_),
    .Y(_3627_)
);

INVX1 _15848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5048_),
    .Y(_5406_)
);

OAI21X1 _15428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4945_),
    .B(_4946_),
    .C(_4652_),
    .Y(_4947_)
);

AOI21X1 _15008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4468_),
    .B(_4474_),
    .C(_4453_),
    .Y(_4486_)
);

OAI22X1 _20661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9986_),
    .B(_10678_),
    .C(_10681_),
    .D(_10675_),
    .Y(_10683_)
);

NAND2X1 _20241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf3),
    .B(areg_29_bF$buf3),
    .Y(_10222_)
);

OAI21X1 _19681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9605_),
    .B(_9608_),
    .C(_9272_),
    .Y(_9610_)
);

NAND2X1 _19261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_29_bF$buf3),
    .Y(_9149_)
);

NAND2X1 _21866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_23_bF$buf0),
    .Y(_95_)
);

OAI21X1 _21446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11543_),
    .B(_11542_),
    .C(_11539_),
    .Y(_11544_)
);

NAND3X1 _21026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11060_),
    .B(_11075_),
    .C(_11082_),
    .Y(_11083_)
);

FILL SFILL74200x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4602_),
    .B(_4674_),
    .C(_4592_),
    .Y(_4676_)
);

FILL SFILL13880x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3273_),
    .B(_3278_),
    .C(_3260_),
    .Y(_3289_)
);

NAND3X1 _16386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5988_),
    .B(_5995_),
    .C(_5745_),
    .Y(_5996_)
);

FILL SFILL13800x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8756_),
    .B(_8762_),
    .C(_8744_),
    .Y(_8810_)
);

AOI21X1 _18532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8343_),
    .B(_8344_),
    .C(_8335_),
    .Y(_8350_)
);

NAND2X1 _18112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf2),
    .B(areg_21_bF$buf2),
    .Y(_7889_)
);

NAND2X1 _20717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_26_bF$buf3),
    .Y(_10744_)
);

INVX1 _23189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1398_),
    .Y(_1541_)
);

AOI21X1 _19737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9658_),
    .B(_9657_),
    .C(_9654_),
    .Y(_9670_)
);

OAI21X1 _19317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9188_),
    .B(_9196_),
    .C(_9198_),
    .Y(_9210_)
);

NAND3X1 _14872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .B(_4043_),
    .C(_4337_),
    .Y(_4338_)
);

OAI21X1 _14452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf0),
    .B(_9104__bF$buf2),
    .C(_3877_),
    .Y(_3878_)
);

OAI21X1 _14032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3415_),
    .B(_3417_),
    .C(_3412_),
    .Y(_3418_)
);

AND2X2 _15657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_25_bF$buf2),
    .Y(_5197_)
);

AOI21X1 _15237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4718_),
    .B(_4722_),
    .C(_4725_),
    .Y(_4737_)
);

XNOR2X1 _20890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10914_),
    .B(_10933_),
    .Y(_10934_)
);

AND2X2 _20470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf2),
    .B(areg_20_bF$buf1),
    .Y(_10473_)
);

OAI21X1 _20050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf0),
    .B(_5668__bF$buf4),
    .C(_9660_),
    .Y(_10012_)
);

OAI21X1 _19490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9025_),
    .B(_9015_),
    .C(_9020_),
    .Y(_9399_)
);

NAND2X1 _19070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_25_bF$buf5),
    .Y(_8938_)
);

NAND2X1 _11997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3296_),
    .B(_3307_),
    .Y(_3318_)
);

NAND3X1 _21675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11751_),
    .B(_11785_),
    .C(_11793_),
    .Y(_11794_)
);

NAND2X1 _21255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf2),
    .B(breg_29_bF$buf4),
    .Y(_11334_)
);

NAND3X1 _17803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7540_),
    .B(_7542_),
    .C(_7535_),
    .Y(_7550_)
);

FILL SFILL54040x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3075_),
    .B(_3074_),
    .C(_3060_),
    .Y(_3080_)
);

NAND3X1 _13303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2580_),
    .B(_2619_),
    .C(_2612_),
    .Y(_2620_)
);

OAI21X1 _23821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9153_),
    .B(_7225__bF$buf1),
    .C(_2227_),
    .Y(_2229_)
);

INVX1 _23401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1771_),
    .Y(_1773_)
);

AND2X2 _16195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_15_bF$buf3),
    .Y(_5786_)
);

OAI21X1 _14928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf0),
    .B(_2362__bF$buf5),
    .C(_4397_),
    .Y(_4398_)
);

OAI21X1 _14508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3935_),
    .B(_3936_),
    .C(_3938_),
    .Y(_3939_)
);

FILL SFILL44040x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8411_),
    .B(_8412_),
    .C(_8281_),
    .Y(_8600_)
);

NAND3X1 _18341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8131_),
    .B(_8135_),
    .C(_8138_),
    .Y(_8140_)
);

NAND3X1 _20946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10691_),
    .B(_10987_),
    .C(_10983_),
    .Y(_10996_)
);

NAND3X1 _20526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10495_),
    .B(_10534_),
    .C(_10527_),
    .Y(_10535_)
);

AOI21X1 _20106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10059_),
    .B(_10064_),
    .C(_10044_),
    .Y(_10074_)
);

NAND2X1 _19966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9914_),
    .B(_9564_),
    .Y(_9921_)
);

OAI21X1 _19546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9459_),
    .B(_9460_),
    .C(_9427_),
    .Y(_9461_)
);

OAI21X1 _19126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8993_),
    .B(_8992_),
    .C(_8990_),
    .Y(_9000_)
);

AOI21X1 _14681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3831_),
    .B(_3809_),
    .C(_3835_),
    .Y(_4128_)
);

OAI21X1 _14261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3667_),
    .B(_3420_),
    .C(_3411_),
    .Y(_3669_)
);

FILL SFILL69160x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5446_),
    .B(_5445_),
    .C(_5447_),
    .Y(_5448_)
);

NOR3X1 _15466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4986_),
    .B(_4972_),
    .C(_4985_),
    .Y(_4987_)
);

FILL SFILL74120x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4527_),
    .B(_4262_),
    .C(_4253_),
    .Y(_4528_)
);

AOI21X1 _21484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11006_),
    .B(_11299_),
    .C(_11585_),
    .Y(_11586_)
);

NAND3X1 _21064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11015_),
    .B(_11118_),
    .C(_11124_),
    .Y(_11125_)
);

NAND3X1 _17612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7336_),
    .B(_7339_),
    .C(_7337_),
    .Y(_7340_)
);

FILL SFILL23720x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(_848_),
    .C(_860_),
    .Y(_996_)
);

OAI21X1 _22269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_532_),
    .C(_531_),
    .Y(_536_)
);

FILL SFILL64120x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8653_),
    .B(_8660_),
    .C(_8638_),
    .Y(_8661_)
);

NAND2X1 _13952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf0),
    .B(breg_10_bF$buf3),
    .Y(_3331_)
);

NAND2X1 _13532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf0),
    .B(areg_12_bF$buf1),
    .Y(_2871_)
);

AOI21X1 _13112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2404_),
    .C(_2403_),
    .Y(_2410_)
);

NOR2X1 _23630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2019_),
    .B(_2020_),
    .Y(_2022_)
);

NAND2X1 _23210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_25_bF$buf1),
    .B(breg_28_bF$buf3),
    .Y(_1564_)
);

FILL SFILL64040x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4183_),
    .B(_4187_),
    .C(_4188_),
    .Y(_4189_)
);

NAND3X1 _14317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3725_),
    .B(_3726_),
    .C(_3724_),
    .Y(_3730_)
);

FILL FILL74040x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8838_),
    .B(_8598_),
    .C(_8833_),
    .Y(_8850_)
);

AOI21X1 _18570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8389_),
    .B(_8388_),
    .C(_8387_),
    .Y(_8390_)
);

OAI21X1 _18150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7493_),
    .B(_7929_),
    .C(_7495_),
    .Y(_7930_)
);

FILL SFILL54120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10780_),
    .B(_10785_),
    .C(_10741_),
    .Y(_10786_)
);

AOI21X1 _20335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10319_),
    .B(_10320_),
    .C(_10318_),
    .Y(_10326_)
);

FILL SFILL18680x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _19775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9690_),
    .Y(_9712_)
);

NAND3X1 _19355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8882_),
    .B(_9245_),
    .C(_9246_),
    .Y(_9252_)
);

AND2X2 _14490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_14_bF$buf0),
    .Y(_3919_)
);

NAND3X1 _14070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3249_),
    .B(_3298_),
    .C(_3303_),
    .Y(_3459_)
);

FILL SFILL59320x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_210_),
    .Y(_242_)
);

AOI21X1 _22901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1227_),
    .C(_1068_),
    .Y(_1229_)
);

NAND2X1 _15695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5236_),
    .B(_5237_),
    .Y(_5238_)
);

AND2X2 _15275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_15_bF$buf1),
    .Y(_4779_)
);

NOR2X1 _21293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11374_),
    .B(_11375_),
    .Y(_11376_)
);

NAND3X1 _17841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7432_),
    .B(_7344_),
    .C(_7431_),
    .Y(_7592_)
);

OAI21X1 _17421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7127_),
    .B(_7126_),
    .C(_7107_),
    .Y(_7132_)
);

NOR3X1 _17001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6668_),
    .B(_6669_),
    .C(_6667_),
    .Y(_6671_)
);

OAI21X1 _22498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_786_),
    .B(_609_),
    .C(_612_),
    .Y(_787_)
);

NAND3X1 _22078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .C(_326_),
    .Y(_327_)
);

NAND3X1 _18626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8450_),
    .B(_8451_),
    .C(_8449_),
    .Y(_8452_)
);

NOR3X1 _18206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7555_),
    .B(_7556_),
    .C(_7554_),
    .Y(_7992_)
);

NAND3X1 _13761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3114_),
    .B(_3120_),
    .C(_3098_),
    .Y(_3121_)
);

INVX2 _13341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .Y(_2662_)
);

FILL SFILL38760x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4134_),
    .Y(_4440_)
);

FILL SFILL74120x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3968_),
    .C(_3970_),
    .Y(_3981_)
);

NAND2X1 _14126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3298_),
    .B(_3459_),
    .Y(_3520_)
);

OAI21X1 _20984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf1),
    .B(_6050__bF$buf2),
    .C(_11026_),
    .Y(_11036_)
);

AOI21X1 _20564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10568_),
    .B(_10566_),
    .C(_10564_),
    .Y(_10577_)
);

XNOR2X1 _20144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10115_),
    .B(_10113_),
    .Y(_10116_)
);

AOI21X1 _19584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9113_),
    .B(_9116_),
    .C(_9108_),
    .Y(_9503_)
);

AOI21X1 _19164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8229_),
    .B(_9041_),
    .C(_8655_),
    .Y(_9042_)
);

FILL SFILL59160x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_29_bF$buf4),
    .Y(_11896_)
);

FILL SFILL64120x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11436_),
    .B(_11435_),
    .C(_11434_),
    .Y(_11437_)
);

NOR2X1 _12612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8599_),
    .B(_10046_),
    .Y(_10057_)
);

OAI21X1 _22710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1015_),
    .C(_980_),
    .Y(_1019_)
);

NAND3X1 _15084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4563_),
    .B(_4526_),
    .C(_4569_),
    .Y(_4570_)
);

AOI21X1 _13817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2916_),
    .B(_2915_),
    .C(_2908_),
    .Y(_3183_)
);

BUFX2 _23915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[33]),
    .Y(y[33])
);

INVX1 _16289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5889_),
    .Y(_5890_)
);

FILL SFILL18760x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf1),
    .B(breg_17_bF$buf0),
    .Y(_7381_)
);

OAI21X1 _17230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6760_),
    .B(_6920_),
    .C(_6750_),
    .Y(_6921_)
);

FILL SFILL54120x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38760x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf2),
    .B(areg_23_bF$buf2),
    .Y(_8703_)
);

NAND2X1 _18435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_20_bF$buf0),
    .Y(_8243_)
);

OAI21X1 _18015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7781_),
    .B(_7593_),
    .C(_7583_),
    .Y(_7782_)
);

NAND3X1 _13990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3362_),
    .B(_3369_),
    .C(_3370_),
    .Y(_3371_)
);

AOI21X1 _13570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2910_),
    .B(_2911_),
    .C(_2864_),
    .Y(_2912_)
);

NOR2X1 _13150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .B(_2451_),
    .Y(_2452_)
);

AOI21X1 _14775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4213_),
    .B(_4217_),
    .C(_4221_),
    .Y(_4231_)
);

XNOR2X1 _14355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3516_),
    .B(_3770_),
    .Y(_0_[20])
);

DFFPOSX1 _24033_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[23]),
    .CLK(clk_bF$buf1),
    .D(a[23])
);

AOI21X1 _20793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10824_),
    .B(_10827_),
    .C(_10822_),
    .Y(_10828_)
);

NOR2X1 _20373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10359_),
    .B(_10360_),
    .Y(_10367_)
);

NAND3X1 _16921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6577_),
    .B(_6581_),
    .C(_6545_),
    .Y(_6583_)
);

AOI21X1 _16501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6116_),
    .B(_6120_),
    .C(_6048_),
    .Y(_6122_)
);

NAND2X1 _19393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_27_bF$buf2),
    .Y(_9293_)
);

OAI21X1 _21998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11879_),
    .B(_238_),
    .C(_237_),
    .Y(_239_)
);

NAND3X1 _21578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11671_),
    .B(_11675_),
    .C(_11683_),
    .Y(_11687_)
);

NAND2X1 _21158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf2),
    .B(areg_29_bF$buf2),
    .Y(_11228_)
);

OAI21X1 _17706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7036_),
    .B(_7025_),
    .C(_7029_),
    .Y(_7443_)
);

FILL SFILL69240x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_648_),
    .C(_484_),
    .Y(_659_)
);

NAND2X1 _12421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7942_),
    .B(_7953_),
    .Y(_7964_)
);

NOR2X1 _12001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3187_),
    .B(_3209_),
    .Y(_3361_)
);

FILL SFILL34040x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2973_),
    .B(_2969_),
    .Y(_2974_)
);

OAI21X1 _13206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2511_),
    .C(_2377_),
    .Y(_2514_)
);

NOR2X1 _23724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2067_),
    .B(_2123_),
    .Y(_2124_)
);

OAI21X1 _23304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf2),
    .B(_6427_),
    .C(_1567_),
    .Y(_1667_)
);

NAND2X1 _16098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5678_),
    .B(_5679_),
    .Y(_5680_)
);

FILL FILL74200x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg_28_bF$buf0),
    .Y(_8493_)
);

OAI21X1 _18244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8025_),
    .B(_8032_),
    .C(_7663_),
    .Y(_8033_)
);

FILL SFILL28760x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10849_),
    .B(_10888_),
    .C(_10882_),
    .Y(_10889_)
);

OAI21X1 _20429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10425_),
    .B(_10426_),
    .C(_10427_),
    .Y(_10428_)
);

NAND3X1 _20009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9642_),
    .B(_9954_),
    .C(_9960_),
    .Y(_9968_)
);

AOI21X1 _19869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9808_),
    .B(_9814_),
    .C(_9793_),
    .Y(_9815_)
);

NAND3X1 _19449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9320_),
    .B(_9353_),
    .C(_9349_),
    .Y(_9354_)
);

INVX1 _19029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8892_),
    .Y(_8893_)
);

OAI21X1 _14584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4004_),
    .B(_4011_),
    .C(_4013_),
    .Y(_4023_)
);

NOR2X1 _14164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3561_),
    .B(_3276_),
    .Y(_3562_)
);

FILL FILL74120x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5083_),
    .B(_5017_),
    .C(_5037_),
    .Y(_5341_)
);

AOI21X1 _15369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4870_),
    .B(_4866_),
    .C(_4853_),
    .Y(_4882_)
);

AND2X2 _20182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9811_),
    .B(_9858_),
    .Y(_10158_)
);

FILL SFILL18760x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33560x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6371_),
    .B(_6372_),
    .Y(_6373_)
);

AOI21X1 _16310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5566_),
    .B(_5562_),
    .C(_5555_),
    .Y(_5913_)
);

NAND2X1 _21387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11474_),
    .B(_11478_),
    .Y(_11479_)
);

NAND3X1 _17935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7679_),
    .B(_7671_),
    .C(_7683_),
    .Y(_7694_)
);

INVX2 _17515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7232_),
    .Y(_7233_)
);

OAI21X1 _12650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf3),
    .B(_4116__bF$buf1),
    .C(_10463_),
    .Y(_10474_)
);

NAND3X1 _12230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4796_),
    .B(_4851_),
    .C(_4829_),
    .Y(_5870_)
);

FILL SFILL23960x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2952_),
    .C(_3224_),
    .Y(_3225_)
);

NOR2X1 _13435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_2763_),
    .Y(_2764_)
);

DFFPOSX1 _23953_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[7]),
    .CLK(clk_bF$buf7),
    .D(_0_[7])
);

AOI21X1 _13015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2298_),
    .C(_2217_),
    .Y(_2310_)
);

INVX2 _23533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1912_),
    .Y(_1917_)
);

NAND2X1 _23113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1457_),
    .B(_1458_),
    .Y(_1459_)
);

NAND2X1 _18893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_26_bF$buf3),
    .Y(_8745_)
);

INVX2 _18473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8284_),
    .Y(_8285_)
);

NAND2X1 _18053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7818_),
    .B(_7823_),
    .Y(_7824_)
);

FILL SFILL13960x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69320x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9992_),
    .B(_10336_),
    .Y(_10679_)
);

AND2X2 _20238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_28_bF$buf1),
    .Y(_10218_)
);

FILL SFILL69240x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2464_),
    .Y(_2486_)
);

NAND3X1 _19678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9276_),
    .B(_9602_),
    .C(_9603_),
    .Y(_9606_)
);

INVX1 _19258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9144_),
    .Y(_9145_)
);

AND2X2 _14393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_15_bF$buf1),
    .Y(_3813_)
);

DFFPOSX1 _24071_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[29]),
    .CLK(clk_bF$buf8),
    .D(b[29])
);

NAND3X1 _12706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10957_),
    .B(_10891_),
    .C(_10935_),
    .Y(_11088_)
);

NAND2X1 _22804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1121_),
    .B(_1116_),
    .Y(_1122_)
);

OAI21X1 _15598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5126_),
    .B(_5127_),
    .C(_5109_),
    .Y(_5132_)
);

NAND2X1 _15178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4433_),
    .B(_4600_),
    .Y(_4672_)
);

FILL SFILL3800x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59320x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11131_),
    .Y(_11270_)
);

OAI21X1 _17744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7145_),
    .B(_7484_),
    .C(_7135_),
    .Y(_7485_)
);

OAI21X1 _17324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6620_),
    .B(_6611_),
    .C(_6614_),
    .Y(_7024_)
);

NAND3X1 _18949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8761_),
    .B(_8750_),
    .C(_8754_),
    .Y(_8806_)
);

NAND2X1 _18529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_29_bF$buf0),
    .Y(_8346_)
);

XOR2X1 _18109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7838_),
    .B(_7884_),
    .Y(_7885_)
);

FILL FILL74200x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3012_),
    .B(_3014_),
    .Y(_3015_)
);

AOI21X1 _13244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2501_),
    .B(_2505_),
    .C(_2377_),
    .Y(_2555_)
);

NOR2X1 _23762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2162_),
    .B(_2164_),
    .Y(_2165_)
);

NAND2X1 _23342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_1619_),
    .Y(_1709_)
);

NAND3X1 _14869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .B(_4332_),
    .C(_4333_),
    .Y(_4334_)
);

OAI21X1 _14449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3616_),
    .B(_3601_),
    .C(_3608_),
    .Y(_3874_)
);

OAI21X1 _14029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_3402__bF$buf1),
    .C(_3399_),
    .Y(_3414_)
);

OAI21X1 _15810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5363_),
    .B(_5362_),
    .C(_5361_),
    .Y(_5364_)
);

NAND2X1 _18282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7768_),
    .B(_7774_),
    .Y(_8075_)
);

OAI21X1 _20887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10929_),
    .B(_10930_),
    .C(_10928_),
    .Y(_10931_)
);

NAND2X1 _20467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf2),
    .B(breg_20_bF$buf1),
    .Y(_10470_)
);

AND2X2 _20047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf0),
    .B(breg_28_bF$buf2),
    .Y(_10009_)
);

AND2X2 _19487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9333_),
    .B(_9394_),
    .Y(_9396_)
);

NAND2X1 _19067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8545_),
    .B(_8552_),
    .Y(_8935_)
);

FILL SFILL23960x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .B(_1642_),
    .C(_1674_),
    .Y(_1685_)
);

NOR2X1 _12515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7591_),
    .B(_8983_),
    .Y(_8994_)
);

NAND3X1 _22613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_912_),
    .B(_913_),
    .C(_910_),
    .Y(_914_)
);

FILL SFILL69000x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _23818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .B(_2223_),
    .Y(_2225_)
);

FILL SFILL74280x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert320 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5315__bF$buf1)
);

BUFX2 BUFX2_insert321 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5315__bF$buf0)
);

BUFX2 BUFX2_insert322 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .Y(_2669__bF$buf3)
);

BUFX2 BUFX2_insert323 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .Y(_2669__bF$buf2)
);

AOI21X1 _17973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7368_),
    .B(_7369_),
    .C(_7352_),
    .Y(_7736_)
);

BUFX2 BUFX2_insert324 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .Y(_2669__bF$buf1)
);

OAI21X1 _17553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6861_),
    .B(_6851_),
    .C(_6855_),
    .Y(_7275_)
);

BUFX2 BUFX2_insert325 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .Y(_2669__bF$buf0)
);

FILL SFILL13960x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert326 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf5)
);

INVX8 _17133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[30]),
    .Y(_6815_)
);

BUFX2 BUFX2_insert327 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf4)
);

BUFX2 BUFX2_insert328 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf3)
);

BUFX2 BUFX2_insert329 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf2)
);

OAI21X1 _18758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8589_),
    .B(_8590_),
    .C(_8586_),
    .Y(_8596_)
);

OAI21X1 _18338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf0),
    .B(_3781__bF$buf2),
    .C(_7721_),
    .Y(_8136_)
);

NAND2X1 _13893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_16_bF$buf1),
    .Y(_3266_)
);

NOR2X1 _13473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf2),
    .B(_8555_),
    .Y(_2806_)
);

DFFPOSX1 _23991_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[45]),
    .CLK(clk_bF$buf8),
    .D(_0_[45])
);

AOI21X1 _23571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2746_),
    .B(_2747_),
    .C(_2745_),
    .Y(_1958_)
);

OAI21X1 _13053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2347_),
    .B(_11494_),
    .C(_2346_),
    .Y(_2348_)
);

XNOR2X1 _23151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1499_),
    .B(_1495_),
    .Y(_1501_)
);

AOI21X1 _14678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_4108_),
    .C(_4112_),
    .Y(_4124_)
);

OAI21X1 _14258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3663_),
    .B(_3664_),
    .C(_3662_),
    .Y(_3665_)
);

FILL SFILL64200x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7478_),
    .B(_7476_),
    .C(_7479_),
    .Y(_7866_)
);

OAI21X1 _20696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf0),
    .B(_5668__bF$buf5),
    .C(_10708_),
    .Y(_10721_)
);

NOR2X1 _20276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10260_),
    .B(_10256_),
    .Y(_10261_)
);

AOI21X1 _16824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_6465_),
    .C(_6443_),
    .Y(_6476_)
);

NAND3X1 _16404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5666_),
    .B(_6010_),
    .C(_6015_),
    .Y(_6016_)
);

NAND3X1 _19296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9176_),
    .B(_9183_),
    .C(_9186_),
    .Y(_9187_)
);

NAND2X1 _17609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6894_),
    .B(_6902_),
    .Y(_7336_)
);

OAI21X1 _12744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11472_),
    .B(_11461_),
    .C(_9981_),
    .Y(_11505_)
);

OAI21X1 _12324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .B(_6878_),
    .C(_6845_),
    .Y(_6900_)
);

NOR2X1 _22842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1154_),
    .Y(_1164_)
);

NAND3X1 _22422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_699_),
    .C(_698_),
    .Y(_705_)
);

INVX2 _22002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .Y(_244_)
);

NAND2X1 _13949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3325_),
    .B(_3326_),
    .Y(_3327_)
);

OAI21X1 _13529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2865_),
    .B(_2866_),
    .C(_2864_),
    .Y(_2867_)
);

NOR2X1 _13109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(_1968_),
    .Y(_2407_)
);

NOR2X1 _23627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2007_),
    .B(_2018_),
    .Y(_2019_)
);

OAI21X1 _23207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1417_),
    .C(_1422_),
    .Y(_1561_)
);

FILL SFILL3720x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7522_),
    .B(_7526_),
    .Y(_7527_)
);

NAND2X1 _17362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_22_bF$buf4),
    .Y(_7067_)
);

FILL SFILL34120x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8415_),
    .B(_8421_),
    .C(_8425_),
    .Y(_8847_)
);

NAND2X1 _18567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8385_),
    .B(_8386_),
    .Y(_8387_)
);

AOI21X1 _18147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7551_),
    .B(_7546_),
    .C(_7513_),
    .Y(_7927_)
);

NAND2X1 _13282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_10_bF$buf3),
    .Y(_2596_)
);

NOR3X1 _23380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .B(_1737_),
    .C(_1741_),
    .Y(_1750_)
);

FILL SFILL8680x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_14_bF$buf0),
    .Y(_3916_)
);

AOI21X1 _14067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3442_),
    .B(_3435_),
    .C(_3357_),
    .Y(_3456_)
);

FILL SFILL8600x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10050_),
    .B(_10049_),
    .C(_10045_),
    .Y(_10051_)
);

OAI21X1 _16633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5887_),
    .B(_6266_),
    .C(_5896_),
    .Y(_6267_)
);

NOR3X1 _16213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5800_),
    .B(_5802_),
    .C(_5799_),
    .Y(_5807_)
);

FILL SFILL74200x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7586_),
    .B(_7587_),
    .C(_7585_),
    .Y(_7588_)
);

OAI21X1 _17418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7127_),
    .B(_7126_),
    .C(_7121_),
    .Y(_7128_)
);

NAND2X1 _12973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2055_),
    .B(_1968_),
    .Y(_2099_)
);

NAND3X1 _12553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9389_),
    .B(_9400_),
    .C(_9378_),
    .Y(_9411_)
);

NOR3X1 _12133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4774_),
    .B(_4763_),
    .C(_4730_),
    .Y(_4807_)
);

NAND2X1 _22651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_762_),
    .Y(_955_)
);

INVX2 _22231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .Y(_495_)
);

OAI21X1 _13758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_2287__bF$buf2),
    .C(_2872_),
    .Y(_3118_)
);

NOR2X1 _13338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2656_),
    .B(_2657_),
    .Y(_2658_)
);

NAND2X1 _23856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2264_),
    .Y(_2265_)
);

NAND2X1 _23436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .B(areg_30_bF$buf4),
    .Y(_1811_)
);

NOR2X1 _23016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1352_),
    .Y(_1353_)
);

FILL SFILL33800x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .B(_6887_),
    .C(_7315_),
    .Y(_7317_)
);

NAND2X1 _17171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_24_bF$buf4),
    .Y(_6857_)
);

NAND2X1 _15904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_14_bF$buf1),
    .Y(_5468_)
);

AOI21X1 _18796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7823_),
    .B(_8637_),
    .C(_8241_),
    .Y(_8638_)
);

OAI21X1 _18376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8176_),
    .B(_8175_),
    .C(_8177_),
    .Y(_8178_)
);

NAND2X1 _13091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_9_bF$buf2),
    .Y(_2388_)
);

NAND3X1 _21922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_152_),
    .C(_151_),
    .Y(_157_)
);

NOR2X1 _21502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf2),
    .B(_7225__bF$buf4),
    .Y(_11605_)
);

AOI21X1 _14296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3706_),
    .B(_3700_),
    .C(_3666_),
    .Y(_3707_)
);

FILL SFILL39000x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10013_),
    .B(_9488_),
    .C(_9422_),
    .Y(_10024_)
);

OAI21X1 _22707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1015_),
    .C(_1011_),
    .Y(_1016_)
);

OAI21X1 _16862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .B(_6138_),
    .C(_6147_),
    .Y(_6518_)
);

OAI21X1 _16442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5713_),
    .B(_6056_),
    .C(_5707_),
    .Y(_6057_)
);

OAI21X1 _16022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5595_),
    .B(_5597_),
    .C(_5594_),
    .Y(_5598_)
);

NAND3X1 _21099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11153_),
    .B(_11152_),
    .C(_11158_),
    .Y(_11163_)
);

NOR2X1 _17647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7372_),
    .B(_7377_),
    .Y(_7378_)
);

NAND3X1 _17227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6915_),
    .B(_6916_),
    .C(_6917_),
    .Y(_6918_)
);

FILL SFILL23640x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10496_),
    .B(_10540_),
    .C(_10562_),
    .Y(_12_)
);

NOR2X1 _12362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7305_),
    .B(_6253_),
    .Y(_7316_)
);

OR2X2 _22880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1204_),
    .Y(_1205_)
);

NOR2X1 _22460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf2),
    .B(_6427_),
    .Y(_745_)
);

AOI21X1 _22040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_281_),
    .C(_255_),
    .Y(_285_)
);

FILL SFILL8680x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3363_),
    .B(_3367_),
    .C(_3366_),
    .Y(_3368_)
);

OAI21X1 _13567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2908_),
    .B(_2900_),
    .C(_2868_),
    .Y(_2909_)
);

NOR2X1 _13147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf2),
    .B(_7711__bF$buf1),
    .Y(_2449_)
);

NAND2X1 _23665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2059_),
    .B(_2044_),
    .Y(_2060_)
);

NAND2X1 _23245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1573_),
    .B(_1602_),
    .Y(_1603_)
);

FILL SFILL48840x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5246_),
    .B(_5247_),
    .C(_5103_),
    .Y(_5259_)
);

FILL SFILL34120x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _18185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf5),
    .B(areg_31_bF$buf1),
    .C(breg_2_bF$buf4),
    .D(areg_30_bF$buf0),
    .Y(_7969_)
);

AOI21X1 _16918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6574_),
    .B(_6575_),
    .C(_6573_),
    .Y(_6579_)
);

NAND3X1 _21731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11599_),
    .B(_11852_),
    .C(_11851_),
    .Y(_11856_)
);

NAND3X1 _21311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11391_),
    .B(_11378_),
    .C(_11382_),
    .Y(_11396_)
);

FILL SFILL64280x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .Y(_626_)
);

NAND3X1 _12418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7876_),
    .B(_7920_),
    .C(_7547_),
    .Y(_7931_)
);

NAND2X1 _22936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1179_),
    .B(_1183_),
    .Y(_1266_)
);

NOR3X1 _22516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_625_),
    .B(_618_),
    .C(_629_),
    .Y(_807_)
);

FILL SFILL64200x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf0),
    .B(areg_26_bF$buf0),
    .Y(_6309_)
);

INVX2 _16251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5847_),
    .Y(_5849_)
);

OAI21X1 _17876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7626_),
    .B(_7627_),
    .C(_7220_),
    .Y(_7630_)
);

NAND3X1 _17456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7163_),
    .B(_7169_),
    .C(_7013_),
    .Y(_7170_)
);

AOI21X1 _17036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6310_),
    .B(_6315_),
    .C(_6320_),
    .Y(_6709_)
);

NAND3X1 _12591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8467_),
    .B(_9817_),
    .C(_9762_),
    .Y(_9828_)
);

OAI21X1 _12171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_3646__bF$buf1),
    .C(_5212_),
    .Y(_5233_)
);

FILL SFILL43960x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3152_),
    .B(_3159_),
    .Y(_3160_)
);

AOI21X1 _13376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2696_),
    .B(_2695_),
    .C(_2693_),
    .Y(_2700_)
);

BUFX2 _23894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[12]),
    .Y(y[12])
);

NOR3X1 _23474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1727_),
    .C(_1844_),
    .Y(_1853_)
);

NAND3X1 _23054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1264_),
    .B(_1386_),
    .C(_1379_),
    .Y(_1395_)
);

NAND3X1 _19602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9483_),
    .B(_9517_),
    .C(_9522_),
    .Y(_9523_)
);

NAND3X1 _15942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5509_),
    .B(_5507_),
    .C(_5506_),
    .Y(_5510_)
);

NAND2X1 _15522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5046_),
    .B(_5048_),
    .Y(_5049_)
);

NAND3X1 _15102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4570_),
    .B(_4576_),
    .C(_4580_),
    .Y(_4590_)
);

AOI21X1 _20599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10602_),
    .B(_10607_),
    .C(_10614_),
    .Y(_10615_)
);

OAI21X1 _20179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_4541__bF$buf0),
    .C(_10148_),
    .Y(_10154_)
);

NAND3X1 _16727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6364_),
    .B(_6369_),
    .C(_6217_),
    .Y(_6370_)
);

NAND3X1 _16307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5896_),
    .B(_5899_),
    .C(_5900_),
    .Y(_5910_)
);

AOI21X1 _21960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11836_),
    .B(_11835_),
    .C(_11830_),
    .Y(_198_)
);

AND2X2 _21540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11642_),
    .B(_11645_),
    .Y(_11646_)
);

AOI21X1 _21120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11175_),
    .B(_11174_),
    .C(_11171_),
    .Y(_11186_)
);

NAND3X1 _19199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9040_),
    .B(_9073_),
    .C(_9076_),
    .Y(_9080_)
);

FILL SFILL13720x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8742_),
    .B(_8775_),
    .C(_8808_),
    .Y(_10441_)
);

NOR3X1 _12227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4204_),
    .B(_5705_),
    .C(_5749_),
    .Y(_5837_)
);

XNOR2X1 _22745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .B(_1057_),
    .Y(_1058_)
);

NAND3X1 _22325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_597_),
    .C(_592_),
    .Y(_598_)
);

FILL SFILL48840x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _16480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6091_),
    .B(_6092_),
    .C(_6094_),
    .Y(_6098_)
);

AOI21X1 _16060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5621_),
    .B(_5625_),
    .C(_5366_),
    .Y(_5639_)
);

FILL SFILL34120x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7044_),
    .B(_7049_),
    .C(_7050_),
    .Y(_7420_)
);

NAND2X1 _17265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6554_),
    .B(_6556_),
    .Y(_6960_)
);

AOI21X1 _20811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10846_),
    .B(_10845_),
    .C(_10844_),
    .Y(_10848_)
);

NOR2X1 _13185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .B(_2490_),
    .Y(_2491_)
);

OAI21X1 _23283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1644_),
    .B(_1640_),
    .C(_1548_),
    .Y(_1645_)
);

NAND2X1 _19831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf2),
    .B(areg_19_bF$buf4),
    .Y(_9774_)
);

OAI21X1 _19411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9311_),
    .B(_9307_),
    .C(_9280_),
    .Y(_9313_)
);

NAND2X1 _11918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_3_bF$buf4),
    .Y(_2453_)
);

FILL SFILL3480x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24068_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[26]),
    .CLK(clk_bF$buf5),
    .D(b[26])
);

INVX1 _15751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5298_),
    .Y(_5300_)
);

NAND3X1 _15331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4834_),
    .B(_4839_),
    .C(_4817_),
    .Y(_4841_)
);

OAI21X1 _16956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6620_),
    .B(_6619_),
    .C(_6611_),
    .Y(_6621_)
);

AOI21X1 _16536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6158_),
    .B(_6159_),
    .C(_6157_),
    .Y(_6160_)
);

NAND3X1 _16116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5675_),
    .B(_5699_),
    .C(_5690_),
    .Y(_5700_)
);

NAND3X1 _12876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11668_),
    .B(_1031_),
    .C(_965_),
    .Y(_1042_)
);

OAI21X1 _12456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8315_),
    .B(_8326_),
    .C(_8337_),
    .Y(_8348_)
);

NAND3X1 _22974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1304_),
    .B(_1300_),
    .C(_1306_),
    .Y(_1307_)
);

NAND2X1 _12036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3591_),
    .B(_3679_),
    .Y(_3745_)
);

NOR2X1 _22554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_627_),
    .Y(_849_)
);

NAND3X1 _22134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_380_),
    .C(_384_),
    .Y(_389_)
);

NOR2X1 _23759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2161_),
    .B(_2160_),
    .Y(_0_[58])
);

AND2X2 _23339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1578_),
    .B(_1703_),
    .Y(_1705_)
);

NAND3X1 _14602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .B(_4039_),
    .C(_3775_),
    .Y(_4042_)
);

NAND3X1 _17494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7197_),
    .B(_7201_),
    .C(_7204_),
    .Y(_7211_)
);

NOR3X1 _17074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6353_),
    .B(_6354_),
    .C(_6351_),
    .Y(_6751_)
);

INVX1 _15807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4996_),
    .Y(_5361_)
);

OAI21X1 _20620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10622_),
    .B(_10629_),
    .C(_10632_),
    .Y(_10638_)
);

AOI21X1 _20200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10175_),
    .B(_10176_),
    .C(_10169_),
    .Y(_10177_)
);

NAND2X1 _18699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_25_bF$buf5),
    .Y(_8531_)
);

OAI21X1 _18279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7696_),
    .B(_7666_),
    .C(_7704_),
    .Y(_8071_)
);

AND2X2 _23092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1431_),
    .B(_1435_),
    .Y(_1436_)
);

NAND3X1 _19640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9556_),
    .B(_9557_),
    .C(_9560_),
    .Y(_9564_)
);

XNOR2X1 _19220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9101_),
    .B(_9099_),
    .Y(_9102_)
);

FILL SFILL69080x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_28_),
    .Y(_50_)
);

OAI21X1 _21405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11490_),
    .B(_11491_),
    .C(_11488_),
    .Y(_11499_)
);

INVX1 _14199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3599_),
    .Y(_3600_)
);

AND2X2 _15980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .B(_5546_),
    .Y(_5551_)
);

AOI21X1 _15560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5088_),
    .B(_5079_),
    .C(_5089_),
    .Y(_5090_)
);

AOI21X1 _15140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4058_),
    .B(_4326_),
    .C(_4630_),
    .Y(_4631_)
);

NAND3X1 _16765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6404_),
    .B(_6411_),
    .C(_6030_),
    .Y(_6412_)
);

NAND3X1 _16345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5940_),
    .B(_5942_),
    .C(_5937_),
    .Y(_5952_)
);

FILL SFILL3560x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert290 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf4)
);

BUFX2 BUFX2_insert291 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf3)
);

BUFX2 BUFX2_insert292 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf2)
);

BUFX2 BUFX2_insert293 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf1)
);

BUFX2 BUFX2_insert294 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf0)
);

BUFX2 BUFX2_insert295 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[21]),
    .Y(breg_21_bF$buf4)
);

BUFX2 BUFX2_insert296 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[21]),
    .Y(breg_21_bF$buf3)
);

FILL SFILL69240x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert297 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[21]),
    .Y(breg_21_bF$buf2)
);

BUFX2 BUFX2_insert298 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[21]),
    .Y(breg_21_bF$buf1)
);

FILL SFILL43960x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10836_),
    .B(_10847_),
    .Y(_10858_)
);

BUFX2 BUFX2_insert299 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[21]),
    .Y(breg_21_bF$buf0)
);

AND2X2 _12265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6231_),
    .B(_6132_),
    .Y(_6253_)
);

OAI21X1 _22783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_953_),
    .C(_975_),
    .Y(_1099_)
);

AOI21X1 _22363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_639_),
    .C(_636_),
    .Y(_640_)
);

FILL SFILL28920x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _18911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8339_),
    .Y(_8765_)
);

FILL SFILL73960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23988_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[42]),
    .CLK(clk_bF$buf7),
    .D(_0_[42])
);

INVX1 _23568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7647_),
    .Y(_1954_)
);

NOR2X1 _23148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1348_),
    .B(_1496_),
    .Y(_1497_)
);

NAND3X1 _14831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4273_),
    .B(_4279_),
    .C(_4283_),
    .Y(_4293_)
);

NAND3X1 _14411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .B(_3831_),
    .C(_3825_),
    .Y(_3833_)
);

OAI21X1 _15616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4815_),
    .B(_5151_),
    .C(_4824_),
    .Y(_5152_)
);

NAND3X1 _18088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7817_),
    .B(_7850_),
    .C(_7853_),
    .Y(_7862_)
);

XNOR2X1 _11956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2858_),
    .B(_2781_),
    .Y(_2869_)
);

OAI21X1 _21634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11735_),
    .B(_11739_),
    .C(_11741_),
    .Y(_11749_)
);

OAI21X1 _21214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11285_),
    .B(_11289_),
    .C(_11009_),
    .Y(_11290_)
);

NAND3X1 _22839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .B(_1159_),
    .C(_1155_),
    .Y(_1160_)
);

OAI21X1 _22419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_697_),
    .B(_700_),
    .C(_492_),
    .Y(_701_)
);

OAI21X1 _16994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_4541__bF$buf3),
    .C(_6654_),
    .Y(_6663_)
);

OAI21X1 _16574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6196_),
    .B(_6197_),
    .C(_6162_),
    .Y(_6202_)
);

NAND3X1 _16154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5739_),
    .B(_5740_),
    .C(_5741_),
    .Y(_5742_)
);

NOR2X1 _17779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7517_),
    .B(_7518_),
    .Y(_7523_)
);

AOI21X1 _17359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6720_),
    .B(_6716_),
    .C(_6679_),
    .Y(_7063_)
);

NOR2X1 _12494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7338_),
    .B(_8753_),
    .Y(_8764_)
);

NAND2X1 _12074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf4),
    .B(breg_4_bF$buf5),
    .Y(_4160_)
);

NAND3X1 _22592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_885_),
    .C(_890_),
    .Y(_891_)
);

NOR3X1 _22172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_401_),
    .B(_416_),
    .C(_421_),
    .Y(_431_)
);

NAND3X1 _18720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8550_),
    .B(_8536_),
    .C(_8540_),
    .Y(_8554_)
);

NAND2X1 _18300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg_28_bF$buf0),
    .Y(_8094_)
);

XNOR2X1 _20905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10605_),
    .B(_10950_),
    .Y(_10951_)
);

NAND2X1 _13699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_12_bF$buf3),
    .Y(_3053_)
);

AOI21X1 _13279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2394_),
    .C(_2592_),
    .Y(_2593_)
);

INVX1 _23797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2202_),
    .Y(_2203_)
);

AOI21X1 _23377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1742_),
    .B(_1746_),
    .C(_1623_),
    .Y(_1747_)
);

AOI21X1 _19925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9491_),
    .B(_9495_),
    .C(_9498_),
    .Y(_9877_)
);

AOI21X1 _19505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9406_),
    .B(_9405_),
    .C(_9402_),
    .Y(_9416_)
);

INVX2 _14640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4075_),
    .Y(_4082_)
);

OAI21X1 _14220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(_3610_),
    .C(_3599_),
    .Y(_3623_)
);

FILL SFILL3640x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5401_),
    .B(_5402_),
    .C(_5400_),
    .Y(_5403_)
);

NAND3X1 _15425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4654_),
    .B(_4937_),
    .C(_4943_),
    .Y(_4944_)
);

OAI21X1 _15005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4206_),
    .B(_4231_),
    .C(_4222_),
    .Y(_4483_)
);

NAND3X1 _21863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_88_),
    .C(_90_),
    .Y(_92_)
);

NAND3X1 _21443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11522_),
    .B(_11540_),
    .C(_11518_),
    .Y(_11541_)
);

OAI21X1 _21023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf2),
    .B(_3781__bF$buf3),
    .C(_10755_),
    .Y(_11080_)
);

FILL SFILL33880x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _22648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .Y(_951_)
);

AOI21X1 _22228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(_470_),
    .C(_246_),
    .Y(_491_)
);

FILL SFILL49080x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3259_),
    .B(_3279_),
    .C(_3284_),
    .Y(_3286_)
);

OAI21X1 _16383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5985_),
    .B(_5986_),
    .C(_5838_),
    .Y(_5993_)
);

NAND3X1 _17588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7310_),
    .B(_7312_),
    .C(_7311_),
    .Y(_7313_)
);

FILL SFILL18840x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_25_bF$buf4),
    .Y(_6853_)
);

FILL SFILL39000x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10431_),
    .B(_10433_),
    .C(_10424_),
    .Y(_10741_)
);

NOR2X1 _13088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .B(_2382_),
    .Y(_2384_)
);

INVX1 _23186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1254_),
    .Y(_1538_)
);

OAI21X1 _19734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_9656_),
    .Y(_9667_)
);

NAND3X1 _19314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9084_),
    .B(_9088_),
    .C(_9090_),
    .Y(_9207_)
);

FILL SFILL29080x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_151_),
    .C(_128_),
    .Y(_153_)
);

FILL SFILL8760x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4855_),
    .B(_4859_),
    .C(_4858_),
    .Y(_5194_)
);

NAND3X1 _15234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4711_),
    .B(_4726_),
    .C(_4733_),
    .Y(_4734_)
);

FILL SFILL53960x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_21_bF$buf0),
    .Y(_6514_)
);

OAI21X1 _16439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5726_),
    .B(_6049_),
    .C(_6052_),
    .Y(_6053_)
);

AOI21X1 _16019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5178_),
    .B(_5222_),
    .C(_5593_),
    .Y(_5594_)
);

XNOR2X1 _11994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3176_),
    .B(_2387_),
    .Y(_3285_)
);

AOI21X1 _21672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11790_),
    .B(_11788_),
    .C(_11781_),
    .Y(_11791_)
);

NOR2X1 _21252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf2),
    .B(_6815__bF$buf0),
    .Y(_11331_)
);

NAND3X1 _17800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7541_),
    .B(_7545_),
    .C(_7527_),
    .Y(_7546_)
);

OAI21X1 _12779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10123_),
    .B(_10233_),
    .C(_11844_),
    .Y(_11887_)
);

INVX2 _12359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7272_),
    .Y(_7283_)
);

AOI21X1 _22877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1200_),
    .B(_1046_),
    .C(_1201_),
    .Y(_1202_)
);

NAND2X1 _22457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_28_bF$buf3),
    .Y(_742_)
);

FILL SFILL3720x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_280_),
    .C(_281_),
    .Y(_282_)
);

FILL SFILL43960x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3075_),
    .B(_3074_),
    .C(_3059_),
    .Y(_3076_)
);

AND2X2 _13300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2433_),
    .Y(_2615_)
);

NAND2X1 _16192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_17_bF$buf3),
    .Y(_5783_)
);

FILL SFILL43880x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_15_bF$buf5),
    .Y(_4395_)
);

AOI21X1 _14505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3923_),
    .B(_3922_),
    .C(_3918_),
    .Y(_3936_)
);

OAI21X1 _17397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7104_),
    .B(_7103_),
    .C(_7094_),
    .Y(_7105_)
);

OAI22X1 _20943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10988_),
    .B(_10992_),
    .C(_10649_),
    .D(_10689_),
    .Y(_10993_)
);

AOI21X1 _20523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10530_),
    .B(_10531_),
    .C(_10523_),
    .Y(_10532_)
);

OAI21X1 _20103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9786_),
    .B(_9788_),
    .C(_9778_),
    .Y(_10071_)
);

NAND3X1 _19963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9897_),
    .B(_9891_),
    .C(_9895_),
    .Y(_9918_)
);

NAND3X1 _19543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9451_),
    .B(_9452_),
    .C(_9453_),
    .Y(_9458_)
);

NAND3X1 _19123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8891_),
    .B(_8991_),
    .C(_8996_),
    .Y(_8997_)
);

FILL SFILL33880x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11601_),
    .B(_11843_),
    .C(_11839_),
    .Y(_11852_)
);

OAI21X1 _21308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11388_),
    .B(_11389_),
    .C(_11391_),
    .Y(_11392_)
);

NAND2X1 _15883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5399_),
    .B(_5403_),
    .Y(_5445_)
);

OAI21X1 _15463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4983_),
    .B(_4704_),
    .C(_4698_),
    .Y(_4984_)
);

OAI21X1 _15043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4523_),
    .B(_4524_),
    .C(_4499_),
    .Y(_4525_)
);

FILL SFILL18600x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6304_),
    .B(_6303_),
    .C(_6294_),
    .Y(_6305_)
);

XNOR2X1 _16248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5844_),
    .B(_5841_),
    .Y(_5845_)
);

AOI21X1 _21481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11581_),
    .B(_11580_),
    .C(_11319_),
    .Y(_11583_)
);

FILL SFILL23880x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10898_),
    .B(_10901_),
    .C(_10899_),
    .Y(_11122_)
);

FILL SFILL54280x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9718_),
    .B(_9641_),
    .C(_9696_),
    .Y(_9795_)
);

INVX8 _12168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .Y(_5190_)
);

OAI21X1 _22686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_841_),
    .C(_847_),
    .Y(_993_)
);

FILL SFILL23800x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _22266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_507_),
    .B(_520_),
    .C(_524_),
    .Y(_533_)
);

AND2X2 _18814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8243_),
    .B(_8286_),
    .Y(_8658_)
);

FILL SFILL8840x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4176_),
    .B(_4170_),
    .C(_4174_),
    .Y(_4186_)
);

AOI21X1 _14314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3725_),
    .B(_3726_),
    .C(_3724_),
    .Y(_3727_)
);

FILL SFILL49000x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5129_),
    .B(_5121_),
    .Y(_5506_)
);

INVX1 _15519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5044_),
    .Y(_5045_)
);

NOR3X1 _20752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10775_),
    .B(_10776_),
    .C(_10778_),
    .Y(_10783_)
);

AOI21X1 _20332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10317_),
    .B(_10322_),
    .C(_9992_),
    .Y(_10323_)
);

AOI21X1 _19772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9392_),
    .B(_9708_),
    .C(_9395_),
    .Y(_9709_)
);

OAI21X1 _19352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .B(_9248_),
    .C(_8881_),
    .Y(_9249_)
);

NAND3X1 _21957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_11826_),
    .C(_185_),
    .Y(_195_)
);

FILL SFILL3720x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11640_),
    .B(_11639_),
    .C(_11638_),
    .Y(_11643_)
);

OAI22X1 _21117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10558_),
    .B(_11181_),
    .C(_11182_),
    .D(_10911_),
    .Y(_11183_)
);

FILL SFILL43960x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_166_),
    .Y(_210_)
);

NAND3X1 _15692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5228_),
    .B(_5234_),
    .C(_5148_),
    .Y(_5235_)
);

NAND2X1 _15272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf4),
    .B(areg_13_bF$buf2),
    .Y(_4776_)
);

NAND3X1 _16897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6551_),
    .B(_6555_),
    .C(_6554_),
    .Y(_6556_)
);

OAI21X1 _16477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6091_),
    .B(_6092_),
    .C(_6094_),
    .Y(_6095_)
);

OAI21X1 _16057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5623_),
    .B(_5624_),
    .C(_5367_),
    .Y(_5636_)
);

NAND2X1 _21290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_26_bF$buf4),
    .Y(_11372_)
);

CLKBUF1 CLKBUF1_insert84 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert85 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert86 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert87 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert88 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert89 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

OR2X2 _12397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_7689_),
    .Y(_7700_)
);

OR2X2 _22495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_553_),
    .B(_783_),
    .Y(_784_)
);

NAND3X1 _22075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_322_),
    .C(_323_),
    .Y(_324_)
);

AOI21X1 _18623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7660_),
    .B(_8043_),
    .C(_8049_),
    .Y(_8449_)
);

OAI21X1 _18203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7978_),
    .C(_7981_),
    .Y(_7989_)
);

XNOR2X1 _20808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10819_),
    .B(_10816_),
    .Y(_10844_)
);

NAND2X1 _19828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9768_),
    .B(_9769_),
    .Y(_9770_)
);

AOI21X1 _19408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9305_),
    .B(_9304_),
    .C(_9282_),
    .Y(_9309_)
);

AOI21X1 _14963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4155_),
    .B(_4197_),
    .C(_4194_),
    .Y(_4437_)
);

AOI21X1 _14543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3969_),
    .B(_3977_),
    .C(_3955_),
    .Y(_3978_)
);

NOR3X1 _14123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3484_),
    .B(_3485_),
    .C(_3483_),
    .Y(_3517_)
);

XNOR2X1 _15748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4963_),
    .B(_5296_),
    .Y(_0_[25])
);

INVX1 _15328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4532_),
    .Y(_4837_)
);

OAI21X1 _20981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11032_),
    .B(_11031_),
    .C(_11023_),
    .Y(_11033_)
);

FILL SFILL23880x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10569_),
    .B(_10572_),
    .C(_10561_),
    .Y(_10574_)
);

INVX2 _20141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10111_),
    .Y(_10113_)
);

NOR2X1 _19581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9492_),
    .B(_9493_),
    .Y(_9500_)
);

NAND2X1 _19161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9033_),
    .B(_9037_),
    .Y(_9039_)
);

NOR2X1 _21766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf1),
    .B(_6815__bF$buf0),
    .Y(_11893_)
);

AND2X2 _21346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11111_),
    .B(_11103_),
    .Y(_11434_)
);

FILL SFILL8840x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4560_),
    .B(_4561_),
    .C(_4559_),
    .Y(_4567_)
);

FILL SFILL74520x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3164_),
    .B(_3169_),
    .C(_3171_),
    .Y(_3180_)
);

BUFX2 _23912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[30]),
    .Y(y[30])
);

NAND2X1 _16286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_20_bF$buf1),
    .Y(_5887_)
);

FILL SFILL13800x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _18852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8657_),
    .B(_8699_),
    .Y(_8700_)
);

NAND3X1 _18432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8239_),
    .B(_8232_),
    .C(_8235_),
    .Y(_8240_)
);

NAND3X1 _18012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7776_),
    .B(_7778_),
    .C(_7775_),
    .Y(_7779_)
);

NAND3X1 _20617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10633_),
    .B(_10634_),
    .C(_10632_),
    .Y(_10635_)
);

FILL SFILL19000x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1428_),
    .B(_1429_),
    .Y(_1432_)
);

AOI21X1 _19637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9557_),
    .B(_9560_),
    .C(_9556_),
    .Y(_9561_)
);

INVX2 _19217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9098_),
    .Y(_9099_)
);

OAI21X1 _14772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4223_),
    .B(_4224_),
    .C(_4227_),
    .Y(_4228_)
);

AOI21X1 _14352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3764_),
    .C(_3517_),
    .Y(_3768_)
);

DFFPOSX1 _24030_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[20]),
    .CLK(clk_bF$buf0),
    .D(a[20])
);

OAI21X1 _15977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_4541__bF$buf3),
    .C(_5545_),
    .Y(_5548_)
);

NAND3X1 _15557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5073_),
    .B(_5066_),
    .C(_5071_),
    .Y(_5087_)
);

NAND3X1 _15137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4349_),
    .B(_4627_),
    .C(_4626_),
    .Y(_4628_)
);

OAI21X1 _20790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253__bF$buf3),
    .B(_3961__bF$buf1),
    .C(_10823_),
    .Y(_10824_)
);

NAND3X1 _20370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10358_),
    .B(_10362_),
    .C(_10361_),
    .Y(_10363_)
);

NAND2X1 _19390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9287_),
    .B(_9288_),
    .Y(_9289_)
);

NAND2X1 _21995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_233_),
    .Y(_236_)
);

OAI21X1 _21575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11680_),
    .B(_11681_),
    .C(_11683_),
    .Y(_11684_)
);

AND2X2 _21155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10932_),
    .B(_10927_),
    .Y(_11225_)
);

NAND2X1 _17703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_19_bF$buf5),
    .Y(_7440_)
);

FILL SFILL54040x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8363_),
    .B(_8760_),
    .C(_8371_),
    .Y(_8761_)
);

NOR2X1 _13623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .B(_2736_),
    .Y(_2971_)
);

AOI21X1 _13203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2495_),
    .B(_2500_),
    .C(_2422_),
    .Y(_2511_)
);

INVX1 _23721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2100_),
    .Y(_2121_)
);

OAI21X1 _23301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_1608_),
    .C(_1605_),
    .Y(_1664_)
);

NOR2X1 _16095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_5676_),
    .Y(_5677_)
);

OAI21X1 _14828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4194_),
    .B(_4189_),
    .C(_4196_),
    .Y(_4289_)
);

AOI21X1 _14408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3827_),
    .B(_3828_),
    .C(_3826_),
    .Y(_3829_)
);

FILL SFILL54040x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8097_),
    .B(_8087_),
    .C(_8091_),
    .Y(_8490_)
);

NAND3X1 _18241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8022_),
    .B(_7782_),
    .C(_8023_),
    .Y(_8030_)
);

FILL SFILL8920x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10884_),
    .B(_10885_),
    .C(_10877_),
    .Y(_10886_)
);

AOI21X1 _20426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10420_),
    .B(_10421_),
    .C(_10418_),
    .Y(_10425_)
);

OAI21X1 _20006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9961_),
    .B(_9964_),
    .C(_9639_),
    .Y(_9965_)
);

AND2X2 _19866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9446_),
    .B(_9485_),
    .Y(_9812_)
);

AOI21X1 _19446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9341_),
    .B(_9336_),
    .C(_9321_),
    .Y(_9351_)
);

OAI21X1 _19026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8889_),
    .B(_8598_),
    .C(_8843_),
    .Y(_8890_)
);

NAND3X1 _14581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3780_),
    .B(_3863_),
    .C(_3862_),
    .Y(_4020_)
);

OAI21X1 _14161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3556_),
    .B(_3557_),
    .C(_3551_),
    .Y(_3559_)
);

FILL SFILL69160x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(_5336_),
    .C(_5337_),
    .Y(_5338_)
);

NOR3X1 _15366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4556_),
    .B(_4550_),
    .C(_4554_),
    .Y(_4879_)
);

FILL SFILL13800x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf3),
    .B(areg_25_bF$buf3),
    .Y(_11476_)
);

NOR3X1 _17932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7690_),
    .B(_7685_),
    .C(_7688_),
    .Y(_7691_)
);

NAND2X1 _17512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6833_),
    .B(_7229_),
    .Y(_7230_)
);

FILL SFILL24040x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23720x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_669_),
    .C(_886_),
    .Y(_887_)
);

NAND3X1 _22169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_399_),
    .B(_426_),
    .C(_422_),
    .Y(_427_)
);

FILL SFILL64120x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8547_),
    .B(_8546_),
    .C(_8550_),
    .Y(_8551_)
);

AOI21X1 _13852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3219_),
    .B(_3221_),
    .C(_2984_),
    .Y(_3222_)
);

INVX1 _13432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .Y(_2761_)
);

DFFPOSX1 _23950_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[4]),
    .CLK(clk_bF$buf7),
    .D(_0_[4])
);

OAI21X1 _13012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2297_),
    .C(_2249_),
    .Y(_2307_)
);

XNOR2X1 _23530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1911_),
    .B(_1897_),
    .Y(_1912_)
);

FILL SFILL28680x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _23110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(_1441_),
    .Y(_1455_)
);

NAND2X1 _14637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf4),
    .B(breg_18_bF$buf5),
    .Y(_4079_)
);

INVX1 _14217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3594_),
    .Y(_3620_)
);

OAI21X1 _18890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8360_),
    .B(_8397_),
    .C(_8388_),
    .Y(_8741_)
);

OAI21X1 _18470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7926_),
    .B(_8280_),
    .C(_8002_),
    .Y(_8281_)
);

NAND2X1 _18050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf2),
    .B(breg_17_bF$buf0),
    .Y(_7820_)
);

AOI21X1 _20655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10657_),
    .B(_10658_),
    .C(_10656_),
    .Y(_10676_)
);

OAI21X1 _20235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9874_),
    .B(_9863_),
    .C(_9867_),
    .Y(_10215_)
);

NAND3X1 _19675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9590_),
    .B(_9584_),
    .C(_9387_),
    .Y(_9603_)
);

AND2X2 _19255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_28_bF$buf5),
    .Y(_9142_)
);

OAI21X1 _14390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3548_),
    .B(_3540_),
    .C(_3543_),
    .Y(_3809_)
);

FILL SFILL19000x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33880x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11000_),
    .B(_11044_),
    .C(_10704_),
    .Y(_11055_)
);

NAND2X1 _22801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf0),
    .B(breg_27_bF$buf1),
    .Y(_1119_)
);

NAND3X1 _15595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5121_),
    .B(_5128_),
    .C(_5108_),
    .Y(_5129_)
);

NOR2X1 _15175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4668_),
    .B(_4666_),
    .Y(_4669_)
);

NOR3X1 _13908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3276_),
    .B(_3271_),
    .C(_3277_),
    .Y(_3282_)
);

FILL SFILL44040x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11118_),
    .B(_11124_),
    .C(_11126_),
    .Y(_11267_)
);

OAI21X1 _17741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7479_),
    .B(_7480_),
    .C(_7478_),
    .Y(_7482_)
);

AND2X2 _17321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6606_),
    .B(_7018_),
    .Y(_7021_)
);

NOR2X1 _22398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_673_),
    .Y(_677_)
);

NOR3X1 _18946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8384_),
    .B(_8390_),
    .C(_8394_),
    .Y(_8803_)
);

OAI21X1 _18526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf2),
    .B(_6686__bF$buf3),
    .C(_8339_),
    .Y(_8343_)
);

NAND2X1 _18106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf3),
    .B(areg_18_bF$buf0),
    .Y(_7882_)
);

NOR2X1 _13661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2765_),
    .Y(_3012_)
);

OAI21X1 _13241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2550_),
    .B(_2359_),
    .C(_2517_),
    .Y(_2552_)
);

FILL SFILL38760x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4327_),
    .B(_4056_),
    .C(_4330_),
    .Y(_4331_)
);

FILL SFILL74120x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_12_bF$buf4),
    .Y(_3871_)
);

NAND3X1 _14026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3406_),
    .B(_3396_),
    .C(_3410_),
    .Y(_3411_)
);

FILL SFILL28920x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29160x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8840x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10564_),
    .B(_10568_),
    .C(_10571_),
    .Y(_10928_)
);

XOR2X1 _20464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10406_),
    .B(_10466_),
    .Y(_10467_)
);

OAI21X1 _20044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9662_),
    .B(_9653_),
    .C(_9657_),
    .Y(_10006_)
);

INVX2 _19484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9392_),
    .Y(_9393_)
);

NAND3X1 _19064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8892_),
    .B(_8931_),
    .C(_8930_),
    .Y(_8932_)
);

FILL SFILL59160x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11497_),
    .B(_11499_),
    .C(_11786_),
    .Y(_11787_)
);

NOR2X1 _21249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf2),
    .B(_7225__bF$buf4),
    .Y(_11327_)
);

INVX1 _12932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1586_),
    .Y(_1653_)
);

NOR2X1 _12512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf3),
    .B(_3646__bF$buf1),
    .Y(_8961_)
);

FILL SFILL28680x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_699_),
    .C(_909_),
    .Y(_910_)
);

OAI21X1 _13717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2815_),
    .B(_3071_),
    .C(_3072_),
    .Y(_3073_)
);

NAND2X1 _23815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2221_),
    .Y(_2222_)
);

OAI21X1 _16189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5434_),
    .B(_5432_),
    .C(_5423_),
    .Y(_5780_)
);

FILL FILL74040x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18760x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7728_),
    .B(_7716_),
    .C(_7720_),
    .Y(_7732_)
);

AOI21X1 _17550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(_6879_),
    .C(_6881_),
    .Y(_7271_)
);

OAI21X1 _17130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6502_),
    .B(_6504_),
    .C(_6506_),
    .Y(_6811_)
);

FILL SFILL38760x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8483_),
    .B(_8587_),
    .C(_8592_),
    .Y(_8593_)
);

OR2X2 _18335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8126_),
    .B(_8127_),
    .Y(_8133_)
);

NAND2X1 _13890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_15_bF$buf1),
    .Y(_3262_)
);

NOR2X1 _13470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2393_),
    .B(_2801_),
    .Y(_2802_)
);

NAND2X1 _13050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .B(_2344_),
    .Y(_2345_)
);

NAND3X1 _14675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4099_),
    .B(_4120_),
    .C(_4113_),
    .Y(_4121_)
);

INVX2 _14255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3641_),
    .Y(_3662_)
);

FILL SFILL44040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10712_),
    .B(_10717_),
    .C(_10705_),
    .Y(_10718_)
);

NOR2X1 _20273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9901_),
    .B(_10257_),
    .Y(_10258_)
);

AOI21X1 _16821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6159_),
    .B(_6157_),
    .C(_6471_),
    .Y(_6473_)
);

AOI21X1 _16401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6007_),
    .B(_6008_),
    .C(_6006_),
    .Y(_6013_)
);

NAND2X1 _19293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9176_),
    .B(_9183_),
    .Y(_9184_)
);

NAND2X1 _21898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf2),
    .B(areg_27_bF$buf0),
    .Y(_130_)
);

AOI21X1 _21478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11570_),
    .B(_11578_),
    .C(_11320_),
    .Y(_11579_)
);

NAND3X1 _21058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11115_),
    .B(_11117_),
    .C(_11111_),
    .Y(_11118_)
);

AOI21X1 _17606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6923_),
    .B(_7008_),
    .C(_7332_),
    .Y(_7333_)
);

FILL SFILL69240x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10002_),
    .B(_11297_),
    .C(_11361_),
    .Y(_11472_)
);

NAND3X1 _12321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6714_),
    .B(_6658_),
    .C(_6692_),
    .Y(_6867_)
);

FILL SFILL34040x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3323_),
    .Y(_3324_)
);

NOR2X1 _13526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2863_),
    .B(_2641_),
    .Y(_2864_)
);

NAND2X1 _13106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2400_),
    .Y(_2404_)
);

NOR2X1 _23624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .B(_2015_),
    .Y(_2016_)
);

NAND2X1 _23204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1414_),
    .B(_1425_),
    .Y(_1558_)
);

FILL FILL74200x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8825_),
    .B(_8832_),
    .C(_8835_),
    .Y(_8844_)
);

AOI21X1 _18564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8383_),
    .B(_8380_),
    .C(_8360_),
    .Y(_8384_)
);

NOR3X1 _18144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7913_),
    .B(_7914_),
    .C(_7908_),
    .Y(_7924_)
);

FILL SFILL59160x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10775_),
    .B(_10776_),
    .C(_10778_),
    .Y(_10779_)
);

OAI21X1 _20329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10314_),
    .B(_10315_),
    .C(_9995_),
    .Y(_10319_)
);

AOI21X1 _19769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9700_),
    .B(_9699_),
    .C(_9698_),
    .Y(_9705_)
);

NAND3X1 _19349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8886_),
    .B(_9241_),
    .C(_9242_),
    .Y(_9245_)
);

NAND2X1 _14484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3907_),
    .B(_3912_),
    .Y(_3913_)
);

OAI21X1 _14064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3441_),
    .C(_3358_),
    .Y(_3453_)
);

FILL SFILL69160x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5226_),
    .B(_5225_),
    .C(_5224_),
    .Y(_5231_)
);

XOR2X1 _15269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4723_),
    .B(_4771_),
    .Y(_4772_)
);

NAND2X1 _20082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_24_bF$buf3),
    .Y(_10048_)
);

FILL SFILL18760x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5953_),
    .B(_5949_),
    .C(_5915_),
    .Y(_6263_)
);

OAI21X1 _16210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5799_),
    .B(_5800_),
    .C(_5802_),
    .Y(_5803_)
);

FILL SFILL33960x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11101_),
    .B(_11098_),
    .C(_11091_),
    .Y(_11369_)
);

AOI21X1 _17835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7062_),
    .B(_7155_),
    .C(_7584_),
    .Y(_7585_)
);

NAND3X1 _17415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf4),
    .B(areg_29_bF$buf5),
    .C(_7124_),
    .Y(_7125_)
);

OAI21X1 _12970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2034_),
    .B(_2045_),
    .C(_2055_),
    .Y(_2066_)
);

AND2X2 _12550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8895_),
    .B(_8928_),
    .Y(_9378_)
);

AOI21X1 _12130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4632_),
    .B(_4588_),
    .C(_4226_),
    .Y(_4774_)
);

FILL SFILL23960x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3107_),
    .B(_3108_),
    .C(_3100_),
    .Y(_3115_)
);

AOI21X1 _23853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_2213_),
    .C(_2261_),
    .Y(_2262_)
);

NAND2X1 _13335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_13_bF$buf1),
    .Y(_2655_)
);

OAI21X1 _23433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .B(_1702_),
    .C(_1807_),
    .Y(_1808_)
);

XNOR2X1 _23013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1349_),
    .B(_1346_),
    .Y(_1350_)
);

NAND2X1 _15901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5121_),
    .B(_5129_),
    .Y(_5465_)
);

OR2X2 _18793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8629_),
    .B(_8634_),
    .Y(_8635_)
);

AOI21X1 _18373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8170_),
    .B(_8169_),
    .C(_8168_),
    .Y(_8175_)
);

FILL SFILL69320x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_11030_)
);

NAND2X1 _20558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_30_bF$buf2),
    .Y(_10570_)
);

OAI21X1 _20138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9854_),
    .B(_9943_),
    .C(_9934_),
    .Y(_10109_)
);

FILL SFILL69240x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9594_),
    .B(_9596_),
    .C(_9955_),
    .Y(_9956_)
);

NAND3X1 _19578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9491_),
    .B(_9495_),
    .C(_9494_),
    .Y(_9496_)
);

NOR3X1 _19158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9029_),
    .B(_9031_),
    .C(_9030_),
    .Y(_9035_)
);

NAND3X1 _14293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3698_),
    .B(_3697_),
    .C(_3696_),
    .Y(_3704_)
);

INVX1 _12606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8676_),
    .Y(_9991_)
);

NAND2X1 _22704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .B(_999_),
    .Y(_1013_)
);

NOR2X1 _15498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4694_),
    .B(_5021_),
    .Y(_5022_)
);

NAND3X1 _15078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4558_),
    .B(_4528_),
    .C(_4562_),
    .Y(_4563_)
);

BUFX2 _23909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[27]),
    .Y(y[27])
);

FILL FILL74200x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11138_),
    .B(_11159_),
    .C(_11151_),
    .Y(_11160_)
);

NAND3X1 _17644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7368_),
    .B(_7352_),
    .C(_7369_),
    .Y(_7375_)
);

NAND2X1 _17224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6493_),
    .B(_6499_),
    .Y(_6915_)
);

NAND2X1 _18849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_8696_)
);

NOR2X1 _18429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7838_),
    .B(_7884_),
    .Y(_8236_)
);

AND2X2 _18009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7321_),
    .B(_7314_),
    .Y(_7775_)
);

AND2X2 _13984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_13_bF$buf0),
    .Y(_3365_)
);

FILL FILL74200x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2905_),
    .B(_2904_),
    .C(_2896_),
    .Y(_2906_)
);

NAND3X1 _13144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2443_),
    .B(_2445_),
    .C(_2444_),
    .Y(_2446_)
);

NAND2X1 _23662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2002_),
    .B(_2025_),
    .Y(_2057_)
);

NOR2X1 _23242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1590_),
    .Y(_1600_)
);

AOI21X1 _14769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4212_),
    .B(_4211_),
    .C(_4208_),
    .Y(_4224_)
);

AOI21X1 _14349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3764_),
    .B(_3763_),
    .C(_3480_),
    .Y(_3765_)
);

DFFPOSX1 _24027_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[17]),
    .CLK(clk_bF$buf5),
    .D(a[17])
);

OAI21X1 _15710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5253_),
    .B(_5254_),
    .C(_5252_),
    .Y(_5255_)
);

OAI21X1 _18182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7529_),
    .B(_7533_),
    .C(_7532_),
    .Y(_7966_)
);

OAI21X1 _20787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10487_),
    .B(_10470_),
    .C(_10478_),
    .Y(_10821_)
);

AND2X2 _20367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_27_bF$buf5),
    .Y(_10360_)
);

NAND3X1 _16915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6573_),
    .B(_6574_),
    .C(_6575_),
    .Y(_6576_)
);

INVX2 _19387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9285_),
    .Y(_9286_)
);

OAI21X1 _12835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10902_),
    .B(_582_),
    .C(_560_),
    .Y(_593_)
);

NOR3X1 _12415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7843_),
    .B(_7832_),
    .C(_7854_),
    .Y(_7898_)
);

OAI21X1 _22933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1126_),
    .B(_1106_),
    .C(_1128_),
    .Y(_1263_)
);

OAI21X1 _22513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .B(_791_),
    .C(_787_),
    .Y(_804_)
);

AOI21X1 _23718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2052_),
    .B(_2103_),
    .C(_2116_),
    .Y(_2117_)
);

AOI21X1 _17873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7611_),
    .B(_7616_),
    .C(_7221_),
    .Y(_7627_)
);

AOI21X1 _17453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7161_),
    .B(_7160_),
    .C(_7159_),
    .Y(_7167_)
);

NOR2X1 _17033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6704_),
    .B(_6705_),
    .Y(_6706_)
);

OAI21X1 _18658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8099_),
    .B(_8085_),
    .C(_8109_),
    .Y(_8486_)
);

NAND3X1 _18238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7768_),
    .B(_7773_),
    .C(_7775_),
    .Y(_8026_)
);

AOI21X1 _13793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2879_),
    .B(_2885_),
    .C(_2887_),
    .Y(_3157_)
);

NAND3X1 _13373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2696_),
    .B(_2695_),
    .C(_2693_),
    .Y(_2697_)
);

BUFX2 _23891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[9]),
    .Y(y[9])
);

NAND3X1 _23471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(_1778_),
    .C(_1845_),
    .Y(_1850_)
);

OAI21X1 _23051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .B(_1390_),
    .C(_1262_),
    .Y(_1392_)
);

OAI21X1 _14998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4472_),
    .B(_4473_),
    .C(_4469_),
    .Y(_4474_)
);

NAND3X1 _14578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4014_),
    .B(_4015_),
    .C(_4013_),
    .Y(_4016_)
);

OAI21X1 _14158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3262_),
    .B(_3554_),
    .C(_3544_),
    .Y(_3555_)
);

FILL SFILL64200x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10611_),
    .B(_10610_),
    .C(_10550_),
    .Y(_10612_)
);

OAI21X1 _20176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_4541__bF$buf0),
    .C(_10143_),
    .Y(_10151_)
);

AOI21X1 _16724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6361_),
    .B(_6360_),
    .C(_6359_),
    .Y(_6367_)
);

OAI21X1 _16304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5906_),
    .B(_5901_),
    .C(_5888_),
    .Y(_5907_)
);

NAND3X1 _19196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9072_),
    .B(_9073_),
    .C(_9076_),
    .Y(_9077_)
);

OAI21X1 _17929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf4),
    .B(_5668__bF$buf3),
    .C(_7674_),
    .Y(_7687_)
);

NOR2X1 _17509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf2),
    .B(_7225__bF$buf1),
    .Y(_7226_)
);

NAND3X1 _12644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8654_),
    .B(_10397_),
    .C(_10386_),
    .Y(_10408_)
);

NAND3X1 _12224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4981_),
    .B(_5793_),
    .C(_5760_),
    .Y(_5804_)
);

NOR2X1 _22742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .B(_868_),
    .Y(_1055_)
);

OAI21X1 _22322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(_590_),
    .C(_542_),
    .Y(_595_)
);

AOI21X1 _13849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3212_),
    .B(_3217_),
    .C(_2985_),
    .Y(_3218_)
);

INVX2 _13429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2756_),
    .Y(_2757_)
);

DFFPOSX1 _23947_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[1]),
    .CLK(clk_bF$buf8),
    .D(_0_[1])
);

OAI21X1 _13009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2303_),
    .C(_2300_),
    .Y(_2304_)
);

XNOR2X1 _23527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1908_),
    .B(_1903_),
    .Y(_1909_)
);

NAND3X1 _23107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_23_bF$buf2),
    .B(areg_27_bF$buf5),
    .C(_1349_),
    .Y(_1452_)
);

OAI21X1 _17682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7412_),
    .B(_7411_),
    .C(_7379_),
    .Y(_7417_)
);

NOR2X1 _17262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6951_),
    .B(_6956_),
    .Y(_6957_)
);

FILL SFILL34120x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8727_),
    .B(_8728_),
    .C(_8723_),
    .Y(_8738_)
);

OAI21X1 _18467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8277_),
    .B(_8276_),
    .C(_8275_),
    .Y(_8278_)
);

OAI21X1 _18047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7405_),
    .B(_7402_),
    .C(_7395_),
    .Y(_7817_)
);

OAI21X1 _13182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2487_),
    .B(_2480_),
    .C(_2447_),
    .Y(_2488_)
);

NAND3X1 _23280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(_1638_),
    .C(_1551_),
    .Y(_1641_)
);

OR2X2 _11915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2419_),
    .Y(_2420_)
);

AND2X2 _14387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .B(_3805_),
    .Y(_3806_)
);

DFFPOSX1 _24065_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[23]),
    .CLK(clk_bF$buf5),
    .D(b[23])
);

FILL SFILL74280x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_20_bF$buf2),
    .Y(_6618_)
);

XNOR2X1 _16533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6135_),
    .B(_6131_),
    .Y(_6157_)
);

OAI21X1 _16113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf0),
    .B(_3781__bF$buf0),
    .C(_5372_),
    .Y(_5697_)
);

NAND2X1 _17738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7038_),
    .B(_7044_),
    .Y(_7478_)
);

NAND2X1 _17318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf3),
    .B(areg_16_bF$buf1),
    .Y(_7017_)
);

AOI21X1 _12873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_987_),
    .C(_921_),
    .Y(_1009_)
);

AOI21X1 _12453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8183_),
    .B(_8227_),
    .C(_8249_),
    .Y(_8315_)
);

NOR2X1 _22971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf1),
    .B(_5676_),
    .Y(_1304_)
);

NAND2X1 _12033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3591_),
    .B(_3701_),
    .Y(_3712_)
);

OR2X2 _22551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_844_),
    .B(_840_),
    .Y(_846_)
);

AOI21X1 _22131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_380_),
    .B(_384_),
    .C(_376_),
    .Y(_386_)
);

NOR2X1 _13658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .B(_2994_),
    .Y(_3008_)
);

AOI21X1 _13238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2547_),
    .C(_2341_),
    .Y(_2548_)
);

INVX2 _23756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2158_),
    .Y(_2159_)
);

NAND2X1 _23336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_26_bF$buf1),
    .B(areg_27_bF$buf4),
    .Y(_1702_)
);

FILL SFILL43720x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7205_),
    .B(_7206_),
    .C(_7204_),
    .Y(_7208_)
);

NAND3X1 _17071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6728_),
    .B(_6734_),
    .C(_6738_),
    .Y(_6748_)
);

AOI21X1 _15804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5009_),
    .B(_5098_),
    .C(_5095_),
    .Y(_5358_)
);

NAND2X1 _18696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8140_),
    .B(_8144_),
    .Y(_8528_)
);

NOR3X1 _18276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8054_),
    .B(_8057_),
    .C(_8060_),
    .Y(_8068_)
);

FILL SFILL33720x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11720_),
    .B(_46_),
    .C(_11722_),
    .Y(_47_)
);

AOI21X1 _21402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11489_),
    .B(_11495_),
    .C(_11475_),
    .Y(_11496_)
);

XOR2X1 _14196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3596_),
    .Y(_3597_)
);

FILL SFILL13640x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1587_),
    .B(_1598_),
    .C(_1609_),
    .Y(_1620_)
);

NAND3X1 _12509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8720_),
    .B(_8917_),
    .C(_8906_),
    .Y(_8928_)
);

AOI21X1 _22607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_906_),
    .C(_726_),
    .Y(_907_)
);

AOI21X1 _16762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6408_),
    .B(_6406_),
    .C(_6400_),
    .Y(_6409_)
);

NAND3X1 _16342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5941_),
    .B(_5948_),
    .C(_5928_),
    .Y(_5949_)
);

FILL SFILL23720x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert260 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .Y(_6300__bF$buf2)
);

BUFX2 BUFX2_insert261 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .Y(_6300__bF$buf1)
);

BUFX2 BUFX2_insert262 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .Y(_6300__bF$buf0)
);

BUFX2 BUFX2_insert263 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf5)
);

OAI21X1 _17967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7726_),
    .B(_7725_),
    .C(_7728_),
    .Y(_7729_)
);

BUFX2 BUFX2_insert264 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf4)
);

NAND3X1 _17547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7255_),
    .B(_7258_),
    .C(_7231_),
    .Y(_7268_)
);

BUFX2 BUFX2_insert265 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf3)
);

BUFX2 BUFX2_insert266 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf2)
);

NOR2X1 _17127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6804_),
    .B(_6807_),
    .Y(_6808_)
);

BUFX2 BUFX2_insert267 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf1)
);

BUFX2 BUFX2_insert268 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[24]),
    .Y(breg_24_bF$buf0)
);

INVX2 _12682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10814_),
    .Y(_10825_)
);

BUFX2 BUFX2_insert269 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217_),
    .Y(_7217__bF$buf4)
);

NAND2X1 _12262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_6_bF$buf2),
    .Y(_6220_)
);

AOI21X1 _22780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_942_),
    .C(_1094_),
    .Y(_1095_)
);

XNOR2X1 _22360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .B(_635_),
    .Y(_636_)
);

FILL SFILL8680x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3258_),
    .B(_3015_),
    .C(_3005_),
    .Y(_3259_)
);

DFFPOSX1 _23985_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[39]),
    .CLK(clk_bF$buf3),
    .D(_0_[39])
);

OAI21X1 _13467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2796_),
    .C(_2798_),
    .Y(_2799_)
);

OAI21X1 _13047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2338_),
    .B(_2339_),
    .C(_1423_),
    .Y(_2342_)
);

INVX1 _23565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7644_),
    .Y(_1951_)
);

NAND3X1 _23145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1492_),
    .B(_1493_),
    .C(_1491_),
    .Y(_1494_)
);

FILL SFILL48840x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4871_),
    .B(_4877_),
    .C(_4847_),
    .Y(_5149_)
);

AOI21X1 _18085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7857_),
    .B(_7858_),
    .C(_7812_),
    .Y(_7859_)
);

OAI21X1 _16818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6459_),
    .B(_6460_),
    .C(_6457_),
    .Y(_6469_)
);

OAI21X1 _11953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_2825__bF$buf2),
    .C(_2540_),
    .Y(_2836_)
);

AOI21X1 _21631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11740_),
    .B(_11744_),
    .C(_11726_),
    .Y(_11746_)
);

NAND3X1 _21211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11280_),
    .B(_11014_),
    .C(_11283_),
    .Y(_11287_)
);

FILL SFILL64280x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9554_),
    .B(_11428_),
    .Y(_11439_)
);

NAND3X1 _12318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6780_),
    .B(_6823_),
    .C(_6110_),
    .Y(_6834_)
);

INVX1 _22836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1049_),
    .Y(_1157_)
);

NAND3X1 _22416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_497_),
    .B(_687_),
    .C(_695_),
    .Y(_698_)
);

FILL SFILL33800x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6653_),
    .B(_6657_),
    .C(_6656_),
    .Y(_6660_)
);

OAI21X1 _16571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6196_),
    .B(_6197_),
    .C(_6193_),
    .Y(_6199_)
);

INVX1 _16151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .Y(_5739_)
);

INVX8 _17776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_28_bF$buf1),
    .Y(_7520_)
);

OAI21X1 _17356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .B(_7053_),
    .C(_7050_),
    .Y(_7060_)
);

INVX1 _12491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8720_),
    .Y(_8731_)
);

NAND2X1 _12071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg_6_bF$buf2),
    .Y(_4127_)
);

OAI21X1 _20902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10941_),
    .B(_10942_),
    .C(_10258_),
    .Y(_10948_)
);

FILL SFILL54200x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2805_),
    .B(_2810_),
    .C(_2829_),
    .Y(_3050_)
);

XNOR2X1 _13276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2589_),
    .B(_2582_),
    .Y(_2590_)
);

INVX1 _23794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .Y(_2200_)
);

OAI21X1 _23374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1739_),
    .C(_1735_),
    .Y(_1744_)
);

NOR2X1 _19922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9865_),
    .B(_9866_),
    .Y(_9874_)
);

NAND3X1 _19502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9407_),
    .B(_9399_),
    .C(_9412_),
    .Y(_9413_)
);

XNOR2X1 _15842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5377_),
    .B(_5370_),
    .Y(_5400_)
);

AOI21X1 _15422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4934_),
    .B(_4935_),
    .C(_4933_),
    .Y(_4941_)
);

OAI21X1 _15002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4472_),
    .B(_4473_),
    .C(_4454_),
    .Y(_4480_)
);

FILL SFILL44200x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf3),
    .B(_5921__bF$buf2),
    .C(_2560__bF$buf1),
    .D(_4541__bF$buf0),
    .Y(_10505_)
);

OAI21X1 _20079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9695_),
    .B(_9691_),
    .C(_9699_),
    .Y(_10044_)
);

NAND3X1 _16627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6244_),
    .B(_6249_),
    .C(_6250_),
    .Y(_6260_)
);

AOI21X1 _16207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5788_),
    .B(_5787_),
    .C(_5784_),
    .Y(_5800_)
);

AND2X2 _21860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11696_),
    .B(_11691_),
    .Y(_88_)
);

OR2X2 _21440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11524_),
    .B(_11535_),
    .Y(_11537_)
);

FILL SFILL38840x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11070_),
    .B(_11069_),
    .C(_11068_),
    .Y(_11076_)
);

NOR3X1 _19099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8619_),
    .B(_8622_),
    .C(_8616_),
    .Y(_8970_)
);

FILL SFILL44120x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2023_),
    .B(_1925_),
    .Y(_2034_)
);

AOI21X1 _12547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9225_),
    .B(_9181_),
    .C(_9027_),
    .Y(_9345_)
);

OAI21X1 _12127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4610_),
    .B(_4621_),
    .C(_4237_),
    .Y(_4741_)
);

INVX1 _22645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_947_),
    .Y(_948_)
);

AOI21X1 _22225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_487_),
    .B(_485_),
    .C(_486_),
    .Y(_488_)
);

NAND3X1 _16380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5746_),
    .B(_5833_),
    .C(_5832_),
    .Y(_5989_)
);

FILL SFILL38920x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(_6866_),
    .Y(_7310_)
);

OAI21X1 _17165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6442_),
    .B(_6849_),
    .C(_6451_),
    .Y(_6850_)
);

FILL SFILL3560x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10701_),
    .B(_10729_),
    .C(_10725_),
    .Y(_10738_)
);

NAND2X1 _13085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_13_bF$buf0),
    .Y(_2381_)
);

NAND3X1 _23183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .B(_1535_),
    .C(_1532_),
    .Y(_1536_)
);

FILL SFILL28920x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9662_),
    .B(_9661_),
    .C(_9653_),
    .Y(_9664_)
);

NAND3X1 _19311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9202_),
    .B(_9198_),
    .C(_9199_),
    .Y(_9204_)
);

AOI21X1 _21916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_149_),
    .C(_129_),
    .Y(_150_)
);

AND2X2 _15651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5183_),
    .B(_5184_),
    .Y(_5191_)
);

OAI21X1 _15231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf2),
    .B(_2586__bF$buf3),
    .C(_4450_),
    .Y(_4731_)
);

FILL SFILL28840x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6373_),
    .B(_6510_),
    .C(_6364_),
    .Y(_6511_)
);

INVX8 _16436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_28_bF$buf2),
    .Y(_6050_)
);

NAND3X1 _16016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5590_),
    .B(_5589_),
    .C(_5588_),
    .Y(_5591_)
);

NOR2X1 _11991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3055_),
    .B(_3241_),
    .Y(_3252_)
);

FILL SFILL54200x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11822_),
    .B(_11844_),
    .Y(_11855_)
);

AND2X2 _12356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7207_),
    .B(_7239_),
    .Y(_7250_)
);

AND2X2 _22874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1198_),
    .Y(_1199_)
);

INVX1 _22454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .Y(_739_)
);

OAI21X1 _22034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_271_),
    .C(_256_),
    .Y(_279_)
);

FILL SFILL18840x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2052_),
    .B(_2050_),
    .Y(_2053_)
);

NAND3X1 _23239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(_1595_),
    .C(_1593_),
    .Y(_1596_)
);

NAND2X1 _14922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_17_bF$buf4),
    .Y(_4392_)
);

OAI21X1 _14502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3929_),
    .B(_3674_),
    .C(_3932_),
    .Y(_3933_)
);

NAND3X1 _17394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7095_),
    .B(_7101_),
    .C(_7099_),
    .Y(_7102_)
);

FILL SFILL48920x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5250_),
    .B(_5251_),
    .Y(_5252_)
);

NAND3X1 _20940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10985_),
    .B(_10692_),
    .C(_10986_),
    .Y(_10989_)
);

AOI21X1 _20520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10144_),
    .B(_10166_),
    .C(_10170_),
    .Y(_10528_)
);

NAND3X1 _20100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10063_),
    .B(_10051_),
    .C(_10055_),
    .Y(_10067_)
);

OAI21X1 _18599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8415_),
    .B(_8421_),
    .C(_8187_),
    .Y(_8422_)
);

AOI22X1 _18179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_29_bF$buf0),
    .C(breg_4_bF$buf1),
    .D(areg_28_bF$buf5),
    .Y(_7962_)
);

XOR2X1 _19960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9911_),
    .B(_9902_),
    .Y(_9914_)
);

AOI21X1 _19540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9452_),
    .B(_9453_),
    .C(_9451_),
    .Y(_9454_)
);

AOI21X1 _19120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8979_),
    .B(_8984_),
    .C(_8933_),
    .Y(_8993_)
);

OAI21X1 _21725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11845_),
    .B(_11848_),
    .C(_11599_),
    .Y(_11849_)
);

NOR3X1 _21305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11372_),
    .B(_11377_),
    .C(_11376_),
    .Y(_11389_)
);

NAND3X1 _14099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3490_),
    .B(_3235_),
    .C(_3487_),
    .Y(_3491_)
);

AOI21X1 _15880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5423_),
    .B(_5429_),
    .C(_5407_),
    .Y(_5441_)
);

INVX2 _15460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4979_),
    .Y(_4980_)
);

NAND3X1 _15040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4515_),
    .B(_4520_),
    .C(_4501_),
    .Y(_4521_)
);

FILL SFILL38920x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6295_),
    .B(_6301_),
    .C(_6299_),
    .Y(_6302_)
);

NAND2X1 _16245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_15_bF$buf2),
    .Y(_5842_)
);

FILL SFILL3560x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69240x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8478_),
    .B(_9707_),
    .C(_9751_),
    .Y(_9762_)
);

XOR2X1 _12165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4423_),
    .B(_5146_),
    .Y(_5157_)
);

OR2X2 _22683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_989_),
    .Y(_990_)
);

AOI21X1 _22263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_525_),
    .C(_504_),
    .Y(_530_)
);

FILL SFILL28920x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8647_),
    .B(_8648_),
    .C(_8639_),
    .Y(_8655_)
);

BUFX2 _23888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[6]),
    .Y(y[6])
);

OAI21X1 _23468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(_1843_),
    .C(_1745_),
    .Y(_1846_)
);

NAND3X1 _23048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1265_),
    .B(_1382_),
    .C(_1385_),
    .Y(_1388_)
);

NAND3X1 _14731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4175_),
    .B(_4181_),
    .C(_4162_),
    .Y(_4183_)
);

NAND2X1 _14311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3722_),
    .B(_3721_),
    .Y(_3724_)
);

AOI21X1 _15936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5152_),
    .B(_5172_),
    .C(_5502_),
    .Y(_5503_)
);

NAND2X1 _15516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_16_bF$buf2),
    .Y(_5042_)
);

NAND3X1 _21954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11889_),
    .B(_91_),
    .C(_90_),
    .Y(_192_)
);

NOR3X1 _21534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11624_),
    .B(_11609_),
    .C(_11631_),
    .Y(_11640_)
);

NAND3X1 _21114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11170_),
    .B(_11178_),
    .C(_11179_),
    .Y(_11180_)
);

FILL SFILL39240x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1050_),
    .B(_1049_),
    .Y(_1051_)
);

OAI21X1 _22319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(_590_),
    .C(_588_),
    .Y(_591_)
);

AND2X2 _16894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf1),
    .B(breg_15_bF$buf4),
    .Y(_6553_)
);

AOI21X1 _16474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6073_),
    .B(_6080_),
    .C(_6059_),
    .Y(_6092_)
);

OAI21X1 _16054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5631_),
    .B(_5632_),
    .C(_5630_),
    .Y(_5633_)
);

OAI21X1 _17679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7412_),
    .B(_7411_),
    .C(_7408_),
    .Y(_7413_)
);

NAND3X1 _17259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6948_),
    .B(_6949_),
    .C(_6932_),
    .Y(_6953_)
);

NAND2X1 _12394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf3),
    .B(areg_8_bF$buf1),
    .Y(_7667_)
);

INVX1 _22492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .Y(_781_)
);

INVX1 _22072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .Y(_321_)
);

OAI21X1 _18620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8429_),
    .B(_8436_),
    .C(_8439_),
    .Y(_8445_)
);

AOI21X1 _18200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7979_),
    .B(_7984_),
    .C(_7955_),
    .Y(_7985_)
);

FILL SFILL69080x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10840_),
    .B(_10839_),
    .C(_10822_),
    .Y(_10841_)
);

NAND3X1 _13599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2925_),
    .B(_2933_),
    .C(_2937_),
    .Y(_2944_)
);

AOI21X1 _13179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2482_),
    .C(_2476_),
    .Y(_2484_)
);

NAND2X1 _23697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .B(_2093_),
    .Y(_2095_)
);

OAI21X1 _23277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1629_),
    .B(_1628_),
    .C(_1553_),
    .Y(_1638_)
);

INVX2 _19825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9766_),
    .Y(_9767_)
);

NAND3X1 _19405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9282_),
    .B(_9305_),
    .C(_9304_),
    .Y(_9306_)
);

NAND3X1 _14960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4431_),
    .B(_4432_),
    .C(_4427_),
    .Y(_4433_)
);

NOR2X1 _14540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .B(_3959_),
    .Y(_3974_)
);

OAI21X1 _14120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .B(_2977_),
    .C(_3512_),
    .Y(_3513_)
);

FILL SFILL3640x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5279_),
    .B(_5285_),
    .C(_5283_),
    .Y(_5294_)
);

NAND3X1 _15325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4824_),
    .B(_4828_),
    .C(_4833_),
    .Y(_4834_)
);

FILL SFILL59080x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf1),
    .B(_7225__bF$buf4),
    .Y(_11890_)
);

AOI21X1 _21343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11221_),
    .B(_11223_),
    .C(_11430_),
    .Y(_11431_)
);

NAND2X1 _22968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf1),
    .B(areg_26_bF$buf0),
    .Y(_1301_)
);

NOR2X1 _22548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_841_),
    .Y(_842_)
);

NOR2X1 _22128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_381_),
    .Y(_382_)
);

FILL SFILL49080x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(_3175_),
    .C(_3171_),
    .Y(_3177_)
);

NAND2X1 _16283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5883_),
    .B(_5878_),
    .Y(_5884_)
);

FILL SFILL39080x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6421_),
    .B(_6786_),
    .C(_7203_),
    .Y(_7204_)
);

OAI21X1 _17068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6642_),
    .B(_6638_),
    .C(_6644_),
    .Y(_6744_)
);

FILL SFILL39000x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10108_),
    .B(_10290_),
    .C(_10631_),
    .Y(_10632_)
);

XOR2X1 _23086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(_1414_),
    .Y(_1429_)
);

NOR3X1 _19634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9546_),
    .B(_9531_),
    .C(_9547_),
    .Y(_9558_)
);

OAI21X1 _19214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8740_),
    .B(_8822_),
    .C(_8799_),
    .Y(_9096_)
);

AOI21X1 _21819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_37_),
    .C(_36_),
    .Y(_43_)
);

FILL SFILL8760x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_22_bF$buf0),
    .Y(_5545_)
);

OAI21X1 _15554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5082_),
    .B(_5083_),
    .C(_5017_),
    .Y(_5084_)
);

NAND3X1 _15134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4350_),
    .B(_4618_),
    .C(_4624_),
    .Y(_4625_)
);

AOI21X1 _16759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5666_),
    .B(_6015_),
    .C(_6018_),
    .Y(_6405_)
);

AOI21X1 _16339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5943_),
    .B(_5944_),
    .C(_5930_),
    .Y(_5945_)
);

NAND3X1 _21992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_233_),
    .C(_230_),
    .Y(_234_)
);

AOI21X1 _21572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11664_),
    .B(_11670_),
    .C(_11649_),
    .Y(_11681_)
);

NAND3X1 _21152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11205_),
    .B(_11217_),
    .C(_11210_),
    .Y(_11222_)
);

OAI21X1 _17700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7159_),
    .B(_7435_),
    .C(_7149_),
    .Y(_7436_)
);

XNOR2X1 _12679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10781_),
    .B(_10726_),
    .Y(_10792_)
);

NAND2X1 _12259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_4_bF$buf5),
    .Y(_6187_)
);

NAND2X1 _22777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1092_),
    .Y(_1093_)
);

NAND3X1 _22357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .B(_632_),
    .C(_631_),
    .Y(_633_)
);

FILL SFILL3720x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8749_),
    .B(_8748_),
    .C(_8746_),
    .Y(_8758_)
);

NAND3X1 _13620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2965_),
    .C(_2966_),
    .Y(_2967_)
);

NOR3X1 _13200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2318_),
    .B(_2319_),
    .C(_2320_),
    .Y(_2507_)
);

NAND2X1 _16092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_24_bF$buf5),
    .Y(_5674_)
);

OAI21X1 _14825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4284_),
    .B(_4285_),
    .C(_4283_),
    .Y(_4286_)
);

INVX1 _14405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3811_),
    .Y(_3826_)
);

AOI21X1 _17297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6983_),
    .B(_6978_),
    .C(_6960_),
    .Y(_6995_)
);

AOI21X1 _20843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10499_),
    .B(_10521_),
    .C(_10524_),
    .Y(_10883_)
);

NAND3X1 _20423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10418_),
    .B(_10420_),
    .C(_10421_),
    .Y(_10422_)
);

NAND3X1 _20003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9957_),
    .B(_9958_),
    .C(_9644_),
    .Y(_9962_)
);

AOI21X1 _19863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9801_),
    .B(_9802_),
    .C(_9794_),
    .Y(_9809_)
);

OAI21X1 _19443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9034_),
    .B(_9036_),
    .C(_9028_),
    .Y(_9348_)
);

NAND2X1 _19023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8587_),
    .B(_8593_),
    .Y(_8887_)
);

FILL SFILL33880x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11736_),
    .B(_11738_),
    .C(_11737_),
    .Y(_11742_)
);

OAI21X1 _21208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11281_),
    .B(_11282_),
    .C(_11130_),
    .Y(_11283_)
);

OAI21X1 _15783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5326_),
    .B(_5327_),
    .C(_5324_),
    .Y(_5335_)
);

NAND3X1 _15363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4867_),
    .B(_4865_),
    .C(_4861_),
    .Y(_4876_)
);

FILL SFILL18600x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .B(areg_23_bF$buf2),
    .Y(_6655_)
);

OAI21X1 _16568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6181_),
    .B(_6182_),
    .C(_6179_),
    .Y(_6195_)
);

AOI21X1 _16148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5368_),
    .B(_5458_),
    .C(_5455_),
    .Y(_5735_)
);

OAI21X1 _21381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11195_),
    .B(_11193_),
    .C(_11184_),
    .Y(_11473_)
);

FILL SFILL23880x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54280x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8687_),
    .B(_8676_),
    .Y(_8698_)
);

NOR2X1 _12068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3394_),
    .B(_4083_),
    .Y(_4094_)
);

AND2X2 _22586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .B(_877_),
    .Y(_884_)
);

FILL SFILL23800x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_420_),
    .C(_417_),
    .Y(_424_)
);

NOR2X1 _18714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8191_),
    .B(_8192_),
    .Y(_8548_)
);

FILL SFILL8760x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9864_),
    .B(_9869_),
    .C(_9867_),
    .Y(_9870_)
);

NAND2X1 _14634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf4),
    .B(breg_19_bF$buf3),
    .Y(_4076_)
);

OAI21X1 _14214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3615_),
    .B(_3616_),
    .C(_3601_),
    .Y(_3617_)
);

FILL SFILL74440x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5386_),
    .B(_5384_),
    .C(_5381_),
    .Y(_5396_)
);

NAND3X1 _15419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4656_),
    .B(_4932_),
    .C(_4936_),
    .Y(_4937_)
);

AOI22X1 _20652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10333_),
    .B(_10331_),
    .C(_10654_),
    .D(_10659_),
    .Y(_10673_)
);

NAND2X1 _20232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_26_bF$buf4),
    .Y(_10212_)
);

NOR3X1 _19672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9205_),
    .B(_9211_),
    .C(_9215_),
    .Y(_9600_)
);

NOR3X1 _19252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9128_),
    .B(_9129_),
    .C(_9123_),
    .Y(_9139_)
);

AOI21X1 _21857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11717_),
    .B(_11803_),
    .C(_11806_),
    .Y(_85_)
);

FILL SFILL3720x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _21437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11531_),
    .B(_11533_),
    .Y(_11534_)
);

AND2X2 _21017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10755_),
    .B(_10818_),
    .Y(_11073_)
);

FILL SFILL43960x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10957_),
    .B(_10979_),
    .C(_10968_),
    .Y(_11022_)
);

AOI21X1 _15592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5123_),
    .B(_5125_),
    .C(_5110_),
    .Y(_5126_)
);

XNOR2X1 _15172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4665_),
    .B(_4657_),
    .Y(_4666_)
);

NAND3X1 _13905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3260_),
    .B(_3273_),
    .C(_3278_),
    .Y(_3279_)
);

AND2X2 _16797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_25_bF$buf3),
    .Y(_6446_)
);

AOI21X1 _16377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5968_),
    .B(_5974_),
    .C(_5884_),
    .Y(_5986_)
);

AND2X2 _21190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11254_),
    .B(_11258_),
    .Y(_11263_)
);

OAI21X1 _12297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5146_),
    .B(_6571_),
    .C(_6593_),
    .Y(_6604_)
);

OAI21X1 _22395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_673_),
    .C(_500_),
    .Y(_674_)
);

OAI21X1 _18943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8783_),
    .B(_8789_),
    .C(_8791_),
    .Y(_8800_)
);

NAND2X1 _18523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8338_),
    .B(_8339_),
    .Y(_8340_)
);

AOI21X1 _18103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7559_),
    .B(_7565_),
    .C(_7485_),
    .Y(_7879_)
);

FILL SFILL33880x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _20708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10731_),
    .B(_10732_),
    .C(_10733_),
    .Y(_10734_)
);

NAND2X1 _19728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_28_bF$buf2),
    .Y(_9660_)
);

NOR2X1 _19308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9184_),
    .B(_9186_),
    .Y(_9200_)
);

OAI21X1 _14863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4323_),
    .B(_4324_),
    .C(_4059_),
    .Y(_4328_)
);

NAND2X1 _14443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3622_),
    .B(_3628_),
    .Y(_3868_)
);

NOR2X1 _14023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3403_),
    .B(_3407_),
    .Y(_3408_)
);

FILL SFILL23480x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .B(_5186_),
    .C(_5185_),
    .Y(_5187_)
);

AOI21X1 _15228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4720_),
    .B(_4721_),
    .C(_4712_),
    .Y(_4727_)
);

OAI21X1 _20881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_8773_),
    .C(_10565_),
    .Y(_10925_)
);

FILL SFILL23880x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf4),
    .B(breg_23_bF$buf1),
    .Y(_10464_)
);

OAI21X1 _20041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9665_),
    .B(_9650_),
    .C(_9675_),
    .Y(_10003_)
);

FILL SFILL44360x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9095_),
    .B(_9388_),
    .C(_9209_),
    .Y(_9390_)
);

OAI21X1 _19061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8927_),
    .B(_8923_),
    .C(_8893_),
    .Y(_8929_)
);

INVX4 _11988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf2),
    .Y(_3220_)
);

OAI21X1 _21666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11783_),
    .B(_11782_),
    .C(_11781_),
    .Y(_11784_)
);

INVX2 _21246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11323_),
    .Y(_11324_)
);

FILL SFILL74200x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3069_),
    .B(_3060_),
    .C(_3067_),
    .Y(_3070_)
);

OAI21X1 _23812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2216_),
    .B(_2182_),
    .C(_2218_),
    .Y(_2219_)
);

FILL SFILL29000x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .B(_5764_),
    .C(_5766_),
    .Y(_5777_)
);

AND2X2 _14919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4386_),
    .B(_4387_),
    .Y(_4388_)
);

AOI21X1 _18752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8572_),
    .B(_8580_),
    .C(_8525_),
    .Y(_8590_)
);

AND2X2 _18332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8126_),
    .B(_8127_),
    .Y(_8130_)
);

NAND3X1 _20937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10695_),
    .B(_10977_),
    .C(_10972_),
    .Y(_10986_)
);

AOI21X1 _20517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10506_),
    .B(_10510_),
    .C(_10513_),
    .Y(_10525_)
);

FILL SFILL43960x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9908_),
    .B(_9910_),
    .Y(_9911_)
);

OAI21X1 _19537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9065_),
    .B(_9432_),
    .C(_9048_),
    .Y(_9451_)
);

OAI21X1 _19117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8689_),
    .B(_8688_),
    .C(_8685_),
    .Y(_8990_)
);

AOI21X1 _14672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4115_),
    .B(_4117_),
    .C(_4114_),
    .Y(_4118_)
);

AOI22X1 _14252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3389_),
    .B(_3391_),
    .C(_3658_),
    .D(_3387_),
    .Y(_3659_)
);

NAND3X1 _15877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5428_),
    .B(_5415_),
    .C(_5418_),
    .Y(_5438_)
);

OAI22X1 _15457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4364_),
    .B(_4679_),
    .C(_4681_),
    .D(_4678_),
    .Y(_4977_)
);

INVX1 _15037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4239_),
    .Y(_4518_)
);

NOR2X1 _20690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10365_),
    .B(_10713_),
    .Y(_10714_)
);

AOI21X1 _20270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10252_),
    .B(_10253_),
    .C(_10251_),
    .Y(_10254_)
);

OAI21X1 _19290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9178_),
    .B(_9179_),
    .C(_9143_),
    .Y(_9180_)
);

OAI21X1 _21895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11783_),
    .B(_11781_),
    .C(_11770_),
    .Y(_127_)
);

AOI21X1 _21475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11564_),
    .B(_11561_),
    .C(_11325_),
    .Y(_11576_)
);

NAND3X1 _21055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11113_),
    .B(_11112_),
    .C(_11114_),
    .Y(_11115_)
);

AOI21X1 _17603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7324_),
    .B(_7323_),
    .C(_7322_),
    .Y(_7330_)
);

FILL SFILL54040x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_3961__bF$buf0),
    .C(_8243_),
    .Y(_8651_)
);

AOI21X1 _13943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3061_),
    .B(_3072_),
    .C(_3063_),
    .Y(_3321_)
);

OAI21X1 _13523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2860_),
    .B(_2859_),
    .C(_2854_),
    .Y(_2861_)
);

NAND2X1 _13103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2400_),
    .Y(_2401_)
);

NAND2X1 _23621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_27_bF$buf3),
    .B(areg_29_bF$buf4),
    .Y(_2013_)
);

OAI21X1 _23201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1479_),
    .B(_1481_),
    .C(_1470_),
    .Y(_1555_)
);

AOI21X1 _14728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4177_),
    .B(_4178_),
    .C(_4164_),
    .Y(_4179_)
);

AOI21X1 _14308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3715_),
    .B(_3719_),
    .C(_3638_),
    .Y(_3720_)
);

NAND3X1 _18981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8483_),
    .B(_8595_),
    .C(_8596_),
    .Y(_8841_)
);

AOI21X1 _18561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7974_),
    .B(_7977_),
    .C(_7971_),
    .Y(_8381_)
);

NAND3X1 _18141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7881_),
    .B(_7919_),
    .C(_7915_),
    .Y(_7921_)
);

AOI21X1 _20746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10758_),
    .B(_10765_),
    .C(_10743_),
    .Y(_10776_)
);

OAI21X1 _20326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10314_),
    .B(_10315_),
    .C(_10313_),
    .Y(_10316_)
);

FILL SFILL8840x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_22_bF$buf0),
    .Y(_9702_)
);

NAND3X1 _19346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8888_),
    .B(_9232_),
    .C(_9227_),
    .Y(_9242_)
);

AOI21X1 _14481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3903_),
    .B(_3904_),
    .C(_3905_),
    .Y(_3910_)
);

OAI21X1 _14061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .B(_3447_),
    .C(_3446_),
    .Y(_3450_)
);

FILL SFILL69560x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74520x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5223_),
    .B(_5227_),
    .C(_5150_),
    .Y(_5228_)
);

NAND2X1 _15266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4468_),
    .B(_4475_),
    .Y(_4769_)
);

FILL SFILL13800x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11330_),
    .B(_11356_),
    .C(_11353_),
    .Y(_11366_)
);

NAND3X1 _17832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7578_),
    .B(_7581_),
    .C(_7579_),
    .Y(_7582_)
);

NAND2X1 _17412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf4),
    .B(areg_29_bF$buf5),
    .Y(_7122_)
);

FILL SFILL49000x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL63880x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf0),
    .B(breg_25_bF$buf1),
    .Y(_777_)
);

AOI21X1 _22069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_316_),
    .C(_98_),
    .Y(_317_)
);

FILL SFILL64120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8440_),
    .B(_8441_),
    .C(_8439_),
    .Y(_8442_)
);

AND2X2 _13752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2872_),
    .B(_2873_),
    .Y(_3112_)
);

OAI21X1 _13332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2478_),
    .B(_2476_),
    .C(_2470_),
    .Y(_2652_)
);

NOR2X1 _23850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2242_),
    .Y(_2258_)
);

NAND2X1 _23430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1710_),
    .B(_1803_),
    .Y(_1804_)
);

NAND2X1 _23010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_23_bF$buf2),
    .B(areg_27_bF$buf5),
    .Y(_1346_)
);

FILL SFILL64040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4420_),
    .B(_4414_),
    .C(_4418_),
    .Y(_4430_)
);

NAND3X1 _14537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3965_),
    .B(_3967_),
    .C(_3966_),
    .Y(_3971_)
);

NAND3X1 _14117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_3497_),
    .C(_3238_),
    .Y(_3510_)
);

NAND3X1 _18790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8623_),
    .B(_8608_),
    .C(_8627_),
    .Y(_8631_)
);

NAND3X1 _18370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8168_),
    .B(_8170_),
    .C(_8169_),
    .Y(_8171_)
);

NAND2X1 _20975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11025_),
    .B(_11026_),
    .Y(_11027_)
);

AOI22X1 _20555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_30_bF$buf2),
    .C(breg_10_bF$buf4),
    .D(areg_29_bF$buf2),
    .Y(_10567_)
);

OAI21X1 _20135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10099_),
    .B(_10098_),
    .C(_10096_),
    .Y(_10106_)
);

AOI21X1 _19995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9952_),
    .B(_9951_),
    .C(_9950_),
    .Y(_9953_)
);

FILL SFILL54040x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_27_bF$buf2),
    .Y(_9493_)
);

OAI21X1 _19155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9030_),
    .B(_9031_),
    .C(_9029_),
    .Y(_9032_)
);

OAI21X1 _14290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3699_),
    .B(_3695_),
    .C(_3669_),
    .Y(_3700_)
);

FILL SFILL59240x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33880x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9641_),
    .Y(_9959_)
);

NAND3X1 _22701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_980_),
    .B(_1004_),
    .C(_1008_),
    .Y(_1010_)
);

INVX2 _15495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5018_),
    .Y(_5019_)
);

OAI21X1 _15075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4554_),
    .B(_4556_),
    .C(_4536_),
    .Y(_4560_)
);

NOR3X1 _13808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3155_),
    .B(_3157_),
    .C(_3149_),
    .Y(_3173_)
);

BUFX2 _23906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[24]),
    .Y(y[24])
);

FILL SFILL44040x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11144_),
    .B(_11141_),
    .Y(_11157_)
);

AOI21X1 _17641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7366_),
    .B(_7370_),
    .C(_7351_),
    .Y(_7372_)
);

AOI21X1 _17221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6512_),
    .B(_6597_),
    .C(_6594_),
    .Y(_6912_)
);

INVX1 _22298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .Y(_568_)
);

AOI21X1 _18846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8398_),
    .B(_8395_),
    .C(_8332_),
    .Y(_8693_)
);

OAI21X1 _18426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf0),
    .B(_2884__bF$buf3),
    .C(_8229_),
    .Y(_8233_)
);

AOI21X1 _18006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7430_),
    .B(_7428_),
    .C(_7771_),
    .Y(_7772_)
);

NAND2X1 _13981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_11_bF$buf0),
    .Y(_3362_)
);

AOI21X1 _13561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_2678_),
    .C(_2681_),
    .Y(_2903_)
);

NOR2X1 _13141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2424_),
    .B(_2034_),
    .Y(_2443_)
);

FILL SFILL69160x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4218_),
    .B(_3952_),
    .C(_4220_),
    .Y(_4221_)
);

FILL SFILL74120x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3753_),
    .B(_3761_),
    .C(_3517_),
    .Y(_3762_)
);

FILL SFILL28920x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24024_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[14]),
    .CLK(clk_bF$buf10),
    .D(a[14])
);

FILL SFILL8840x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf3),
    .B(breg_21_bF$buf1),
    .Y(_10818_)
);

NAND2X1 _20364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf0),
    .B(breg_29_bF$buf0),
    .Y(_10357_)
);

AOI21X1 _16912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5786_),
    .B(_6552_),
    .C(_6181_),
    .Y(_6573_)
);

INVX2 _19384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9282_),
    .Y(_9283_)
);

AOI21X1 _21989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11597_),
    .B(_11857_),
    .C(_11880_),
    .Y(_230_)
);

OAI21X1 _21569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11445_),
    .B(_11676_),
    .C(_11468_),
    .Y(_11677_)
);

OAI21X1 _21149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11214_),
    .B(_11215_),
    .C(_11217_),
    .Y(_11218_)
);

OAI21X1 _12832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_549__bF$buf4),
    .C(_516_),
    .Y(_560_)
);

OAI21X1 _12412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7854_),
    .B(_7843_),
    .C(_7832_),
    .Y(_7865_)
);

INVX1 _22930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1258_),
    .Y(_1259_)
);

OAI21X1 _22510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_616_),
    .C(_638_),
    .Y(_800_)
);

NAND3X1 _13617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2958_),
    .B(_2963_),
    .C(_2753_),
    .Y(_2964_)
);

OAI21X1 _23715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_1984_),
    .C(_2113_),
    .Y(_2114_)
);

AOI21X1 _16089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(_5336_),
    .C(_5341_),
    .Y(_5670_)
);

FILL FILL74040x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7617_),
    .B(_7220_),
    .C(_7621_),
    .Y(_7622_)
);

NAND3X1 _17450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7156_),
    .B(_7162_),
    .C(_7015_),
    .Y(_7163_)
);

NAND3X1 _17030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6696_),
    .B(_6701_),
    .C(_6699_),
    .Y(_6702_)
);

FILL SFILL54120x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8162_),
    .B(_8167_),
    .Y(_8483_)
);

NAND3X1 _18235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8005_),
    .B(_8011_),
    .C(_7878_),
    .Y(_8023_)
);

OAI21X1 _13790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf0),
    .B(_3146__bF$buf3),
    .C(_3152_),
    .Y(_3153_)
);

AND2X2 _13370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2645_),
    .B(_2649_),
    .Y(_2693_)
);

OAI21X1 _14995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_2287__bF$buf2),
    .C(_4457_),
    .Y(_4471_)
);

AOI21X1 _14575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3724_),
    .B(_3726_),
    .C(_3731_),
    .Y(_4013_)
);

INVX2 _14155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .Y(_3552_)
);

FILL SFILL44040x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10555_),
    .B(_10608_),
    .Y(_10609_)
);

AND2X2 _20173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_22_bF$buf3),
    .Y(_10148_)
);

NAND3X1 _16721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .B(_6219_),
    .C(_6362_),
    .Y(_6364_)
);

AOI21X1 _16301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5895_),
    .B(_5894_),
    .C(_5890_),
    .Y(_5904_)
);

NOR3X1 _19193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9058_),
    .B(_9055_),
    .C(_9057_),
    .Y(_9074_)
);

OAI21X1 _21798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_16_),
    .C(_15_),
    .Y(_20_)
);

OAI21X1 _21378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11454_),
    .B(_11458_),
    .C(_11460_),
    .Y(_11469_)
);

AOI21X1 _17926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7679_),
    .B(_7683_),
    .C(_7671_),
    .Y(_7684_)
);

OAI21X1 _17506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7187_),
    .B(_7222_),
    .C(_7177_),
    .Y(_7223_)
);

FILL SFILL69240x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10364_),
    .B(_10321_),
    .C(_8665_),
    .Y(_10375_)
);

OAI21X1 _12221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5738_),
    .B(_5727_),
    .C(_5716_),
    .Y(_5771_)
);

NAND3X1 _13846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3208_),
    .B(_3210_),
    .C(_3207_),
    .Y(_3215_)
);

AOI21X1 _13426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2721_),
    .B(_2718_),
    .C(_2556_),
    .Y(_2754_)
);

BUFX2 _23944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[62]),
    .Y(y[62])
);

NAND2X1 _13006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2292_),
    .B(_2289_),
    .Y(_2301_)
);

INVX2 _23524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .Y(_1906_)
);

OR2X2 _23104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1301_),
    .B(_1448_),
    .Y(_1449_)
);

FILL SFILL3800x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8695_),
    .B(_8734_),
    .C(_8729_),
    .Y(_8735_)
);

AND2X2 _18464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7868_),
    .B(_7862_),
    .Y(_8275_)
);

AOI21X1 _18044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7801_),
    .B(_7805_),
    .C(_7793_),
    .Y(_7814_)
);

FILL SFILL59160x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9251_),
    .B(_9258_),
    .Y(_10669_)
);

AND2X2 _20229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9884_),
    .B(_9876_),
    .Y(_10209_)
);

NOR2X1 _11912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_2376__bF$buf0),
    .Y(_2387_)
);

OAI21X1 _19669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9577_),
    .B(_9583_),
    .C(_9586_),
    .Y(_9596_)
);

NAND3X1 _19249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9097_),
    .B(_9134_),
    .C(_9130_),
    .Y(_9135_)
);

NAND2X1 _14384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3785_),
    .B(_3800_),
    .Y(_3803_)
);

DFFPOSX1 _24062_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[20]),
    .CLK(clk_bF$buf4),
    .D(b[20])
);

FILL SFILL9000x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4777_),
    .B(_4781_),
    .C(_4784_),
    .Y(_5122_)
);

AND2X2 _15169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4661_),
    .B(_4659_),
    .Y(_4662_)
);

FILL FILL74040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18760x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6229_),
    .B(_6613_),
    .Y(_6614_)
);

OAI21X1 _16530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6144_),
    .B(_6140_),
    .C(_6138_),
    .Y(_6153_)
);

OAI21X1 _16110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5315__bF$buf1),
    .C(_5678_),
    .Y(_5693_)
);

OAI21X1 _21187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10952_),
    .B(_11131_),
    .C(_11259_),
    .Y(_11260_)
);

AOI21X1 _17735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7086_),
    .B(_7083_),
    .C(_7088_),
    .Y(_7475_)
);

AOI21X1 _17315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6728_),
    .B(_6734_),
    .C(_6650_),
    .Y(_7014_)
);

AOI21X1 _12870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11264_),
    .B(_11253_),
    .C(_11231_),
    .Y(_976_)
);

AOI21X1 _12450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8260_),
    .B(_8271_),
    .C(_8249_),
    .Y(_8282_)
);

XNOR2X1 _12030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3668_),
    .B(_3624_),
    .Y(_3679_)
);

FILL SFILL23960x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2999_),
    .B(_3004_),
    .C(_2995_),
    .Y(_3005_)
);

AOI21X1 _13235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2537_),
    .B(_1412_),
    .C(_2544_),
    .Y(_2545_)
);

INVX1 _23753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2155_),
    .Y(_2156_)
);

INVX1 _23333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .Y(_1699_)
);

OAI21X1 _15801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5097_),
    .B(_5090_),
    .C(_5099_),
    .Y(_5355_)
);

AND2X2 _18693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8520_),
    .B(_8524_),
    .Y(_8525_)
);

NAND3X1 _18273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8060_),
    .B(_8061_),
    .C(_8065_),
    .Y(_8066_)
);

FILL SFILL69320x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_8773_),
    .C(_10570_),
    .Y(_10921_)
);

NAND2X1 _20458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10455_),
    .B(_10459_),
    .Y(_10460_)
);

AND2X2 _20038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9736_),
    .B(_9728_),
    .Y(_9999_)
);

FILL SFILL69240x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9844_),
    .B(_9843_),
    .C(_9846_),
    .Y(_9847_)
);

NAND3X1 _19478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9383_),
    .B(_9384_),
    .C(_9385_),
    .Y(_9386_)
);

AOI21X1 _19058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8920_),
    .B(_8921_),
    .C(_8896_),
    .Y(_8925_)
);

NOR2X1 _14193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf1),
    .B(_2379_),
    .Y(_3594_)
);

NAND2X1 _12926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_9_bF$buf2),
    .Y(_1587_)
);

OAI21X1 _12506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8884_),
    .B(_8852_),
    .C(_8731_),
    .Y(_8895_)
);

AOI21X1 _22604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_903_),
    .B(_898_),
    .C(_727_),
    .Y(_904_)
);

OAI21X1 _15398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4912_),
    .B(_4913_),
    .C(_4909_),
    .Y(_4914_)
);

OAI21X1 _23809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2169_),
    .B(_2193_),
    .C(_2214_),
    .Y(_2215_)
);

FILL SFILL59240x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert230 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf1)
);

BUFX2 BUFX2_insert231 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf0)
);

BUFX2 BUFX2_insert232 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[20]),
    .Y(areg_20_bF$buf4)
);

BUFX2 BUFX2_insert233 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[20]),
    .Y(areg_20_bF$buf3)
);

NOR3X1 _17964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7712_),
    .B(_7714_),
    .C(_7715_),
    .Y(_7726_)
);

BUFX2 BUFX2_insert234 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[20]),
    .Y(areg_20_bF$buf2)
);

NOR3X1 _17544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7262_),
    .B(_7263_),
    .C(_7264_),
    .Y(_7265_)
);

BUFX2 BUFX2_insert235 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[20]),
    .Y(areg_20_bF$buf1)
);

BUFX2 BUFX2_insert236 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[20]),
    .Y(areg_20_bF$buf0)
);

NOR2X1 _17124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6416_),
    .B(_6803_),
    .Y(_6805_)
);

BUFX2 BUFX2_insert237 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf5)
);

BUFX2 BUFX2_insert238 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf4)
);

BUFX2 BUFX2_insert239 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf3)
);

OAI21X1 _18749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8276_),
    .B(_8275_),
    .C(_8273_),
    .Y(_8586_)
);

NAND2X1 _18329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_25_bF$buf5),
    .Y(_8126_)
);

OAI21X1 _13884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2990_),
    .B(_3251_),
    .C(_3255_),
    .Y(_3256_)
);

FILL FILL74200x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23982_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[36]),
    .CLK(clk_bF$buf3),
    .D(_0_[36])
);

NAND2X1 _13464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_13_bF$buf0),
    .Y(_2796_)
);

AOI21X1 _13044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2331_),
    .C(_1467_),
    .Y(_2339_)
);

NAND2X1 _23562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_1943_),
    .Y(_1949_)
);

AND2X2 _23142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .B(_1324_),
    .Y(_1491_)
);

FILL SFILL33960x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4100_),
    .Y(_4114_)
);

AOI21X1 _14249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3650_),
    .B(_3651_),
    .C(_3649_),
    .Y(_3655_)
);

FILL SFILL18760x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5129_),
    .B(_5134_),
    .C(_5136_),
    .Y(_5145_)
);

AOI21X1 _18082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7848_),
    .B(_7855_),
    .C(_7816_),
    .Y(_7856_)
);

OAI21X1 _20687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf0),
    .B(_5668__bF$buf5),
    .C(_10365_),
    .Y(_10711_)
);

NAND2X1 _20267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9876_),
    .B(_9884_),
    .Y(_10251_)
);

NAND3X1 _16815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6443_),
    .B(_6458_),
    .C(_6465_),
    .Y(_6466_)
);

NOR2X1 _11950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2792_),
    .Y(_2803_)
);

NAND3X1 _19287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9168_),
    .B(_9169_),
    .C(_9171_),
    .Y(_9177_)
);

FILL SFILL23960x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11373_),
    .B(_11395_),
    .C(_11384_),
    .Y(_11406_)
);

NOR3X1 _12315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6758_),
    .C(_6714_),
    .Y(_6802_)
);

OAI21X1 _22833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .B(_1153_),
    .C(_1049_),
    .Y(_1154_)
);

OAI21X1 _22413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_694_),
    .C(_499_),
    .Y(_695_)
);

NOR2X1 _23618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1885_),
    .B(_1888_),
    .Y(_2009_)
);

NAND2X1 _17773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_27_bF$buf1),
    .Y(_7517_)
);

NAND3X1 _17353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7016_),
    .B(_7051_),
    .C(_7056_),
    .Y(_7057_)
);

NAND3X1 _18978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8836_),
    .B(_8837_),
    .C(_8835_),
    .Y(_8838_)
);

NAND3X1 _18558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8375_),
    .B(_8377_),
    .C(_8376_),
    .Y(_8378_)
);

NAND3X1 _18138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7900_),
    .B(_7907_),
    .C(_7886_),
    .Y(_7917_)
);

NAND2X1 _13693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3041_),
    .B(_3046_),
    .Y(_3047_)
);

OAI21X1 _13273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf3),
    .B(_2586__bF$buf0),
    .C(_2381_),
    .Y(_2587_)
);

NAND2X1 _23791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2194_),
    .B(_2195_),
    .Y(_2197_)
);

NOR3X1 _23371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1739_),
    .B(_1735_),
    .C(_1738_),
    .Y(_1741_)
);

XOR2X1 _14898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4068_),
    .B(_4364_),
    .Y(_4365_)
);

NAND3X1 _14478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3903_),
    .B(_3904_),
    .C(_3905_),
    .Y(_3906_)
);

NAND2X1 _14058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3444_),
    .B(_3445_),
    .Y(_3446_)
);

FILL SFILL64200x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_23_bF$buf1),
    .Y(_10502_)
);

AND2X2 _20076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10037_),
    .B(_10040_),
    .Y(_10041_)
);

OAI21X1 _16624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6256_),
    .B(_6251_),
    .C(_6221_),
    .Y(_6257_)
);

OAI22X1 _16204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5106_),
    .B(_5468_),
    .C(_5796_),
    .D(_5466_),
    .Y(_5797_)
);

NAND3X1 _19096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8959_),
    .B(_8964_),
    .C(_8966_),
    .Y(_8967_)
);

NAND2X1 _17829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7574_),
    .B(_7577_),
    .Y(_7578_)
);

OAI21X1 _17409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7117_),
    .B(_7113_),
    .C(_7108_),
    .Y(_7118_)
);

NAND2X1 _12964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(_1968_),
    .Y(_2001_)
);

OAI21X1 _12544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9203_),
    .B(_9214_),
    .C(_9038_),
    .Y(_9312_)
);

NOR2X1 _12124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3438_),
    .B(_3460_),
    .Y(_4708_)
);

INVX1 _22642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_944_),
    .Y(_945_)
);

NOR2X1 _22222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_236_),
    .Y(_485_)
);

OAI21X1 _13749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_10869__bF$buf1),
    .C(_3102_),
    .Y(_3108_)
);

OAI21X1 _13329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2641_),
    .B(_2642_),
    .C(_2636_),
    .Y(_2648_)
);

INVX2 _23847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2255_),
    .Y(_2256_)
);

XNOR2X1 _23427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .B(_1787_),
    .Y(_1801_)
);

OAI21X1 _23007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(_1337_),
    .C(_1216_),
    .Y(_1343_)
);

AOI21X1 _17582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6954_),
    .B(_6952_),
    .C(_7306_),
    .Y(_7307_)
);

OAI21X1 _17162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6846_),
    .B(_6441_),
    .C(_6482_),
    .Y(_6847_)
);

FILL SFILL33800x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8622_),
    .B(_8623_),
    .C(_8627_),
    .Y(_8628_)
);

NAND2X1 _18367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8120_),
    .B(_8116_),
    .Y(_8168_)
);

AOI21X1 _13082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1565_),
    .B(_1631_),
    .C(_1772_),
    .Y(_2378_)
);

NAND2X1 _23180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1394_),
    .Y(_1532_)
);

FILL SFILL8680x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11814_),
    .Y(_147_)
);

NAND3X1 _14287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3693_),
    .B(_3692_),
    .C(_3677_),
    .Y(_3697_)
);

FILL SFILL74280x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6504_),
    .B(_6507_),
    .C(_6506_),
    .Y(_6508_)
);

OAI21X1 _16433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6006_),
    .B(_6046_),
    .C(_5996_),
    .Y(_6047_)
);

NAND2X1 _16013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5586_),
    .B(_5587_),
    .Y(_5588_)
);

NAND3X1 _17638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7362_),
    .B(_7364_),
    .C(_7363_),
    .Y(_7368_)
);

NAND3X1 _17218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6902_),
    .B(_6907_),
    .C(_6906_),
    .Y(_6908_)
);

FILL SFILL69000x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10090_),
    .B(_10221_),
    .C(_10123_),
    .Y(_11822_)
);

INVX8 _12353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .Y(_7217_)
);

NOR2X1 _22871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1194_),
    .B(_1193_),
    .Y(_1196_)
);

OAI21X1 _22451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_520_),
    .B(_507_),
    .C(_528_),
    .Y(_736_)
);

AOI21X1 _22031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_274_),
    .C(_258_),
    .Y(_276_)
);

OAI21X1 _13978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3127_),
    .B(_3186_),
    .C(_3179_),
    .Y(_3358_)
);

AOI21X1 _13558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2889_),
    .B(_2886_),
    .C(_2877_),
    .Y(_2898_)
);

INVX1 _13138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .Y(_2439_)
);

NOR2X1 _23656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .B(_1994_),
    .Y(_2051_)
);

NAND2X1 _23236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1590_),
    .Y(_1593_)
);

FILL SFILL64200x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _17391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7096_),
    .B(_7097_),
    .Y(_7099_)
);

NAND3X1 _15704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5242_),
    .B(_5248_),
    .C(_5101_),
    .Y(_5249_)
);

NAND3X1 _18596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8411_),
    .B(_8412_),
    .C(_8281_),
    .Y(_8419_)
);

INVX1 _18176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7958_),
    .Y(_7959_)
);

FILL SFILL33720x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6245_),
    .B(_6568_),
    .C(_6567_),
    .Y(_6569_)
);

NAND3X1 _21722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11842_),
    .B(_11602_),
    .C(_11841_),
    .Y(_11846_)
);

OAI22X1 _21302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10818_),
    .B(_11135_),
    .C(_11385_),
    .D(_11134_),
    .Y(_11386_)
);

OAI21X1 _14096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3484_),
    .B(_3485_),
    .C(_3245_),
    .Y(_3488_)
);

NAND2X1 _12829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_13_bF$buf1),
    .Y(_527_)
);

XNOR2X1 _12409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7624_),
    .B(_7569_),
    .Y(_7832_)
);

NAND2X1 _22927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1255_),
    .B(_1254_),
    .Y(_1256_)
);

NAND2X1 _22507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_794_),
    .Y(_797_)
);

OR2X2 _16662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6296_),
    .B(_6298_),
    .Y(_6299_)
);

NAND2X1 _16242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .B(_5491_),
    .Y(_5839_)
);

OAI21X1 _17867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .B(_7615_),
    .C(_7223_),
    .Y(_7619_)
);

OAI21X1 _17447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7152_),
    .B(_7154_),
    .C(_7064_),
    .Y(_7160_)
);

NAND2X1 _17027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6697_),
    .B(_6698_),
    .Y(_6699_)
);

OAI21X1 _12582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9674_),
    .B(_9685_),
    .C(_8500_),
    .Y(_9729_)
);

INVX2 _12162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5113_),
    .Y(_5124_)
);

OAI21X1 _22680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf3),
    .B(_5676_),
    .C(_985_),
    .Y(_986_)
);

OAI21X1 _22260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_523_),
    .B(_522_),
    .C(_521_),
    .Y(_526_)
);

FILL SFILL8680x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3141_),
    .Y(_3150_)
);

AOI21X1 _13367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2675_),
    .B(_2678_),
    .C(_2659_),
    .Y(_2690_)
);

BUFX2 _23885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[3]),
    .Y(y[3])
);

AOI21X1 _23465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1829_),
    .B(_1833_),
    .C(_1779_),
    .Y(_1843_)
);

OAI21X1 _23045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_1384_),
    .C(_1267_),
    .Y(_1385_)
);

FILL SFILL74280x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .B(_5493_),
    .C(_5492_),
    .Y(_5500_)
);

AOI21X1 _15513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5037_),
    .B(_5038_),
    .C(_5035_),
    .Y(_5039_)
);

FILL SFILL34120x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6353_),
    .B(_6354_),
    .C(_6265_),
    .Y(_6360_)
);

NAND3X1 _21951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_185_),
    .C(_11829_),
    .Y(_189_)
);

AOI21X1 _21531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11635_),
    .B(_11632_),
    .C(_11607_),
    .Y(_11637_)
);

NAND3X1 _21111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11171_),
    .B(_11175_),
    .C(_11174_),
    .Y(_11177_)
);

FILL SFILL64280x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10035_),
    .B(_10178_),
    .C(_10244_),
    .Y(_10342_)
);

NOR3X1 _12218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5409_),
    .B(_5343_),
    .C(_5640_),
    .Y(_5738_)
);

XNOR2X1 _22736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1047_),
    .B(_1044_),
    .Y(_1048_)
);

AOI21X1 _22316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(_334_),
    .C(_587_),
    .Y(_588_)
);

FILL SFILL33800x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_17_bF$buf0),
    .Y(_6550_)
);

OAI21X1 _16471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5752_),
    .B(_6086_),
    .C(_5776_),
    .Y(_6089_)
);

NAND2X1 _16051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5627_),
    .B(_5628_),
    .Y(_5630_)
);

OAI21X1 _17676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7396_),
    .B(_7397_),
    .C(_7394_),
    .Y(_7410_)
);

NAND3X1 _17256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6947_),
    .B(_6948_),
    .C(_6949_),
    .Y(_6950_)
);

XNOR2X1 _12391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7624_),
    .B(_7580_),
    .Y(_7635_)
);

NAND2X1 _20802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf4),
    .B(areg_22_bF$buf1),
    .Y(_10838_)
);

FILL SFILL54200x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2790_),
    .B(_2934_),
    .C(_2940_),
    .Y(_2941_)
);

AOI21X1 _13176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2298_),
    .C(_2302_),
    .Y(_2481_)
);

INVX1 _23694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .Y(_2092_)
);

OAI21X1 _23274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1634_),
    .C(_1551_),
    .Y(_1635_)
);

XNOR2X1 _19822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9763_),
    .B(_9758_),
    .Y(_9764_)
);

OAI21X1 _19402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9302_),
    .B(_9297_),
    .C(_9283_),
    .Y(_9303_)
);

DFFPOSX1 _24059_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[17]),
    .CLK(clk_bF$buf5),
    .D(b[17])
);

OAI21X1 _15742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5288_),
    .B(_5290_),
    .C(_5285_),
    .Y(_5291_)
);

AND2X2 _15322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_20_bF$buf1),
    .Y(_4831_)
);

NAND2X1 _20399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf0),
    .B(breg_26_bF$buf3),
    .Y(_10395_)
);

NAND2X1 _16947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_18_bF$buf0),
    .Y(_6611_)
);

OAI21X1 _16527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .B(_6149_),
    .C(_6137_),
    .Y(_6150_)
);

NAND3X1 _16107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5684_),
    .B(_5689_),
    .C(_5687_),
    .Y(_5690_)
);

INVX2 _21760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11885_),
    .Y(_11886_)
);

AOI21X1 _21340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11421_),
    .B(_11422_),
    .C(_11420_),
    .Y(_11427_)
);

FILL SFILL44120x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_845_),
    .C(_144_),
    .Y(_943_)
);

INVX2 _12447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6955_),
    .Y(_8249_)
);

NAND2X1 _22965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1296_),
    .B(_1297_),
    .Y(_1298_)
);

INVX8 _12027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .Y(_3646_)
);

NOR2X1 _22545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_657_),
    .B(_664_),
    .Y(_839_)
);

NAND2X1 _22125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_26_bF$buf2),
    .Y(_379_)
);

OAI21X1 _16280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5874_),
    .B(_5875_),
    .C(_5876_),
    .Y(_5880_)
);

FILL SFILL38920x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7199_),
    .B(_7200_),
    .C(_7198_),
    .Y(_7201_)
);

OAI21X1 _17065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6739_),
    .B(_6740_),
    .C(_6738_),
    .Y(_6741_)
);

FILL SFILL3560x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10627_),
    .B(_10626_),
    .C(_10625_),
    .Y(_10629_)
);

XNOR2X1 _23083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(_1414_),
    .Y(_1426_)
);

NOR3X1 _19631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9549_),
    .B(_9173_),
    .C(_9553_),
    .Y(_9555_)
);

NOR3X1 _19211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9082_),
    .B(_9078_),
    .C(_9083_),
    .Y(_9093_)
);

NAND2X1 _21816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf2),
    .B(breg_22_bF$buf3),
    .Y(_40_)
);

OAI21X1 _15971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5540_),
    .B(_5213_),
    .C(_5206_),
    .Y(_5542_)
);

NAND3X1 _15551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5037_),
    .B(_5035_),
    .C(_5038_),
    .Y(_5081_)
);

AOI21X1 _15131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4616_),
    .B(_4615_),
    .C(_4614_),
    .Y(_4622_)
);

FILL SFILL28840x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6391_),
    .B(_6384_),
    .C(_6047_),
    .Y(_6402_)
);

AOI21X1 _16336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .B(_5561_),
    .C(_5565_),
    .Y(_5942_)
);

FILL SFILL18840x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10737_),
    .B(_10748_),
    .Y(_10759_)
);

OAI21X1 _12256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5453__bF$buf1),
    .C(_5442_),
    .Y(_6154_)
);

INVX1 _22774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1084_),
    .Y(_1090_)
);

OAI21X1 _22354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(_625_),
    .C(_619_),
    .Y(_630_)
);

OAI22X1 _18902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8368_),
    .B(_8369_),
    .C(_8372_),
    .D(_8362_),
    .Y(_8755_)
);

DFFPOSX1 _23979_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[33]),
    .CLK(clk_bF$buf3),
    .D(_0_[33])
);

OAI21X1 _23559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1941_),
    .B(_1940_),
    .C(_1939_),
    .Y(_1945_)
);

AOI21X1 _23139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(_1476_),
    .C(_1436_),
    .Y(_1487_)
);

AOI21X1 _14822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3993_),
    .B(_3995_),
    .C(_4282_),
    .Y(_4283_)
);

AOI21X1 _14402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3594_),
    .B(_3822_),
    .C(_3820_),
    .Y(_3823_)
);

NAND3X1 _17294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6969_),
    .B(_6982_),
    .C(_6973_),
    .Y(_6992_)
);

FILL SFILL44200x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5141_),
    .B(_5137_),
    .C(_5104_),
    .Y(_5142_)
);

AOI21X1 _20840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10860_),
    .B(_10864_),
    .C(_10867_),
    .Y(_10879_)
);

INVX1 _20420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10394_),
    .Y(_10418_)
);

NAND3X1 _20000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9938_),
    .B(_9945_),
    .C(_9754_),
    .Y(_9958_)
);

OAI21X1 _18499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8296_),
    .B(_8300_),
    .C(_8302_),
    .Y(_8313_)
);

AOI21X1 _18079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7827_),
    .B(_7830_),
    .C(_7840_),
    .Y(_7852_)
);

OAI21X1 _19860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_5921__bF$buf2),
    .C(_9446_),
    .Y(_9805_)
);

NAND3X1 _19440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9340_),
    .B(_9328_),
    .C(_9332_),
    .Y(_9344_)
);

INVX2 _19020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8882_),
    .Y(_8883_)
);

NOR2X1 _11947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2573_),
    .B(_2759_),
    .Y(_2770_)
);

AOI21X1 _21625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11738_),
    .B(_11737_),
    .C(_11736_),
    .Y(_11739_)
);

NAND3X1 _21205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11272_),
    .B(_11273_),
    .C(_11269_),
    .Y(_11280_)
);

NAND3X1 _15780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4974_),
    .B(_5325_),
    .C(_5330_),
    .Y(_5331_)
);

INVX2 _15360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4848_),
    .Y(_4872_)
);

FILL SFILL38920x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6266_),
    .B(_6651_),
    .C(_6273_),
    .Y(_6652_)
);

NAND3X1 _16565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6162_),
    .B(_6186_),
    .C(_6191_),
    .Y(_6192_)
);

NAND3X1 _16145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5731_),
    .B(_5725_),
    .C(_5730_),
    .Y(_5732_)
);

FILL SFILL69240x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8654_),
    .Y(_8665_)
);

NAND3X1 _12065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3799_),
    .B(_3493_),
    .C(_3832_),
    .Y(_4061_)
);

OAI21X1 _22583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_833_),
    .B(_838_),
    .C(_880_),
    .Y(_881_)
);

NOR3X1 _22163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(_417_),
    .C(_419_),
    .Y(_421_)
);

NAND3X1 _18711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8536_),
    .B(_8540_),
    .C(_8543_),
    .Y(_8545_)
);

NAND2X1 _23788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2192_),
    .Y(_2193_)
);

AOI21X1 _23368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_1732_),
    .C(_1736_),
    .Y(_1737_)
);

NAND2X1 _19916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9865_),
    .B(_9866_),
    .Y(_9867_)
);

AOI21X1 _14631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3794_),
    .B(_3796_),
    .C(_3791_),
    .Y(_4073_)
);

NAND3X1 _14211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3607_),
    .B(_3609_),
    .C(_3608_),
    .Y(_3614_)
);

FILL SFILL18920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5388_),
    .B(_5392_),
    .C(_5379_),
    .Y(_5393_)
);

OAI21X1 _15416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4930_),
    .C(_4676_),
    .Y(_4934_)
);

FILL SFILL18840x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_81_),
    .C(_75_),
    .Y(_82_)
);

XNOR2X1 _21434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11530_),
    .B(_11526_),
    .Y(_11531_)
);

OAI21X1 _21014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf2),
    .B(_5315__bF$buf1),
    .C(_11062_),
    .Y(_11070_)
);

FILL SFILL38920x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13960x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_934_),
    .C(_940_),
    .Y(_941_)
);

NAND3X1 _22219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_480_),
    .B(_481_),
    .C(_479_),
    .Y(_482_)
);

NOR2X1 _13902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3275_),
    .B(_3268_),
    .Y(_3276_)
);

OAI21X1 _16794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5685_),
    .B(_6442_),
    .C(_6066_),
    .Y(_6443_)
);

NOR3X1 _16374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5595_),
    .B(_5597_),
    .C(_5594_),
    .Y(_5983_)
);

NAND3X1 _17999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7761_),
    .B(_7762_),
    .C(_7763_),
    .Y(_7764_)
);

AOI21X1 _17579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7297_),
    .B(_7298_),
    .C(_7296_),
    .Y(_7303_)
);

NAND3X1 _17159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6435_),
    .B(_6839_),
    .C(_6842_),
    .Y(_6843_)
);

NAND2X1 _12294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_9_bF$buf1),
    .Y(_6571_)
);

NAND3X1 _22392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_605_),
    .C(_606_),
    .Y(_671_)
);

NAND3X1 _18940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8734_),
    .B(_8736_),
    .C(_8729_),
    .Y(_8796_)
);

INVX1 _18520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8335_),
    .Y(_8336_)
);

NOR3X1 _18100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7856_),
    .B(_7864_),
    .C(_7866_),
    .Y(_7875_)
);

AOI21X1 _20705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10354_),
    .B(_10378_),
    .C(_10376_),
    .Y(_10731_)
);

FILL SFILL69240x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2794_),
    .B(_2833_),
    .C(_2828_),
    .Y(_2834_)
);

INVX2 _13079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .Y(_2374_)
);

OAI21X1 _23597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1972_),
    .B(_1981_),
    .C(_1985_),
    .Y(_1986_)
);

NOR3X1 _23177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1406_),
    .C(_1519_),
    .Y(_1529_)
);

NAND2X1 _19725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9655_),
    .B(_9656_),
    .Y(_9657_)
);

FILL SFILL38600x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9188_),
    .B(_9196_),
    .C(_9096_),
    .Y(_9197_)
);

AOI21X1 _14860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4309_),
    .B(_4315_),
    .C(_4063_),
    .Y(_4324_)
);

NAND3X1 _14440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3861_),
    .B(_3863_),
    .C(_3862_),
    .Y(_3864_)
);

OAI21X1 _14020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_3402__bF$buf1),
    .C(_3403_),
    .Y(_3404_)
);

FILL SFILL3640x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48760x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_22_bF$buf1),
    .Y(_5184_)
);

AND2X2 _15225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4450_),
    .B(_4451_),
    .Y(_4724_)
);

AOI21X1 _11985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .B(_3176_),
    .C(_3143_),
    .Y(_3187_)
);

INVX2 _21663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11755_),
    .Y(_11781_)
);

AOI21X1 _21243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11280_),
    .B(_11283_),
    .C(_11014_),
    .Y(_11321_)
);

FILL SFILL28920x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf4),
    .B(areg_28_bF$buf2),
    .Y(_1192_)
);

AND2X2 _22448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_592_),
    .B(_585_),
    .Y(_732_)
);

AOI21X1 _22028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11897_),
    .B(_11903_),
    .C(_11906_),
    .Y(_272_)
);

NAND2X1 _13711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3061_),
    .B(_3065_),
    .Y(_3067_)
);

AOI21X1 _16183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5765_),
    .B(_5773_),
    .C(_5752_),
    .Y(_5774_)
);

FILL SFILL39080x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4384_),
    .B(_4380_),
    .Y(_4385_)
);

INVX1 _17388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7094_),
    .Y(_7095_)
);

FILL SFILL18760x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10982_),
    .B(_10978_),
    .C(_10692_),
    .Y(_10983_)
);

NAND3X1 _20514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10499_),
    .B(_10514_),
    .C(_10521_),
    .Y(_10522_)
);

OAI21X1 _19954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9906_),
    .B(_9907_),
    .C(_9903_),
    .Y(_9908_)
);

OAI22X1 _19534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8699_),
    .B(_9446_),
    .C(_9447_),
    .D(_9098_),
    .Y(_9448_)
);

OAI21X1 _19114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8981_),
    .B(_8982_),
    .C(_8934_),
    .Y(_8987_)
);

OAI21X1 _21719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11830_),
    .B(_11827_),
    .C(_11715_),
    .Y(_11842_)
);

FILL SFILL8760x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5433_),
    .B(_5434_),
    .C(_5432_),
    .Y(_5435_)
);

NOR2X1 _15454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4658_),
    .B(_4973_),
    .Y(_4974_)
);

NAND3X1 _15034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4514_),
    .B(_4507_),
    .C(_4512_),
    .Y(_4515_)
);

FILL SFILL53960x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53880x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6294_),
    .Y(_6295_)
);

NAND2X1 _16239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5834_),
    .B(_5830_),
    .Y(_5835_)
);

OAI21X1 _21892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_114_),
    .C(_116_),
    .Y(_124_)
);

AOI21X1 _21472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11010_),
    .B(_11288_),
    .C(_11572_),
    .Y(_11573_)
);

NAND2X1 _21052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11056_),
    .B(_11052_),
    .Y(_11112_)
);

AOI21X1 _17600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6997_),
    .B(_7002_),
    .C(_7003_),
    .Y(_7326_)
);

NAND2X1 _12999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_14_bF$buf4),
    .Y(_2294_)
);

OAI21X1 _12579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9674_),
    .B(_9685_),
    .C(_9663_),
    .Y(_9696_)
);

XNOR2X1 _12159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5080_),
    .B(_5025_),
    .Y(_5091_)
);

OAI21X1 _22677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf3),
    .B(_5315__bF$buf2),
    .C(_777_),
    .Y(_983_)
);

NOR3X1 _22257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .B(_511_),
    .C(_513_),
    .Y(_523_)
);

FILL SFILL3720x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_3402__bF$buf0),
    .C(_8637_),
    .Y(_8648_)
);

AND2X2 _13940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3314_),
    .B(_3315_),
    .Y(_3317_)
);

INVX1 _13520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2844_),
    .Y(_2857_)
);

NAND2X1 _13100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2396_),
    .Y(_2397_)
);

FILL SFILL3640x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .B(_3884_),
    .C(_3890_),
    .Y(_4176_)
);

NAND3X1 _14305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3711_),
    .B(_3710_),
    .C(_3713_),
    .Y(_3717_)
);

NOR3X1 _17197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6529_),
    .B(_6531_),
    .C(_6525_),
    .Y(_6885_)
);

FILL SFILL49080x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10468_),
    .B(_10772_),
    .C(_10492_),
    .Y(_10773_)
);

AOI21X1 _20323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9640_),
    .B(_9963_),
    .C(_10312_),
    .Y(_10313_)
);

OR2X2 _19763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9692_),
    .B(_9693_),
    .Y(_9699_)
);

NOR3X1 _19343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8839_),
    .B(_8845_),
    .C(_8848_),
    .Y(_9239_)
);

FILL SFILL33880x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_182_),
    .C(_184_),
    .Y(_185_)
);

OAI21X1 _21528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11629_),
    .B(_11630_),
    .C(_11626_),
    .Y(_11633_)
);

AND2X2 _21108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf3),
    .B(areg_26_bF$buf4),
    .Y(_11173_)
);

OAI21X1 _15683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5220_),
    .B(_5221_),
    .C(_5181_),
    .Y(_5225_)
);

NAND2X1 _15263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4765_),
    .B(_4759_),
    .Y(_4766_)
);

FILL SFILL18600x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6190_),
    .B(_6188_),
    .C(_6180_),
    .Y(_6546_)
);

OAI21X1 _16468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .B(_6075_),
    .C(_6072_),
    .Y(_6084_)
);

NAND3X1 _16048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5366_),
    .B(_5621_),
    .C(_5625_),
    .Y(_5626_)
);

NOR3X1 _21281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11358_),
    .B(_11359_),
    .C(_11360_),
    .Y(_11363_)
);

FILL SFILL23880x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL63960x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6385_),
    .B(_7591_),
    .Y(_7602_)
);

OAI21X1 _22486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_554_),
    .B(_561_),
    .C(_550_),
    .Y(_774_)
);

AOI21X1 _22066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_309_),
    .B(_307_),
    .C(_306_),
    .Y(_314_)
);

AOI21X1 _18614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8028_),
    .B(_8031_),
    .C(_8438_),
    .Y(_8439_)
);

FILL SFILL8760x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9702_),
    .B(_9759_),
    .Y(_9760_)
);

NAND3X1 _14954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4419_),
    .B(_4426_),
    .C(_4388_),
    .Y(_4427_)
);

AOI21X1 _14534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3967_),
    .B(_3966_),
    .C(_3965_),
    .Y(_3968_)
);

AOI22X1 _14114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11582_),
    .B(_11625_),
    .C(_3506_),
    .D(_3505_),
    .Y(_3507_)
);

FILL SFILL29000x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5264_),
    .B(_5272_),
    .C(_5269_),
    .Y(_5287_)
);

OAI21X1 _15319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_3146__bF$buf0),
    .C(_4820_),
    .Y(_4827_)
);

INVX2 _20972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11023_),
    .Y(_11024_)
);

INVX2 _20552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10563_),
    .Y(_10564_)
);

NAND3X1 _20132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10097_),
    .B(_9999_),
    .C(_10102_),
    .Y(_10103_)
);

NAND2X1 _19992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9949_),
    .B(_9947_),
    .Y(_9950_)
);

NAND2X1 _19572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf2),
    .B(areg_25_bF$buf4),
    .Y(_9490_)
);

AOI21X1 _19152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8609_),
    .B(_8618_),
    .C(_8625_),
    .Y(_9029_)
);

AOI21X1 _21757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11842_),
    .B(_11841_),
    .C(_11602_),
    .Y(_11883_)
);

FILL SFILL3720x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11205_),
    .B(_11210_),
    .C(_11217_),
    .Y(_11424_)
);

FILL SFILL43960x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7109_),
    .B(_8359_),
    .C(_9915_),
    .Y(_9926_)
);

NOR2X1 _15492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5013_),
    .B(_5015_),
    .Y(_5016_)
);

OAI21X1 _15072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4554_),
    .B(_4556_),
    .C(_4550_),
    .Y(_4557_)
);

OAI21X1 _13805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3164_),
    .B(_3169_),
    .C(_3128_),
    .Y(_3170_)
);

BUFX2 _23903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[21]),
    .Y(y[21])
);

AOI21X1 _16697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5928_),
    .B(_5948_),
    .C(_6336_),
    .Y(_6337_)
);

NOR3X1 _16277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5874_),
    .B(_5875_),
    .C(_5876_),
    .Y(_5877_)
);

NAND3X1 _21090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11147_),
    .B(_11149_),
    .C(_11148_),
    .Y(_11153_)
);

FILL SFILL64360x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5497_),
    .B(_5486_),
    .Y(_5508_)
);

AOI21X1 _22295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_550_),
    .C(_545_),
    .Y(_565_)
);

NOR3X1 _18843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8674_),
    .B(_8679_),
    .C(_8680_),
    .Y(_8690_)
);

NAND2X1 _18423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8224_),
    .B(_8229_),
    .Y(_8230_)
);

AOI21X1 _18003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7762_),
    .B(_7763_),
    .C(_7761_),
    .Y(_7769_)
);

FILL SFILL33880x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10624_),
    .B(_10623_),
    .Y(_10625_)
);

NAND3X1 _19628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9530_),
    .B(_9544_),
    .C(_9539_),
    .Y(_9551_)
);

NAND3X1 _19208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9006_),
    .B(_9088_),
    .C(_9084_),
    .Y(_9089_)
);

INVX1 _14763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3949_),
    .Y(_4218_)
);

AOI21X1 _14343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3746_),
    .B(_3747_),
    .C(_3522_),
    .Y(_3759_)
);

DFFPOSX1 _24021_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[11]),
    .CLK(clk_bF$buf1),
    .D(a[11])
);

NAND3X1 _15968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5536_),
    .B(_5535_),
    .C(_5537_),
    .Y(_5538_)
);

AOI21X1 _15548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5059_),
    .B(_5065_),
    .C(_5043_),
    .Y(_5077_)
);

NAND3X1 _15128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4613_),
    .B(_4617_),
    .C(_4352_),
    .Y(_4618_)
);

NAND2X1 _20781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10527_),
    .B(_10535_),
    .Y(_10815_)
);

FILL SFILL23880x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf3),
    .B(_6815__bF$buf2),
    .Y(_10354_)
);

FILL SFILL54280x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _19381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9278_),
    .Y(_9280_)
);

OAI21X1 _21986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_217_),
    .C(_220_),
    .Y(_227_)
);

FILL SFILL23800x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11665_),
    .B(_11666_),
    .C(_11663_),
    .Y(_11674_)
);

AOI21X1 _21146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11204_),
    .B(_11197_),
    .C(_11167_),
    .Y(_11215_)
);

FILL SFILL8840x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2954_),
    .B(_2955_),
    .C(_2756_),
    .Y(_2961_)
);

OAI21X1 _23712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(_1654_),
    .C(_1767_),
    .Y(_2111_)
);

OAI21X1 _16086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5632_),
    .B(_5630_),
    .C(_5621_),
    .Y(_5667_)
);

FILL SFILL13800x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4276_),
    .B(_4278_),
    .C(_4277_),
    .Y(_4279_)
);

FILL SFILL74040x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19080x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8479_),
    .Y(_8480_)
);

NOR3X1 _18232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7586_),
    .B(_7587_),
    .C(_7585_),
    .Y(_8020_)
);

NAND3X1 _20837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10852_),
    .B(_10868_),
    .C(_10875_),
    .Y(_10876_)
);

AOI21X1 _20417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10113_),
    .B(_10414_),
    .C(_10413_),
    .Y(_10415_)
);

FILL SFILL43960x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_4551__bF$buf0),
    .C(_9792_),
    .Y(_9802_)
);

OAI21X1 _19437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9338_),
    .B(_9337_),
    .C(_9340_),
    .Y(_9341_)
);

AOI21X1 _19017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8861_),
    .B(_8862_),
    .C(_8477_),
    .Y(_8880_)
);

FILL SFILL64440x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4462_),
    .B(_4454_),
    .C(_4467_),
    .Y(_4468_)
);

OAI21X1 _14572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3990_),
    .B(_3996_),
    .C(_4000_),
    .Y(_4010_)
);

OAI21X1 _14152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3548_),
    .B(_3546_),
    .C(_3540_),
    .Y(_3549_)
);

OAI21X1 _15777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_3781__bF$buf3),
    .C(_4679_),
    .Y(_5328_)
);

AOI21X1 _15357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4860_),
    .B(_4858_),
    .C(_4856_),
    .Y(_4869_)
);

NAND3X1 _20590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10596_),
    .B(_10594_),
    .C(_10590_),
    .Y(_10605_)
);

OAI21X1 _20170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9816_),
    .B(_10143_),
    .C(_9800_),
    .Y(_10144_)
);

OAI21X1 _19190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9064_),
    .B(_9069_),
    .C(_9040_),
    .Y(_9070_)
);

NOR3X1 _21795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_11894_),
    .C(_8_),
    .Y(_17_)
);

INVX2 _21375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11441_),
    .Y(_11466_)
);

NOR2X1 _17923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7243_),
    .B(_7680_),
    .Y(_7681_)
);

OAI21X1 _17503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7200_),
    .B(_7198_),
    .C(_7191_),
    .Y(_7220_)
);

NAND2X1 _18708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_22_bF$buf0),
    .Y(_8541_)
);

OAI21X1 _13843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3204_),
    .B(_3211_),
    .C(_2987_),
    .Y(_3212_)
);

OAI21X1 _13423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .B(_2750_),
    .C(_2744_),
    .Y(_2751_)
);

BUFX2 _23941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[59]),
    .Y(y[59])
);

OAI21X1 _13003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2296_),
    .B(_2297_),
    .C(_2238_),
    .Y(_2298_)
);

NAND2X1 _23521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_26_bF$buf1),
    .B(areg_29_bF$buf5),
    .Y(_1903_)
);

OAI21X1 _23101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300__bF$buf2),
    .B(_5676_),
    .C(_1444_),
    .Y(_1446_)
);

INVX2 _14628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf3),
    .Y(_4069_)
);

OAI21X1 _14208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_9104__bF$buf0),
    .C(_3331_),
    .Y(_3609_)
);

NAND3X1 _18881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8714_),
    .B(_8722_),
    .C(_8701_),
    .Y(_8732_)
);

OAI21X1 _18461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7923_),
    .B(_7922_),
    .C(_7919_),
    .Y(_8272_)
);

NAND3X1 _18041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7809_),
    .B(_7806_),
    .C(_7791_),
    .Y(_7811_)
);

FILL SFILL8920x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9252_),
    .B(_9253_),
    .C(_9251_),
    .Y(_10666_)
);

NAND2X1 _20226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9918_),
    .B(_9919_),
    .Y(_10206_)
);

NAND3X1 _19666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .B(_9384_),
    .C(_9385_),
    .Y(_9593_)
);

NAND3X1 _19246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9122_),
    .B(_9118_),
    .C(_9102_),
    .Y(_9132_)
);

NAND2X1 _14381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .B(_3797_),
    .Y(_3800_)
);

FILL SFILL69560x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74520x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5112_),
    .B(_5114_),
    .Y(_5119_)
);

INVX1 _15166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4658_),
    .Y(_4659_)
);

FILL SFILL74120x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38680x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11252_),
    .Y(_11257_)
);

NAND3X1 _17732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7471_),
    .B(_7464_),
    .C(_7469_),
    .Y(_7472_)
);

OAI21X1 _17312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7005_),
    .B(_7006_),
    .C(_7003_),
    .Y(_7011_)
);

FILL SFILL49000x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _22389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_667_),
    .Y(_668_)
);

NAND2X1 _18937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8791_),
    .B(_8792_),
    .Y(_8793_)
);

NAND2X1 _18517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_26_bF$buf3),
    .Y(_8333_)
);

NOR2X1 _13652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2797_),
    .B(_3001_),
    .Y(_3002_)
);

AND2X2 _13232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2533_),
    .B(_2532_),
    .Y(_2542_)
);

XNOR2X1 _23750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2151_),
    .B(_2126_),
    .Y(_2152_)
);

NAND3X1 _23330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .B(_1588_),
    .C(_1581_),
    .Y(_1695_)
);

FILL SFILL64040x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4320_),
    .C(_4059_),
    .Y(_4321_)
);

AND2X2 _14437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3572_),
    .B(_3566_),
    .Y(_3861_)
);

NAND2X1 _14017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3399_),
    .B(_3400_),
    .Y(_3401_)
);

FILL SFILL38920x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8518_),
    .B(_8517_),
    .C(_8516_),
    .Y(_8521_)
);

NOR3X1 _18270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8039_),
    .B(_8044_),
    .C(_8047_),
    .Y(_8062_)
);

INVX1 _20875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10917_),
    .Y(_10918_)
);

NAND3X1 _20455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10447_),
    .B(_10453_),
    .C(_10443_),
    .Y(_10457_)
);

NAND2X1 _20035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9743_),
    .B(_9748_),
    .Y(_9996_)
);

FILL SFILL18680x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9822_),
    .B(_9790_),
    .C(_9829_),
    .Y(_9844_)
);

AND2X2 _19475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8985_),
    .B(_8979_),
    .Y(_9383_)
);

NAND3X1 _19055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8896_),
    .B(_8920_),
    .C(_8921_),
    .Y(_8922_)
);

NAND2X1 _14190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3589_),
    .B(_3584_),
    .Y(_3590_)
);

FILL SFILL19000x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11756_),
    .B(_11778_),
    .C(_1543_),
    .Y(_1554_)
);

NAND2X1 _12503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8786_),
    .B(_8830_),
    .Y(_8863_)
);

NAND3X1 _22601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_895_),
    .C(_896_),
    .Y(_901_)
);

NAND3X1 _15395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4885_),
    .B(_4891_),
    .C(_4894_),
    .Y(_4911_)
);

NOR2X1 _13708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .B(_3062_),
    .Y(_3063_)
);

INVX1 _23806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2211_),
    .Y(_2212_)
);

BUFX2 BUFX2_insert200 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520_),
    .Y(_7520__bF$buf3)
);

BUFX2 BUFX2_insert201 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520_),
    .Y(_7520__bF$buf2)
);

BUFX2 BUFX2_insert202 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520_),
    .Y(_7520__bF$buf1)
);

BUFX2 BUFX2_insert203 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520_),
    .Y(_7520__bF$buf0)
);

OAI22X1 _17961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6927_),
    .B(_7721_),
    .C(_7373_),
    .D(_7348_),
    .Y(_7723_)
);

BUFX2 BUFX2_insert204 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100_),
    .Y(_7100__bF$buf3)
);

AOI21X1 _17541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6816_),
    .B(_7260_),
    .C(_6832_),
    .Y(_7262_)
);

BUFX2 BUFX2_insert205 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100_),
    .Y(_7100__bF$buf2)
);

BUFX2 BUFX2_insert206 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100_),
    .Y(_7100__bF$buf1)
);

NAND2X1 _17121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6801_),
    .B(_6798_),
    .Y(_6803_)
);

BUFX2 BUFX2_insert207 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100_),
    .Y(_7100__bF$buf0)
);

BUFX2 BUFX2_insert208 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[26]),
    .Y(areg_26_bF$buf4)
);

BUFX2 BUFX2_insert209 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[26]),
    .Y(areg_26_bF$buf3)
);

NAND3X1 _22198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_457_),
    .C(_452_),
    .Y(_459_)
);

OAI21X1 _18746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8578_),
    .B(_8579_),
    .C(_8527_),
    .Y(_8583_)
);

NAND2X1 _18326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7724_),
    .B(_7730_),
    .Y(_8123_)
);

INVX8 _13881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .Y(_3253_)
);

OAI21X1 _13461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2707_),
    .B(_2791_),
    .C(_2698_),
    .Y(_2793_)
);

NAND3X1 _13041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .B(_2335_),
    .C(_1423_),
    .Y(_2336_)
);

FILL SFILL69160x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3869_),
    .B(_4110_),
    .C(_4109_),
    .Y(_4111_)
);

FILL SFILL74120x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3650_),
    .B(_3651_),
    .C(_3649_),
    .Y(_3652_)
);

FILL SFILL28920x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf5)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf4)
);

FILL SFILL8840x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[27]),
    .Y(areg_27_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf1)
);

AND2X2 _20684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_10708_)
);

AOI21X1 _20264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10229_),
    .B(_10237_),
    .C(_10214_),
    .Y(_10248_)
);

OAI21X1 _16812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf0),
    .B(_3781__bF$buf2),
    .C(_6070_),
    .Y(_6463_)
);

OAI21X1 _19284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf0),
    .B(_8759_),
    .C(_8772_),
    .Y(_9174_)
);

FILL SFILL28760x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_115_),
    .C(_102_),
    .Y(_120_)
);

AOI21X1 _21469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11567_),
    .B(_11568_),
    .C(_11323_),
    .Y(_11569_)
);

FILL SFILL64120x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11096_),
    .B(_11091_),
    .C(_11059_),
    .Y(_11108_)
);

INVX2 _12732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10002_),
    .Y(_11373_)
);

OAI21X1 _12312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6758_),
    .C(_6714_),
    .Y(_6769_)
);

XNOR2X1 _22830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1147_),
    .Y(_1150_)
);

NAND2X1 _22410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_689_),
    .B(_688_),
    .Y(_690_)
);

NAND2X1 _13937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_13_bF$buf0),
    .Y(_3314_)
);

AOI21X1 _13517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .B(_2853_),
    .C(_2656_),
    .Y(_2854_)
);

NOR2X1 _23615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(_2005_),
    .Y(_2006_)
);

FILL FILL74040x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7512_),
    .B(_7130_),
    .C(_7119_),
    .Y(_7513_)
);

AOI21X1 _17350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7038_),
    .B(_7042_),
    .C(_7023_),
    .Y(_7053_)
);

FILL SFILL54120x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8418_),
    .B(_8420_),
    .C(_8834_),
    .Y(_8835_)
);

INVX1 _18555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8361_),
    .Y(_8375_)
);

AOI21X1 _18135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7507_),
    .B(_7505_),
    .C(_7508_),
    .Y(_7914_)
);

NAND3X1 _13690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .B(_3029_),
    .C(_3039_),
    .Y(_3043_)
);

NAND2X1 _13270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_12_bF$buf3),
    .Y(_2583_)
);

AND2X2 _14895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4134_),
    .B(_4126_),
    .Y(_4362_)
);

NAND3X1 _14475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3897_),
    .B(_3899_),
    .C(_3896_),
    .Y(_3903_)
);

NAND3X1 _14055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3357_),
    .B(_3442_),
    .C(_3435_),
    .Y(_3443_)
);

OAI21X1 _20493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10143_),
    .B(_10498_),
    .C(_10152_),
    .Y(_10499_)
);

OAI21X1 _20073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10034_),
    .B(_10033_),
    .C(_10032_),
    .Y(_10038_)
);

AOI21X1 _16621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6238_),
    .B(_6243_),
    .C(_6225_),
    .Y(_6254_)
);

NAND3X1 _16201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5783_),
    .B(_5790_),
    .C(_5791_),
    .Y(_5794_)
);

NAND3X1 _19093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8960_),
    .B(_8962_),
    .C(_8963_),
    .Y(_8964_)
);

NAND2X1 _21698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11817_),
    .B(_11810_),
    .Y(_11819_)
);

AOI21X1 _21278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11019_),
    .B(_11042_),
    .C(_11040_),
    .Y(_11358_)
);

NAND3X1 _17826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7475_),
    .B(_7464_),
    .C(_7469_),
    .Y(_7575_)
);

NAND3X1 _17406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7110_),
    .B(_7114_),
    .C(_7112_),
    .Y(_7115_)
);

XNOR2X1 _12961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1957_),
    .B(_1925_),
    .Y(_1968_)
);

FILL SFILL69240x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9257_),
    .B(_9268_),
    .C(_9247_),
    .Y(_9279_)
);

AOI21X1 _12121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4533_),
    .B(_4577_),
    .C(_4237_),
    .Y(_4675_)
);

FILL SFILL38760x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_10869__bF$buf3),
    .C(_2849_),
    .Y(_3105_)
);

NAND3X1 _13326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2644_),
    .B(_2629_),
    .C(_2637_),
    .Y(_2645_)
);

XOR2X1 _23844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2245_),
    .B(_2252_),
    .Y(_2253_)
);

XNOR2X1 _23424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1797_),
    .B(_1793_),
    .Y(_1798_)
);

NAND3X1 _23004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1268_),
    .B(_1335_),
    .C(_1339_),
    .Y(_1340_)
);

FILL SFILL3800x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8211_),
    .B(_8624_),
    .Y(_8625_)
);

AOI21X1 _18364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8151_),
    .B(_8155_),
    .C(_8123_),
    .Y(_8165_)
);

INVX2 _20969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11019_),
    .Y(_11020_)
);

XNOR2X1 _20549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10559_),
    .B(_10557_),
    .Y(_10560_)
);

AOI21X1 _20129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10089_),
    .B(_10083_),
    .C(_10041_),
    .Y(_10099_)
);

AOI21X1 _21910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_137_),
    .B(_138_),
    .C(_136_),
    .Y(_143_)
);

AOI21X1 _19989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9938_),
    .B(_9945_),
    .C(_9754_),
    .Y(_9946_)
);

XOR2X1 _19569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9446_),
    .B(_9485_),
    .Y(_9486_)
);

NOR2X1 _19149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9018_),
    .B(_9019_),
    .Y(_9025_)
);

NAND3X1 _14284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3691_),
    .B(_3693_),
    .C(_3692_),
    .Y(_3694_)
);

NAND2X1 _15489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_21_bF$buf2),
    .Y(_5012_)
);

OAI21X1 _15069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_4541__bF$buf4),
    .C(_4245_),
    .Y(_4553_)
);

FILL SFILL18760x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6111_),
    .B(_6102_),
    .Y(_6504_)
);

OAI21X1 _16430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6019_),
    .B(_6017_),
    .C(_6010_),
    .Y(_6043_)
);

NAND3X1 _16010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5578_),
    .B(_5583_),
    .C(_5539_),
    .Y(_5584_)
);

AOI21X1 _21087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11149_),
    .B(_11148_),
    .C(_11147_),
    .Y(_11150_)
);

AOI21X1 _17635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7364_),
    .B(_7363_),
    .C(_7362_),
    .Y(_7365_)
);

NAND3X1 _17215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6888_),
    .B(_6893_),
    .C(_6897_),
    .Y(_6905_)
);

OAI21X1 _12770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10112_),
    .B(_11767_),
    .C(_11778_),
    .Y(_11789_)
);

NAND2X1 _12350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6055_),
    .B(_6087_),
    .Y(_7185_)
);

FILL SFILL23960x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3343_),
    .B(_3339_),
    .C(_3344_),
    .Y(_3355_)
);

INVX2 _13555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2871_),
    .Y(_2895_)
);

XOR2X1 _13135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1936_),
    .B(_2435_),
    .Y(_2436_)
);

XNOR2X1 _23653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_1997_),
    .Y(_2048_)
);

XOR2X1 _23233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1589_),
    .B(_1577_),
    .Y(_1590_)
);

FILL SFILL69320x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24018_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[8]),
    .CLK(clk_bF$buf5),
    .D(a[8])
);

AOI21X1 _15701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5240_),
    .B(_5239_),
    .C(_5238_),
    .Y(_5246_)
);

OAI21X1 _18593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8277_),
    .B(_8276_),
    .C(_8188_),
    .Y(_8416_)
);

AOI21X1 _18173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7540_),
    .B(_7535_),
    .C(_7528_),
    .Y(_7956_)
);

NAND2X1 _20778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10806_),
    .B(_10810_),
    .Y(_10811_)
);

NOR2X1 _20358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf2),
    .B(_7225__bF$buf3),
    .Y(_10350_)
);

AOI21X1 _16906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6555_),
    .B(_6554_),
    .C(_6551_),
    .Y(_6566_)
);

NAND2X1 _19798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9686_),
    .B(_9682_),
    .Y(_9737_)
);

OAI21X1 _19378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9275_),
    .B(_9002_),
    .C(_9223_),
    .Y(_9276_)
);

AOI21X1 _14093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3474_),
    .B(_3466_),
    .C(_3246_),
    .Y(_3485_)
);

INVX2 _12826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_484_),
    .Y(_494_)
);

AOI21X1 _12406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7722_),
    .B(_7700_),
    .C(_7678_),
    .Y(_7799_)
);

XNOR2X1 _22924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1095_),
    .B(_1253_),
    .Y(_0_[49])
);

OAI21X1 _22504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .B(_791_),
    .C(_793_),
    .Y(_794_)
);

AOI21X1 _15298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4499_),
    .B(_4520_),
    .C(_4523_),
    .Y(_4804_)
);

FILL SFILL3800x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _23709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1542_),
    .B(_2106_),
    .C(_1400_),
    .Y(_2107_)
);

FILL SFILL59240x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49320x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .B(_7615_),
    .C(_7613_),
    .Y(_7616_)
);

NAND3X1 _17444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7058_),
    .B(_7051_),
    .C(_7056_),
    .Y(_7157_)
);

INVX2 _17024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .Y(_6696_)
);

AOI21X1 _18649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8440_),
    .B(_8441_),
    .C(_8078_),
    .Y(_8476_)
);

OAI21X1 _18229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7998_),
    .B(_8004_),
    .C(_8007_),
    .Y(_8017_)
);

AND2X2 _13784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_17_bF$buf2),
    .Y(_3147_)
);

FILL FILL74200x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _23882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[0]),
    .Y(y[0])
);

OAI21X1 _13364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2676_),
    .C(_2662_),
    .Y(_2687_)
);

OAI21X1 _23462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1837_),
    .B(_1839_),
    .C(_1733_),
    .Y(_1840_)
);

NAND3X1 _23042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1377_),
    .C(_1376_),
    .Y(_1382_)
);

NOR2X1 _14989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4460_),
    .B(_4463_),
    .Y(_4464_)
);

NAND3X1 _14569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3902_),
    .B(_3906_),
    .C(_3908_),
    .Y(_4006_)
);

NAND3X1 _14149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3541_),
    .B(_3544_),
    .C(_3543_),
    .Y(_3545_)
);

FILL SFILL18760x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5160_),
    .B(_5163_),
    .C(_5165_),
    .Y(_5496_)
);

XNOR2X1 _15510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5016_),
    .B(_5010_),
    .Y(_5035_)
);

OAI21X1 _20587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10601_),
    .B(_10597_),
    .C(_10270_),
    .Y(_10602_)
);

NOR2X1 _20167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10136_),
    .B(_10140_),
    .Y(_10141_)
);

NAND3X1 _16715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6221_),
    .B(_6259_),
    .C(_6260_),
    .Y(_6357_)
);

NAND3X1 _19187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9048_),
    .B(_9052_),
    .C(_9062_),
    .Y(_9067_)
);

FILL SFILL23960x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8731_),
    .B(_8852_),
    .C(_8917_),
    .Y(_10310_)
);

AOI21X1 _12215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5694_),
    .B(_5651_),
    .C(_4992_),
    .Y(_5705_)
);

NAND2X1 _22733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_30_bF$buf4),
    .Y(_1045_)
);

NAND3X1 _22313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_579_),
    .C(_584_),
    .Y(_585_)
);

FILL SFILL69320x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _23938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[56]),
    .Y(y[56])
);

NAND2X1 _23518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1808_),
    .B(_1817_),
    .Y(_1899_)
);

NAND3X1 _17673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7401_),
    .B(_7406_),
    .C(_7379_),
    .Y(_7407_)
);

AOI21X1 _17253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6519_),
    .B(_6528_),
    .C(_6534_),
    .Y(_6947_)
);

AOI21X1 _18878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8334_),
    .B(_8353_),
    .C(_8356_),
    .Y(_8728_)
);

OAI21X1 _18458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8262_),
    .B(_8266_),
    .C(_8267_),
    .Y(_8268_)
);

NOR3X1 _18038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7794_),
    .B(_7803_),
    .C(_7804_),
    .Y(_7807_)
);

AOI21X1 _13593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(_2932_),
    .C(_2930_),
    .Y(_2938_)
);

AOI21X1 _13173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2467_),
    .C(_2458_),
    .Y(_2478_)
);

NAND3X1 _23691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .B(_2031_),
    .C(_2036_),
    .Y(_2089_)
);

OR2X2 _23271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1627_),
    .Y(_1632_)
);

NOR3X1 _14798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4243_),
    .B(_4247_),
    .C(_4251_),
    .Y(_4255_)
);

OAI21X1 _14378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf2),
    .B(_3253__bF$buf2),
    .C(_3790_),
    .Y(_3796_)
);

DFFPOSX1 _24056_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[14]),
    .CLK(clk_bF$buf9),
    .D(b[14])
);

FILL SFILL64200x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10081_),
    .B(_10078_),
    .C(_10072_),
    .Y(_10392_)
);

OAI21X1 _16944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6223_),
    .B(_6606_),
    .C(_6607_),
    .Y(_6608_)
);

NAND2X1 _16524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .B(_6142_),
    .Y(_6147_)
);

OAI21X1 _16104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_5676_),
    .C(_5686_),
    .Y(_5687_)
);

NAND3X1 _17729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7457_),
    .B(_7451_),
    .C(_7455_),
    .Y(_7468_)
);

OAI21X1 _17309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7005_),
    .B(_7006_),
    .C(_7007_),
    .Y(_7008_)
);

NAND3X1 _12864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_133_),
    .B(_856_),
    .C(_900_),
    .Y(_911_)
);

NAND3X1 _12444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8084_),
    .B(_8117_),
    .C(_8139_),
    .Y(_8216_)
);

OAI21X1 _22962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1161_),
    .C(_1155_),
    .Y(_1295_)
);

NOR2X1 _12024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf0),
    .B(_2508_),
    .Y(_3613_)
);

NAND3X1 _22542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_829_),
    .B(_827_),
    .C(_822_),
    .Y(_836_)
);

NOR2X1 _22122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_6300__bF$buf3),
    .Y(_376_)
);

OAI21X1 _13649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2765_),
    .B(_2996_),
    .C(_2997_),
    .Y(_2998_)
);

NOR2X1 _13229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .B(_2345_),
    .Y(_2538_)
);

XNOR2X1 _23747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2147_),
    .B(_2148_),
    .Y(_2149_)
);

NAND2X1 _23327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1688_),
    .B(_1691_),
    .Y(_1692_)
);

FILL SFILL63800x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _17482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6811_),
    .Y(_7198_)
);

AOI21X1 _17062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6291_),
    .B(_6340_),
    .C(_6737_),
    .Y(_6738_)
);

FILL SFILL74280x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8503_),
    .B(_8488_),
    .C(_8509_),
    .Y(_8518_)
);

NOR3X1 _18267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7626_),
    .B(_7627_),
    .C(_7625_),
    .Y(_8059_)
);

OR2X2 _23080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(_1421_),
    .Y(_1422_)
);

OR2X2 _21813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_31_),
    .Y(_37_)
);

NAND3X1 _14187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3572_),
    .B(_3582_),
    .C(_3576_),
    .Y(_3587_)
);

FILL SFILL74280x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .B(_6392_),
    .C(_6398_),
    .Y(_6399_)
);

NOR2X1 _16333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5564_),
    .B(_5938_),
    .Y(_5939_)
);

BUFX2 BUFX2_insert170 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .Y(_2884__bF$buf2)
);

BUFX2 BUFX2_insert171 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .Y(_2884__bF$buf1)
);

BUFX2 BUFX2_insert172 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .Y(_2884__bF$buf0)
);

BUFX2 BUFX2_insert173 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582_),
    .Y(_6582__bF$buf3)
);

OAI21X1 _17958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf2),
    .B(_5315__bF$buf3),
    .C(_7278_),
    .Y(_7719_)
);

BUFX2 BUFX2_insert174 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582_),
    .Y(_6582__bF$buf2)
);

BUFX2 BUFX2_insert175 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582_),
    .Y(_6582__bF$buf1)
);

NAND3X1 _17538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7232_),
    .B(_7256_),
    .C(_7257_),
    .Y(_7258_)
);

BUFX2 BUFX2_insert176 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582_),
    .Y(_6582__bF$buf0)
);

OAI21X1 _17118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6795_),
    .B(_6796_),
    .C(_6420_),
    .Y(_6799_)
);

FILL SFILL69000x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert177 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_549__bF$buf4)
);

BUFX2 BUFX2_insert178 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_549__bF$buf3)
);

INVX2 _12673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10715_),
    .Y(_10726_)
);

BUFX2 BUFX2_insert179 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_549__bF$buf2)
);

OAI21X1 _12253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4127_),
    .B(_5442_),
    .C(_5552_),
    .Y(_6121_)
);

NAND2X1 _22771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_1080_),
    .Y(_1087_)
);

NAND2X1 _22351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_28_bF$buf2),
    .Y(_627_)
);

OAI21X1 _13878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3020_),
    .B(_2990_),
    .C(_3032_),
    .Y(_3249_)
);

NAND3X1 _13458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2788_),
    .C(_2787_),
    .Y(_2789_)
);

DFFPOSX1 _23976_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[30]),
    .CLK(clk_bF$buf6),
    .D(_0_[30])
);

FILL SFILL18760x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_2328_),
    .C(_2330_),
    .Y(_2333_)
);

NOR3X1 _23556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1940_),
    .C(_1941_),
    .Y(_1942_)
);

OAI21X1 _23136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(_1475_),
    .C(_1437_),
    .Y(_1484_)
);

OAI21X1 _17291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6986_),
    .B(_6987_),
    .C(_6985_),
    .Y(_6989_)
);

AOI21X1 _15604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5128_),
    .B(_5121_),
    .C(_5108_),
    .Y(_5139_)
);

AOI21X1 _18496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8301_),
    .B(_8309_),
    .C(_8288_),
    .Y(_8310_)
);

AOI21X1 _18076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7380_),
    .B(_7400_),
    .C(_7403_),
    .Y(_7849_)
);

AOI21X1 _16809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6452_),
    .B(_6453_),
    .C(_6444_),
    .Y(_6459_)
);

XOR2X1 _11944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2419_),
    .B(_2727_),
    .Y(_2738_)
);

INVX2 _21622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11728_),
    .Y(_11736_)
);

NAND2X1 _21202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10955_),
    .B(_10962_),
    .Y(_11277_)
);

FILL SFILL39000x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10419_),
    .B(_11187_),
    .C(_11231_),
    .Y(_11350_)
);

NAND3X1 _12309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6450_),
    .B(_6549_),
    .C(_6505_),
    .Y(_6736_)
);

NAND2X1 _22827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1142_),
    .Y(_1147_)
);

NAND3X1 _22407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_681_),
    .C(_682_),
    .Y(_687_)
);

AOI21X1 _16982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6334_),
    .B(_6329_),
    .C(_6293_),
    .Y(_6649_)
);

NOR3X1 _16562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6182_),
    .B(_6184_),
    .C(_6181_),
    .Y(_6189_)
);

NAND3X1 _16142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5712_),
    .B(_5717_),
    .C(_5721_),
    .Y(_5729_)
);

OAI21X1 _17767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7508_),
    .B(_7509_),
    .C(_7507_),
    .Y(_7510_)
);

OAI21X1 _17347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6666_),
    .B(_6673_),
    .C(_6675_),
    .Y(_7050_)
);

XNOR2X1 _12482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8621_),
    .B(_8577_),
    .Y(_8632_)
);

AOI21X1 _12062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3964_),
    .B(_3997_),
    .C(_3350_),
    .Y(_4030_)
);

NAND2X1 _22580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_876_),
    .Y(_877_)
);

INVX2 _22160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .Y(_417_)
);

FILL SFILL8680x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3038_),
    .B(_3037_),
    .C(_3039_),
    .Y(_3040_)
);

AOI21X1 _13267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2391_),
    .B(_2396_),
    .C(_2410_),
    .Y(_2580_)
);

OAI21X1 _23785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2129_),
    .B(_2149_),
    .C(_2189_),
    .Y(_2190_)
);

OAI22X1 _23365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4069_),
    .B(_8773_),
    .C(_5369_),
    .D(_8759_),
    .Y(_1734_)
);

INVX2 _19913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9863_),
    .Y(_9864_)
);

FILL SFILL74280x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5385_),
    .B(_5389_),
    .Y(_5390_)
);

OAI21X1 _15413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4930_),
    .C(_4925_),
    .Y(_4931_)
);

FILL SFILL43800x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5908_),
    .B(_5901_),
    .C(_5910_),
    .Y(_6250_)
);

NAND3X1 _21851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_63_),
    .B(_71_),
    .C(_68_),
    .Y(_79_)
);

NAND2X1 _21431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf2),
    .B(areg_30_bF$buf1),
    .Y(_11528_)
);

OAI21X1 _21011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11065_),
    .B(_11064_),
    .C(_11061_),
    .Y(_11067_)
);

NAND2X1 _12958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf1),
    .B(areg_8_bF$buf4),
    .Y(_1936_)
);

XNOR2X1 _12538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9016_),
    .B(_8961_),
    .Y(_9247_)
);

NAND3X1 _12118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4226_),
    .B(_4632_),
    .C(_4588_),
    .Y(_4642_)
);

NAND2X1 _22636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_937_),
    .B(_715_),
    .Y(_938_)
);

AOI21X1 _22216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11881_),
    .B(_227_),
    .C(_478_),
    .Y(_479_)
);

FILL SFILL64200x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6097_),
    .B(_6100_),
    .C(_6090_),
    .Y(_6440_)
);

NAND3X1 _16371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5961_),
    .B(_5967_),
    .C(_5971_),
    .Y(_5980_)
);

NAND2X1 _17996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7705_),
    .B(_7702_),
    .Y(_7761_)
);

AOI21X1 _17576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6948_),
    .B(_6949_),
    .C(_6932_),
    .Y(_7300_)
);

INVX1 _17156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6839_),
    .Y(_6840_)
);

AND2X2 _12291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5179_),
    .B(_6483_),
    .Y(_6538_)
);

NAND3X1 _20702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10712_),
    .B(_10705_),
    .C(_10717_),
    .Y(_10728_)
);

AND2X2 _13496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2634_),
    .B(_2636_),
    .Y(_2831_)
);

NAND2X1 _13076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1816_),
    .B(_1762_),
    .Y(_2371_)
);

AOI21X1 _23594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1862_),
    .B(_1863_),
    .C(_1949_),
    .Y(_1983_)
);

AOI21X1 _23174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(_1520_),
    .C(_1405_),
    .Y(_1526_)
);

INVX2 _19722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9653_),
    .Y(_9654_)
);

NAND3X1 _19302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9176_),
    .B(_9183_),
    .C(_9193_),
    .Y(_9194_)
);

FILL SFILL23720x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf2),
    .B(_8773_),
    .C(_11528_),
    .Y(_140_)
);

OAI21X1 _15642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5180_),
    .B(_4874_),
    .C(_4866_),
    .Y(_5181_)
);

OAI21X1 _15222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf0),
    .B(_2362__bF$buf5),
    .C(_4714_),
    .Y(_4721_)
);

OR2X2 _20299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10273_),
    .B(_10208_),
    .Y(_10286_)
);

OAI21X1 _16847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6213_),
    .B(_6206_),
    .C(_6215_),
    .Y(_6501_)
);

NAND2X1 _16427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5301_),
    .B(_6039_),
    .Y(_6040_)
);

AOI21X1 _16007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5576_),
    .B(_5575_),
    .C(_5573_),
    .Y(_5581_)
);

INVX2 _11982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3099_),
    .Y(_3154_)
);

AOI21X1 _21660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11525_),
    .B(_11529_),
    .C(_11776_),
    .Y(_11777_)
);

OAI21X1 _21240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11316_),
    .B(_11007_),
    .C(_11298_),
    .Y(_11317_)
);

FILL SFILL13720x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf3),
    .B(_8555_),
    .Y(_11756_)
);

NAND3X1 _12347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7120_),
    .B(_7142_),
    .C(_7131_),
    .Y(_7153_)
);

INVX1 _22865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .Y(_1189_)
);

NAND2X1 _22445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_670_),
    .Y(_729_)
);

NOR2X1 _22025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_261_),
    .Y(_269_)
);

FILL SFILL48840x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5757_),
    .B(_5755_),
    .Y(_5770_)
);

NAND3X1 _14913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4375_),
    .B(_4377_),
    .C(_4376_),
    .Y(_4382_)
);

AOI21X1 _17385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6707_),
    .B(_6702_),
    .C(_6694_),
    .Y(_7092_)
);

NAND3X1 _20931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10976_),
    .B(_10975_),
    .C(_10697_),
    .Y(_10980_)
);

OAI21X1 _20511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf1),
    .B(_6686__bF$buf3),
    .C(_10157_),
    .Y(_10519_)
);

FILL SFILL38840x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_31_bF$buf0),
    .Y(_9905_)
);

AOI21X1 _19531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9434_),
    .B(_9431_),
    .C(_9429_),
    .Y(_9445_)
);

OAI21X1 _19111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8981_),
    .B(_8982_),
    .C(_8980_),
    .Y(_8984_)
);

OAI21X1 _21716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11831_),
    .B(_11838_),
    .C(_11602_),
    .Y(_11839_)
);

FILL SFILL64200x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4715_),
    .B(_5411_),
    .C(_5060_),
    .Y(_5432_)
);

NAND2X1 _15451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4657_),
    .B(_4665_),
    .Y(_4971_)
);

NAND3X1 _15031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4509_),
    .B(_4510_),
    .C(_4508_),
    .Y(_4512_)
);

FILL SFILL28840x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5940_),
    .B(_5937_),
    .C(_5929_),
    .Y(_6292_)
);

OAI21X1 _16236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5825_),
    .B(_5827_),
    .C(_5828_),
    .Y(_5832_)
);

FILL SFILL54200x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_2280_),
    .Y(_2291_)
);

AOI21X1 _12576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8194_),
    .B(_8172_),
    .C(_9652_),
    .Y(_9663_)
);

NOR2X1 _12156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5036_),
    .B(_5047_),
    .Y(_5058_)
);

NAND2X1 _22674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_802_),
    .B(_810_),
    .Y(_980_)
);

AOI21X1 _22254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_519_),
    .C(_508_),
    .Y(_520_)
);

OAI21X1 _18802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_3402__bF$buf0),
    .C(_8644_),
    .Y(_8645_)
);

XOR2X1 _23879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3263_),
    .B(_3252_),
    .Y(_0_[2])
);

NAND2X1 _23459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1823_),
    .Y(_1836_)
);

AOI21X1 _23039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1377_),
    .B(_1376_),
    .C(_1266_),
    .Y(_1378_)
);

NOR2X1 _14722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4166_),
    .B(_4167_),
    .Y(_4173_)
);

AOI21X1 _14302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3711_),
    .B(_3713_),
    .C(_3710_),
    .Y(_3714_)
);

NAND3X1 _17194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(_6881_),
    .C(_6879_),
    .Y(_6882_)
);

FILL SFILL48920x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .B(_5489_),
    .C(_5472_),
    .Y(_5493_)
);

OAI21X1 _15507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5023_),
    .B(_5022_),
    .C(_5020_),
    .Y(_5032_)
);

OAI21X1 _20740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10761_),
    .B(_10760_),
    .C(_10757_),
    .Y(_10769_)
);

NAND3X1 _20320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10306_),
    .B(_10307_),
    .C(_10308_),
    .Y(_10309_)
);

INVX2 _18399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8197_),
    .Y(_8203_)
);

AND2X2 _19760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9692_),
    .B(_9693_),
    .Y(_9695_)
);

OAI21X1 _19340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9219_),
    .B(_9226_),
    .C(_9229_),
    .Y(_9235_)
);

AOI21X1 _21945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_174_),
    .C(_172_),
    .Y(_182_)
);

AOI21X1 _21525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11618_),
    .B(_11616_),
    .C(_11612_),
    .Y(_11630_)
);

NAND2X1 _21105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf3),
    .B(areg_24_bF$buf4),
    .Y(_11170_)
);

OAI21X1 _15680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5220_),
    .B(_5221_),
    .C(_5219_),
    .Y(_5222_)
);

OAI21X1 _15260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4756_),
    .B(_4755_),
    .C(_4757_),
    .Y(_4762_)
);

FILL SFILL38920x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6525_),
    .B(_6529_),
    .C(_6531_),
    .Y(_6543_)
);

NAND3X1 _16465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6059_),
    .B(_6073_),
    .C(_6080_),
    .Y(_6081_)
);

AOI21X1 _16045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5619_),
    .B(_5617_),
    .C(_5616_),
    .Y(_5623_)
);

FILL SFILL3560x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69320x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69240x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf1),
    .B(_4258__bF$buf2),
    .Y(_7569_)
);

AOI21X1 _22483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_567_),
    .C(_573_),
    .Y(_771_)
);

NAND2X1 _22063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf3),
    .B(areg_23_bF$buf0),
    .Y(_311_)
);

FILL SFILL28920x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8433_),
    .B(_8434_),
    .C(_8432_),
    .Y(_8436_)
);

NOR2X1 _23688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2028_),
    .B(_2084_),
    .Y(_2085_)
);

NOR2X1 _23268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1513_),
    .Y(_1628_)
);

NAND2X1 _19816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9465_),
    .B(_9471_),
    .Y(_9757_)
);

AOI21X1 _14951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4421_),
    .B(_4422_),
    .C(_4415_),
    .Y(_4424_)
);

INVX2 _14531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3957_),
    .Y(_3965_)
);

OAI21X1 _14111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3502_),
    .B(_1391_),
    .C(_2537_),
    .Y(_3504_)
);

FILL SFILL18920x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4965_),
    .B(_5279_),
    .C(_5283_),
    .Y(_5284_)
);

NAND3X1 _15316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4819_),
    .B(_4823_),
    .C(_4822_),
    .Y(_4824_)
);

BUFX2 BUFX2_insert80 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[22]),
    .Y(breg_22_bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[22]),
    .Y(breg_22_bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[22]),
    .Y(breg_22_bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[22]),
    .Y(breg_22_bF$buf0)
);

NOR3X1 _21754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11845_),
    .B(_11850_),
    .C(_11848_),
    .Y(_11880_)
);

OAI21X1 _21334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11416_),
    .B(_11415_),
    .C(_11369_),
    .Y(_11421_)
);

FILL SFILL38920x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf3),
    .B(_7225__bF$buf0),
    .Y(_1291_)
);

OAI21X1 _22539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(_831_),
    .C(_829_),
    .Y(_832_)
);

NOR2X1 _22119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_370_),
    .Y(_371_)
);

NAND3X1 _13802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3158_),
    .B(_3140_),
    .C(_3162_),
    .Y(_3167_)
);

BUFX2 _23900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[18]),
    .Y(y[18])
);

NAND3X1 _16694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6331_),
    .B(_6333_),
    .C(_6332_),
    .Y(_6334_)
);

AOI21X1 _16274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5868_),
    .B(_5869_),
    .C(_5867_),
    .Y(_5874_)
);

FILL SFILL53880x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7653_),
    .B(_6843_),
    .C(_7622_),
    .Y(_7654_)
);

AOI21X1 _17479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7177_),
    .B(_7182_),
    .C(_6919_),
    .Y(_7194_)
);

NAND3X1 _17059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6733_),
    .B(_6732_),
    .C(_6731_),
    .Y(_6734_)
);

OAI21X1 _12194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4127_),
    .B(_5442_),
    .C(_5464_),
    .Y(_5475_)
);

OAI21X1 _22292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf3),
    .B(_5318_),
    .C(_548_),
    .Y(_562_)
);

NAND3X1 _18840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8602_),
    .B(_8685_),
    .C(_8681_),
    .Y(_8686_)
);

NAND2X1 _18420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_17_bF$buf1),
    .Y(_8226_)
);

AOI21X1 _18000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7414_),
    .B(_7419_),
    .C(_7421_),
    .Y(_7765_)
);

AOI21X1 _20605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10616_),
    .B(_10621_),
    .C(_10460_),
    .Y(_10622_)
);

AOI21X1 _13399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2719_),
    .B(_2720_),
    .C(_2576_),
    .Y(_2725_)
);

AND2X2 _23497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(_1788_),
    .Y(_1877_)
);

OAI21X1 _23077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1416_),
    .B(_1417_),
    .C(_1418_),
    .Y(_1419_)
);

OAI21X1 _19625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9547_),
    .B(_9546_),
    .C(_9530_),
    .Y(_9548_)
);

NAND3X1 _19205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9070_),
    .B(_9039_),
    .C(_9077_),
    .Y(_9086_)
);

OAI21X1 _14760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf4),
    .B(_2465__bF$buf0),
    .C(_4210_),
    .Y(_4214_)
);

AOI21X1 _14340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3246_),
    .B(_3474_),
    .C(_3754_),
    .Y(_3755_)
);

FILL SFILL48760x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _15965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .Y(_5535_)
);

NAND3X1 _15545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5064_),
    .B(_5051_),
    .C(_5054_),
    .Y(_5074_)
);

OAI21X1 _15125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4609_),
    .B(_4611_),
    .C(_4361_),
    .Y(_4615_)
);

FILL SFILL48680x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_223_),
    .C(_220_),
    .Y(_224_)
);

NAND3X1 _21563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11649_),
    .B(_11664_),
    .C(_11670_),
    .Y(_11671_)
);

AOI21X1 _21143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10910_),
    .B(_10943_),
    .C(_11211_),
    .Y(_11212_)
);

FILL SFILL49000x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_947_),
    .B(_1082_),
    .C(_1081_),
    .Y(_1083_)
);

OAI21X1 _22348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_7520__bF$buf1),
    .C(_378_),
    .Y(_623_)
);

NAND3X1 _13611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2953_),
    .B(_2956_),
    .C(_2755_),
    .Y(_2958_)
);

NOR3X1 _16083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5652_),
    .B(_5650_),
    .C(_5647_),
    .Y(_5664_)
);

FILL SFILL39080x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4274_),
    .B(_4275_),
    .Y(_4276_)
);

INVX2 _17288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6960_),
    .Y(_6985_)
);

FILL SFILL18760x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf2),
    .B(_7100__bF$buf1),
    .C(_10511_),
    .Y(_10873_)
);

NOR3X1 _20414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10395_),
    .B(_10399_),
    .C(_10400_),
    .Y(_10412_)
);

OAI22X1 _19854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_4551__bF$buf0),
    .C(_2560__bF$buf2),
    .D(_3961__bF$buf0),
    .Y(_9799_)
);

NOR3X1 _19434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9322_),
    .B(_9326_),
    .C(_9327_),
    .Y(_9338_)
);

INVX1 _19014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8471_),
    .Y(_8877_)
);

AND2X2 _21619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_25_bF$buf3),
    .Y(_11732_)
);

NAND3X1 _15774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5317_),
    .B(_5322_),
    .C(_5324_),
    .Y(_5325_)
);

NAND3X1 _15354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4865_),
    .B(_4861_),
    .C(_4854_),
    .Y(_4866_)
);

NAND3X1 _16979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6630_),
    .B(_6635_),
    .C(_6636_),
    .Y(_6646_)
);

OAI21X1 _16559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6181_),
    .B(_6182_),
    .C(_6184_),
    .Y(_6185_)
);

NAND3X1 _16139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5669_),
    .B(_5718_),
    .C(_5724_),
    .Y(_5725_)
);

AOI21X1 _21792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_13_),
    .B(_9_),
    .C(_11892_),
    .Y(_14_)
);

OAI21X1 _21372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11453_),
    .B(_11449_),
    .C(_11447_),
    .Y(_11463_)
);

OAI21X1 _17920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf0),
    .B(_5668__bF$buf3),
    .C(_7243_),
    .Y(_7677_)
);

NAND2X1 _17500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7197_),
    .B(_7201_),
    .Y(_7216_)
);

AOI21X1 _12899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11636_),
    .B(_1271_),
    .C(_1282_),
    .Y(_1293_)
);

NAND2X1 _12479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg_10_bF$buf5),
    .Y(_8599_)
);

OAI21X1 _22997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1327_),
    .B(_1328_),
    .C(_1295_),
    .Y(_1332_)
);

NAND2X1 _12059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3372_),
    .B(_3986_),
    .Y(_3997_)
);

NOR2X1 _22577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_872_),
    .Y(_874_)
);

INVX1 _22157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .Y(_414_)
);

FILL SFILL3720x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _18705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8531_),
    .B(_8532_),
    .Y(_8538_)
);

NAND3X1 _13840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3199_),
    .B(_3202_),
    .C(_3049_),
    .Y(_3208_)
);

NAND3X1 _13420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2745_),
    .B(_2746_),
    .C(_2747_),
    .Y(_2748_)
);

OAI21X1 _13000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_527_),
    .B(_2294_),
    .C(_2288_),
    .Y(_2295_)
);

FILL SFILL3640x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3845_),
    .B(_3846_),
    .Y(_4066_)
);

AOI21X1 _14205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3603_),
    .B(_3605_),
    .C(_3601_),
    .Y(_3606_)
);

AOI21X1 _17097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6756_),
    .B(_6763_),
    .C(_6511_),
    .Y(_6776_)
);

OAI21X1 _20643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8068_),
    .B(_10662_),
    .C(_8466_),
    .Y(_10663_)
);

NAND3X1 _20223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10190_),
    .B(_10181_),
    .C(_10192_),
    .Y(_10203_)
);

NAND3X1 _19663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9588_),
    .B(_9589_),
    .C(_9586_),
    .Y(_9590_)
);

AOI21X1 _19243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8766_),
    .B(_8762_),
    .C(_8767_),
    .Y(_9129_)
);

FILL SFILL33880x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_74_),
    .C(_24_),
    .Y(_75_)
);

AOI21X1 _21428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11234_),
    .B(_11523_),
    .C(_11243_),
    .Y(_11524_)
);

NAND2X1 _21008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf5),
    .B(breg_24_bF$buf1),
    .Y(_11063_)
);

OAI21X1 _15583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_2669__bF$buf2),
    .C(_4783_),
    .Y(_5116_)
);

OAI21X1 _15163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4655_),
    .B(_4614_),
    .C(_4606_),
    .Y(_4656_)
);

FILL SFILL39080x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6435_),
    .Y(_6436_)
);

OAI21X1 _16368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5877_),
    .B(_5873_),
    .C(_5879_),
    .Y(_5977_)
);

OAI21X1 _21181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11219_),
    .B(_11224_),
    .C(_11252_),
    .Y(_11254_)
);

FILL SFILL23880x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6472_),
    .B(_6494_),
    .Y(_6505_)
);

AOI21X1 _22386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_651_),
    .C(_641_),
    .Y(_665_)
);

OAI21X1 _18934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8783_),
    .B(_8789_),
    .C(_8741_),
    .Y(_8790_)
);

NAND2X1 _18514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8324_),
    .B(_8329_),
    .Y(_8330_)
);

FILL SFILL8760x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _19719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9649_),
    .Y(_9650_)
);

OAI21X1 _14854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4312_),
    .B(_4313_),
    .C(_4065_),
    .Y(_4318_)
);

AOI21X1 _14434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3593_),
    .B(_3627_),
    .C(_3636_),
    .Y(_3858_)
);

INVX2 _14014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3397_),
    .Y(_3398_)
);

FILL SFILL29000x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5174_),
    .B(_5175_),
    .C(_5176_),
    .Y(_5177_)
);

OAI22X1 _15219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf3),
    .B(_2560__bF$buf4),
    .C(_6582__bF$buf2),
    .D(_2362__bF$buf5),
    .Y(_4717_)
);

XNOR2X1 _20872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10914_),
    .B(_10911_),
    .Y(_10915_)
);

OAI21X1 _20452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10451_),
    .B(_10450_),
    .C(_10453_),
    .Y(_10454_)
);

OAI21X1 _20032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9677_),
    .B(_9647_),
    .C(_9684_),
    .Y(_9993_)
);

AOI21X1 _19892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9483_),
    .B(_9522_),
    .C(_9840_),
    .Y(_9841_)
);

AOI21X1 _19472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9006_),
    .B(_9084_),
    .C(_9093_),
    .Y(_9380_)
);

OAI21X1 _19052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8918_),
    .B(_8911_),
    .C(_8897_),
    .Y(_8919_)
);

OAI21X1 _11979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2661_),
    .C(_2475_),
    .Y(_3131_)
);

AOI21X1 _21657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11772_),
    .B(_11773_),
    .C(_11771_),
    .Y(_11774_)
);

FILL SFILL3720x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10688_),
    .B(_11313_),
    .Y(_11314_)
);

FILL SFILL43960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _12920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11712_),
    .B(_1511_),
    .Y(_1522_)
);

NAND3X1 _12500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8797_),
    .B(_8819_),
    .C(_8808_),
    .Y(_8830_)
);

NOR3X1 _15392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4581_),
    .B(_4582_),
    .C(_4580_),
    .Y(_4908_)
);

INVX1 _13705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3059_),
    .Y(_3060_)
);

OR2X2 _23803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2208_),
    .B(_2118_),
    .Y(_2209_)
);

NAND2X1 _16597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_17_bF$buf4),
    .Y(_6227_)
);

NAND3X1 _16177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5761_),
    .B(_5763_),
    .C(_5762_),
    .Y(_5767_)
);

NAND2X1 _12097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_4401_),
    .Y(_4412_)
);

XOR2X1 _22195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_203_),
    .Y(_456_)
);

OAI21X1 _18743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8578_),
    .B(_8579_),
    .C(_8574_),
    .Y(_8580_)
);

NAND3X1 _18323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8080_),
    .B(_8119_),
    .C(_8118_),
    .Y(_8120_)
);

FILL SFILL33880x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10963_),
    .B(_10811_),
    .C(_10958_),
    .Y(_10976_)
);

AOI21X1 _20508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10508_),
    .B(_10509_),
    .C(_10500_),
    .Y(_10515_)
);

NAND2X1 _19948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_30_bF$buf2),
    .Y(_9901_)
);

AOI21X1 _19528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9099_),
    .B(_9440_),
    .C(_9439_),
    .Y(_9441_)
);

AOI21X1 _19108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8528_),
    .B(_8565_),
    .C(_8569_),
    .Y(_8980_)
);

OAI21X1 _14663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf2),
    .B(_2763_),
    .C(_4107_),
    .Y(_4108_)
);

INVX1 _14243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3642_),
    .Y(_3649_)
);

AOI21X1 _15868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5130_),
    .B(_5427_),
    .C(_5426_),
    .Y(_5428_)
);

NOR2X1 _15448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4671_),
    .B(_4966_),
    .Y(_4967_)
);

INVX1 _15028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4502_),
    .Y(_4508_)
);

OAI21X1 _20681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10367_),
    .B(_10357_),
    .C(_10361_),
    .Y(_10705_)
);

FILL SFILL23880x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10210_),
    .B(_10238_),
    .C(_10243_),
    .Y(_10245_)
);

FILL SFILL39000x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9161_),
    .B(_9162_),
    .C(_9158_),
    .Y(_9171_)
);

NAND3X1 _21886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_113_),
    .C(_112_),
    .Y(_117_)
);

AOI21X1 _21466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11565_),
    .B(_11558_),
    .C(_11324_),
    .Y(_11566_)
);

NAND3X1 _21046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11083_),
    .B(_11087_),
    .C(_11095_),
    .Y(_11105_)
);

FILL FILL73960x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3070_),
    .B(_3078_),
    .Y(_3311_)
);

OAI21X1 _13514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2638_),
    .B(_2849_),
    .C(_2850_),
    .Y(_2851_)
);

OAI21X1 _23612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1882_),
    .B(_1883_),
    .C(_1889_),
    .Y(_2003_)
);

FILL SFILL53960x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _14719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_549__bF$buf3),
    .C(_7217__bF$buf0),
    .D(_10869__bF$buf3),
    .Y(_4169_)
);

AOI21X1 _18972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8829_),
    .B(_8831_),
    .C(_8828_),
    .Y(_8832_)
);

AND2X2 _18552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8346_),
    .B(_8364_),
    .Y(_8372_)
);

NAND3X1 _18132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7902_),
    .B(_7888_),
    .C(_7906_),
    .Y(_7911_)
);

NAND3X1 _20737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10743_),
    .B(_10758_),
    .C(_10765_),
    .Y(_10766_)
);

INVX2 _20317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9996_),
    .Y(_10306_)
);

FILL SFILL43960x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_25_bF$buf5),
    .Y(_9692_)
);

NAND3X1 _19337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9231_),
    .B(_9230_),
    .C(_9229_),
    .Y(_9232_)
);

XOR2X1 _14892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4358_),
    .B(_4356_),
    .Y(_4359_)
);

AOI21X1 _14472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3899_),
    .B(_3897_),
    .C(_3896_),
    .Y(_3900_)
);

AOI21X1 _14052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3439_),
    .B(_3437_),
    .C(_3431_),
    .Y(_3440_)
);

AOI21X1 _15677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4853_),
    .B(_4870_),
    .C(_5218_),
    .Y(_5219_)
);

OAI21X1 _15257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4758_),
    .B(_4754_),
    .C(_4677_),
    .Y(_4759_)
);

NOR2X1 _20490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10490_),
    .B(_10494_),
    .Y(_10495_)
);

NOR3X1 _20070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10019_),
    .B(_10005_),
    .C(_10026_),
    .Y(_10034_)
);

INVX1 _19090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8936_),
    .Y(_8960_)
);

NOR2X1 _21695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11814_),
    .B(_11815_),
    .Y(_11816_)
);

NAND3X1 _21275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11340_),
    .B(_11344_),
    .C(_11333_),
    .Y(_11355_)
);

OAI21X1 _17823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7570_),
    .B(_7571_),
    .C(_7568_),
    .Y(_7572_)
);

NAND2X1 _17403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6698_),
    .B(_7111_),
    .Y(_7112_)
);

NAND2X1 _18608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8431_),
    .B(_8430_),
    .Y(_8432_)
);

AND2X2 _13743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf5),
    .B(areg_11_bF$buf0),
    .Y(_3102_)
);

NOR2X1 _13323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2630_),
    .B(_2640_),
    .Y(_2642_)
);

NOR2X1 _23841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815__bF$buf3),
    .B(_8773_),
    .Y(_2250_)
);

NAND2X1 _23421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_27_bF$buf1),
    .B(breg_28_bF$buf5),
    .Y(_1795_)
);

AOI21X1 _23001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1333_),
    .B(_1332_),
    .C(_1331_),
    .Y(_1337_)
);

AOI21X1 _14948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4099_),
    .B(_4120_),
    .C(_4123_),
    .Y(_4420_)
);

INVX8 _14528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf3),
    .Y(_3961_)
);

NAND3X1 _14108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2538_),
    .B(_2745_),
    .C(_3499_),
    .Y(_3500_)
);

AOI21X1 _18781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8203_),
    .B(_8206_),
    .C(_8212_),
    .Y(_8622_)
);

NAND3X1 _18361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8156_),
    .B(_8160_),
    .C(_8122_),
    .Y(_8162_)
);

FILL SFILL23800x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11016_),
    .Y(_11017_)
);

NAND2X1 _20546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf0),
    .B(areg_25_bF$buf3),
    .Y(_10557_)
);

OAI21X1 _20126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9849_),
    .B(_9851_),
    .C(_9847_),
    .Y(_10096_)
);

NOR2X1 _19986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9855_),
    .B(_9928_),
    .Y(_9943_)
);

NAND2X1 _19566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9125_),
    .B(_9131_),
    .Y(_9483_)
);

NAND3X1 _19146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9017_),
    .B(_9021_),
    .C(_9020_),
    .Y(_9022_)
);

AOI21X1 _14281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3398_),
    .B(_3404_),
    .C(_3408_),
    .Y(_3691_)
);

FILL SFILL13880x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4739_),
    .B(_4747_),
    .Y(_5009_)
);

AOI21X1 _15066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4244_),
    .B(_4248_),
    .C(_4251_),
    .Y(_4550_)
);

FILL SFILL74120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _21084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11140_),
    .Y(_11147_)
);

INVX2 _17632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7353_),
    .Y(_7362_)
);

NAND3X1 _17212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6894_),
    .B(_6844_),
    .C(_6901_),
    .Y(_6902_)
);

FILL SFILL3960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _22289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .Y(_558_)
);

NAND3X1 _18837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8667_),
    .B(_8673_),
    .C(_8635_),
    .Y(_8683_)
);

OAI21X1 _18417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7852_),
    .B(_7819_),
    .C(_7845_),
    .Y(_8223_)
);

INVX1 _13972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3070_),
    .Y(_3352_)
);

AOI21X1 _13552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2885_),
    .B(_2883_),
    .C(_2879_),
    .Y(_2892_)
);

OAI22X1 _13132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_2432_),
    .C(_2163_),
    .D(_2196_),
    .Y(_2433_)
);

XNOR2X1 _23650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2043_),
    .B(_2000_),
    .Y(_2044_)
);

NAND2X1 _23230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .B(_1581_),
    .Y(_1585_)
);

FILL SFILL28680x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4209_),
    .B(_4210_),
    .Y(_4211_)
);

AOI21X1 _14337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3751_),
    .B(_3750_),
    .C(_3520_),
    .Y(_3752_)
);

DFFPOSX1 _24015_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[5]),
    .CLK(clk_bF$buf10),
    .D(a[5])
);

NAND3X1 _18590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8392_),
    .B(_8399_),
    .C(_8330_),
    .Y(_8412_)
);

OAI21X1 _18170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7945_),
    .B(_7946_),
    .C(_7943_),
    .Y(_7952_)
);

NAND3X1 _20775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10798_),
    .B(_10804_),
    .C(_10794_),
    .Y(_10808_)
);

AOI21X1 _20355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10282_),
    .B(_10275_),
    .C(_10109_),
    .Y(_10347_)
);

OAI22X1 _16903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6177_),
    .B(_6561_),
    .C(_6562_),
    .D(_6222_),
    .Y(_6563_)
);

AOI21X1 _19795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9722_),
    .B(_9717_),
    .C(_9689_),
    .Y(_9734_)
);

NAND2X1 _19375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8991_),
    .B(_8997_),
    .Y(_9273_)
);

NOR3X1 _14090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3204_),
    .B(_3211_),
    .C(_3214_),
    .Y(_3481_)
);

FILL SFILL59240x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_451_),
    .Y(_462_)
);

OAI21X1 _12403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7755_),
    .B(_7744_),
    .C(_7667_),
    .Y(_7766_)
);

OAI21X1 _22921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1248_),
    .B(_1249_),
    .C(_1100_),
    .Y(_1251_)
);

NOR3X1 _22501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_776_),
    .C(_778_),
    .Y(_791_)
);

AOI21X1 _15295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4793_),
    .B(_4799_),
    .C(_4800_),
    .Y(_4801_)
);

OAI21X1 _13608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2950_),
    .B(_2951_),
    .C(_2760_),
    .Y(_2954_)
);

AND2X2 _23706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2104_),
    .B(_2103_),
    .Y(_2105_)
);

FILL SFILL44040x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6919_),
    .B(_7182_),
    .C(_7612_),
    .Y(_7613_)
);

AOI21X1 _17441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7135_),
    .B(_7140_),
    .C(_7091_),
    .Y(_7154_)
);

AND2X2 _17021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6688_),
    .B(_6691_),
    .Y(_6693_)
);

NAND2X1 _22098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_292_),
    .B(_289_),
    .Y(_349_)
);

OAI21X1 _18646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8472_),
    .B(_8072_),
    .C(_8454_),
    .Y(_8473_)
);

NAND3X1 _18226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7873_),
    .B(_7867_),
    .C(_7871_),
    .Y(_8014_)
);

AND2X2 _13781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_3144_)
);

OAI21X1 _13361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2681_),
    .B(_2682_),
    .C(_2680_),
    .Y(_2684_)
);

FILL SFILL69160x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_2287__bF$buf0),
    .C(_4460_),
    .Y(_4461_)
);

NAND3X1 _14566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .B(_4002_),
    .C(_4000_),
    .Y(_4003_)
);

NAND2X1 _14146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_15_bF$buf1),
    .Y(_3542_)
);

FILL SFILL28920x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10586_),
    .B(_10589_),
    .C(_10556_),
    .Y(_10599_)
);

NAND3X1 _20164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10132_),
    .B(_10117_),
    .C(_10133_),
    .Y(_10138_)
);

AOI21X1 _16712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6335_),
    .B(_6340_),
    .C(_6291_),
    .Y(_6354_)
);

AOI21X1 _19184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9056_),
    .B(_9063_),
    .C(_9042_),
    .Y(_9064_)
);

FILL SFILL59160x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6_),
    .B(_7_),
    .C(_3_),
    .Y(_10_)
);

OAI21X1 _21369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11454_),
    .B(_11458_),
    .C(_11446_),
    .Y(_11459_)
);

FILL SFILL64120x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_28_bF$buf0),
    .Y(_7674_)
);

OAI21X1 _12632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10189_),
    .B(_10233_),
    .C(_10068_),
    .Y(_10277_)
);

NAND3X1 _12212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5003_),
    .B(_5289_),
    .C(_5332_),
    .Y(_5672_)
);

OR2X2 _22730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .B(_853_),
    .Y(_1041_)
);

NAND3X1 _22310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_572_),
    .C(_577_),
    .Y(_581_)
);

NAND3X1 _13837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3042_),
    .B(_3036_),
    .C(_3040_),
    .Y(_3205_)
);

NAND3X1 _13417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2350_),
    .B(_2531_),
    .C(_2527_),
    .Y(_2745_)
);

BUFX2 _23935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[53]),
    .Y(y[53])
);

NAND2X1 _23515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1894_),
    .B(_1895_),
    .Y(_1896_)
);

FILL FILL74040x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _17670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7397_),
    .B(_7399_),
    .C(_7396_),
    .Y(_7403_)
);

OAI21X1 _17250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf0),
    .B(_3529__bF$buf1),
    .C(_6533_),
    .Y(_6943_)
);

FILL SFILL54120x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8716_),
    .B(_8702_),
    .C(_8721_),
    .Y(_8725_)
);

OAI21X1 _18455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8247_),
    .B(_8253_),
    .C(_8255_),
    .Y(_8265_)
);

NOR2X1 _18035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7796_),
    .B(_7797_),
    .Y(_7804_)
);

NAND3X1 _13590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2933_),
    .B(_2925_),
    .C(_2793_),
    .Y(_2934_)
);

NAND3X1 _13170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2470_),
    .C(_2473_),
    .Y(_2474_)
);

OAI21X1 _14795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4251_),
    .B(_4247_),
    .C(_4243_),
    .Y(_4252_)
);

OAI21X1 _14375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3792_),
    .B(_3791_),
    .C(_3789_),
    .Y(_3793_)
);

DFFPOSX1 _24053_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[11]),
    .CLK(clk_bF$buf1),
    .D(b[11])
);

FILL SFILL44040x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10352_),
    .B(_10380_),
    .C(_10377_),
    .Y(_10389_)
);

NOR2X1 _16941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_2465__bF$buf1),
    .Y(_6605_)
);

NOR2X1 _16521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6141_),
    .B(_6142_),
    .Y(_6144_)
);

NAND3X1 _16101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5677_),
    .B(_5682_),
    .C(_5680_),
    .Y(_5684_)
);

INVX1 _21598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11411_),
    .Y(_11709_)
);

OR2X2 _21178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11246_),
    .B(_11235_),
    .Y(_11250_)
);

INVX2 _17726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7439_),
    .Y(_7465_)
);

AOI21X1 _17306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7000_),
    .B(_7001_),
    .C(_6998_),
    .Y(_7005_)
);

AOI21X1 _12861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_823_),
    .B(_834_),
    .C(_812_),
    .Y(_878_)
);

FILL SFILL69240x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7185_),
    .B(_8172_),
    .C(_8128_),
    .Y(_8183_)
);

NOR2X1 _12021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_3569_),
    .Y(_3580_)
);

FILL SFILL69160x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .B(_2994_),
    .Y(_2995_)
);

NAND2X1 _13226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2535_),
    .B(_2534_),
    .Y(_2536_)
);

XNOR2X1 _23744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2145_),
    .B(_2134_),
    .Y(_2146_)
);

OR2X2 _23324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1671_),
    .B(_1684_),
    .Y(_1689_)
);

FILL SFILL3800x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8514_),
    .B(_8510_),
    .C(_8486_),
    .Y(_8515_)
);

OAI21X1 _18264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8039_),
    .B(_8044_),
    .C(_8047_),
    .Y(_8056_)
);

FILL SFILL59160x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf0),
    .B(areg_26_bF$buf4),
    .Y(_10911_)
);

AOI21X1 _20449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10445_),
    .B(_10446_),
    .C(_10444_),
    .Y(_10450_)
);

OAI21X1 _20029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9632_),
    .B(_9988_),
    .C(_9986_),
    .Y(_9989_)
);

AOI22X1 _21810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf1),
    .B(breg_25_bF$buf2),
    .C(areg_20_bF$buf4),
    .D(breg_24_bF$buf0),
    .Y(_33_)
);

OAI21X1 _19889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9815_),
    .B(_9821_),
    .C(_9823_),
    .Y(_9837_)
);

NAND3X1 _19469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9374_),
    .B(_9375_),
    .C(_9370_),
    .Y(_9376_)
);

AOI21X1 _19049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8913_),
    .B(_8914_),
    .C(_8899_),
    .Y(_8915_)
);

NAND3X1 _14184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3578_),
    .B(_3523_),
    .C(_3583_),
    .Y(_3584_)
);

FILL FILL74120x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11866_),
    .B(_11811_),
    .Y(_1489_)
);

AOI21X1 _15389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4885_),
    .B(_4891_),
    .C(_4814_),
    .Y(_4904_)
);

FILL SFILL49160x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6390_),
    .B(_6389_),
    .C(_6388_),
    .Y(_6395_)
);

INVX2 _16330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5934_),
    .Y(_5935_)
);

FILL SFILL18680x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert140 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf6)
);

BUFX2 BUFX2_insert141 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf5)
);

BUFX2 BUFX2_insert142 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf4)
);

BUFX2 BUFX2_insert143 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf3)
);

OAI21X1 _17955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7715_),
    .B(_7714_),
    .C(_7712_),
    .Y(_7716_)
);

BUFX2 BUFX2_insert144 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf2)
);

OAI21X1 _17535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7254_),
    .B(_7247_),
    .C(_7233_),
    .Y(_7255_)
);

BUFX2 BUFX2_insert145 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf1)
);

BUFX2 BUFX2_insert146 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(breg_1_bF$buf0)
);

AOI21X1 _17115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6786_),
    .B(_6778_),
    .C(_6421_),
    .Y(_6796_)
);

BUFX2 BUFX2_insert147 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .Y(_2376__bF$buf3)
);

BUFX2 BUFX2_insert148 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .Y(_2376__bF$buf2)
);

NAND2X1 _12670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10639_),
    .B(_10682_),
    .Y(_10693_)
);

BUFX2 BUFX2_insert149 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .Y(_2376__bF$buf1)
);

XNOR2X1 _12250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6087_),
    .B(_6055_),
    .Y(_6088_)
);

FILL SFILL23960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3036_),
    .B(_3041_),
    .Y(_3246_)
);

NAND3X1 _13455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2761_),
    .B(_2782_),
    .C(_2785_),
    .Y(_2786_)
);

DFFPOSX1 _23973_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[27]),
    .CLK(clk_bF$buf7),
    .D(_0_[27])
);

AOI21X1 _13035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2317_),
    .B(_2321_),
    .C(_1881_),
    .Y(_2330_)
);

INVX2 _23553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .Y(_1939_)
);

AOI21X1 _23133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1464_),
    .B(_1469_),
    .C(_1437_),
    .Y(_1481_)
);

OAI21X1 _15601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4817_),
    .B(_4843_),
    .C(_4834_),
    .Y(_5136_)
);

NOR2X1 _18493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8294_),
    .B(_8291_),
    .Y(_8307_)
);

OAI21X1 _18073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7836_),
    .B(_7837_),
    .C(_7834_),
    .Y(_7846_)
);

OAI21X1 _20678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10369_),
    .B(_10355_),
    .C(_10379_),
    .Y(_10701_)
);

OAI21X1 _20258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10235_),
    .B(_10236_),
    .C(_10215_),
    .Y(_10241_)
);

AND2X2 _16806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6070_),
    .B(_6134_),
    .Y(_6456_)
);

FILL SFILL69240x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2694_),
    .C(_2628_),
    .Y(_2705_)
);

NAND3X1 _19698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9626_),
    .B(_9627_),
    .C(_9625_),
    .Y(_9628_)
);

INVX1 _19278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .Y(_9167_)
);

NOR3X1 _12726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9455_),
    .B(_9444_),
    .C(_9433_),
    .Y(_11308_)
);

NAND3X1 _12306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6352_),
    .B(_6658_),
    .C(_6692_),
    .Y(_6703_)
);

NAND2X1 _22824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf2),
    .B(areg_25_bF$buf1),
    .Y(_1144_)
);

OAI21X1 _22404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_679_),
    .C(_497_),
    .Y(_684_)
);

NAND2X1 _15198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_19_bF$buf2),
    .Y(_4694_)
);

FILL SFILL3800x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _23609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1818_),
    .C(_1911_),
    .Y(_1999_)
);

FILL SFILL59240x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7085_),
    .B(_7493_),
    .C(_7073_),
    .Y(_7507_)
);

OAI21X1 _17344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7040_),
    .B(_7041_),
    .C(_7024_),
    .Y(_7047_)
);

NAND2X1 _18969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8827_),
    .B(_8826_),
    .Y(_8828_)
);

NAND2X1 _18549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_29_bF$buf0),
    .Y(_8368_)
);

NAND3X1 _18129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7901_),
    .B(_7902_),
    .C(_7906_),
    .Y(_7907_)
);

AOI21X1 _13684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3032_),
    .B(_3031_),
    .C(_3030_),
    .Y(_3037_)
);

FILL FILL74200x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2576_),
    .Y(_2577_)
);

INVX1 _23782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2186_),
    .Y(_2187_)
);

NAND2X1 _23362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1692_),
    .B(_1721_),
    .Y(_1731_)
);

XNOR2X1 _19910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9859_),
    .B(_9857_),
    .Y(_9860_)
);

FILL SFILL49240x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4095_),
    .B(_4353_),
    .Y(_4355_)
);

XNOR2X1 _14469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .B(_3895_),
    .Y(_3896_)
);

AOI21X1 _14049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3180_),
    .B(_3126_),
    .C(_3185_),
    .Y(_3436_)
);

FILL SFILL18760x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf3),
    .B(_3529__bF$buf3),
    .C(_5385_),
    .Y(_5386_)
);

NAND3X1 _15410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4909_),
    .B(_4899_),
    .C(_4905_),
    .Y(_4927_)
);

NAND3X1 _20487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10483_),
    .B(_10469_),
    .C(_10488_),
    .Y(_10492_)
);

AOI21X1 _20067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10030_),
    .B(_10027_),
    .C(_10003_),
    .Y(_10031_)
);

OAI21X1 _16615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6240_),
    .B(_6241_),
    .C(_6226_),
    .Y(_6247_)
);

AOI21X1 _19087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8604_),
    .B(_8956_),
    .C(_8955_),
    .Y(_8957_)
);

NOR2X1 _12955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10463_),
    .B(_177_),
    .Y(_1913_)
);

AOI21X1 _12535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9115_),
    .B(_9103_),
    .C(_9060_),
    .Y(_9214_)
);

NOR3X1 _12115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4544_),
    .B(_4566_),
    .C(_4555_),
    .Y(_4610_)
);

OAI21X1 _22633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_904_),
    .C(_910_),
    .Y(_935_)
);

AOI21X1 _22213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_474_),
    .B(_475_),
    .C(_243_),
    .Y(_476_)
);

NAND2X1 _23838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_30_bF$buf0),
    .B(breg[31]),
    .Y(_2246_)
);

NOR2X1 _23418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1678_),
    .B(_1681_),
    .Y(_1791_)
);

BUFX2 BUFX2_insert520 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .Y(_3958__bF$buf0)
);

BUFX2 BUFX2_insert521 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .Y(_2562__bF$buf4)
);

BUFX2 BUFX2_insert522 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .Y(_2562__bF$buf3)
);

BUFX2 BUFX2_insert523 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .Y(_2562__bF$buf2)
);

AOI21X1 _17993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7743_),
    .B(_7738_),
    .C(_7709_),
    .Y(_7758_)
);

BUFX2 BUFX2_insert524 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .Y(_2562__bF$buf1)
);

BUFX2 BUFX2_insert525 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .Y(_2562__bF$buf0)
);

NAND3X1 _17573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7292_),
    .B(_7280_),
    .C(_7285_),
    .Y(_7297_)
);

AOI21X1 _17153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6835_),
    .B(_6836_),
    .C(_6833_),
    .Y(_6837_)
);

BUFX2 BUFX2_insert526 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .Y(_2465__bF$buf4)
);

FILL SFILL13960x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert527 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .Y(_2465__bF$buf3)
);

BUFX2 BUFX2_insert528 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .Y(_2465__bF$buf2)
);

BUFX2 BUFX2_insert529 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .Y(_2465__bF$buf1)
);

OAI22X1 _18778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf3),
    .B(_3253__bF$buf1),
    .C(_2669__bF$buf1),
    .D(_3529__bF$buf4),
    .Y(_8618_)
);

NAND3X1 _18358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8144_),
    .B(_8148_),
    .C(_8154_),
    .Y(_8158_)
);

NAND3X1 _13493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2820_),
    .B(_2824_),
    .C(_2827_),
    .Y(_2828_)
);

FILL SFILL59320x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .B(_2366_),
    .Y(_2368_)
);

AOI21X1 _23591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1973_),
    .B(_11873_),
    .C(_1978_),
    .Y(_1980_)
);

OAI21X1 _23171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1517_),
    .C(_1516_),
    .Y(_1523_)
);

OAI21X1 _21904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf3),
    .B(_7520__bF$buf1),
    .C(_131_),
    .Y(_137_)
);

NAND3X1 _14698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4067_),
    .B(_4141_),
    .C(_4145_),
    .Y(_4146_)
);

INVX2 _14278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3682_),
    .Y(_3687_)
);

NAND3X1 _20296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10282_),
    .B(_10275_),
    .C(_10109_),
    .Y(_10283_)
);

NOR3X1 _16844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6491_),
    .B(_6496_),
    .C(_6497_),
    .Y(_6498_)
);

AND2X2 _16424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6036_),
    .B(_6029_),
    .Y(_6037_)
);

NAND3X1 _16004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5542_),
    .B(_5577_),
    .C(_5572_),
    .Y(_5578_)
);

AND2X2 _17629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_18_bF$buf2),
    .Y(_7358_)
);

AOI21X1 _17209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6891_),
    .B(_6892_),
    .C(_6890_),
    .Y(_6898_)
);

NOR2X1 _12764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10035_),
    .B(_11712_),
    .Y(_11723_)
);

OR2X2 _12344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5903_),
    .B(_5892_),
    .Y(_7120_)
);

NAND3X1 _22862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1060_),
    .B(_1178_),
    .C(_1174_),
    .Y(_1186_)
);

OAI21X1 _22442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .B(_503_),
    .C(_537_),
    .Y(_726_)
);

NAND3X1 _22022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_265_),
    .C(_262_),
    .Y(_266_)
);

AOI21X1 _13969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3120_),
    .B(_3122_),
    .C(_3123_),
    .Y(_3348_)
);

OAI21X1 _13549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2888_),
    .B(_2887_),
    .C(_2878_),
    .Y(_2889_)
);

OAI21X1 _13129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2012_),
    .B(_2427_),
    .C(_2428_),
    .Y(_2429_)
);

NAND2X1 _23647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2039_),
    .B(_2027_),
    .Y(_2041_)
);

NOR2X1 _23227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686__bF$buf1),
    .B(_5676_),
    .Y(_1582_)
);

AOI21X1 _14910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4377_),
    .B(_4376_),
    .C(_4375_),
    .Y(_4378_)
);

AOI21X1 _17382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7073_),
    .B(_7077_),
    .C(_7078_),
    .Y(_7089_)
);

NOR3X1 _18587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7985_),
    .B(_7990_),
    .C(_7993_),
    .Y(_8409_)
);

NAND3X1 _18167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7930_),
    .B(_7944_),
    .C(_7948_),
    .Y(_7949_)
);

OAI21X1 _21713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11829_),
    .B(_11828_),
    .C(_11541_),
    .Y(_11836_)
);

NAND3X1 _14087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3458_),
    .B(_3465_),
    .C(_3468_),
    .Y(_3478_)
);

NAND3X1 _22918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1099_),
    .B(_1241_),
    .C(_1242_),
    .Y(_1247_)
);

NAND3X1 _16653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .B(_6278_),
    .C(_6280_),
    .Y(_6289_)
);

FILL SFILL13960x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _16233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5825_),
    .B(_5827_),
    .C(_5828_),
    .Y(_5829_)
);

FILL SFILL74200x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7609_),
    .B(_7607_),
    .C(_7608_),
    .Y(_7610_)
);

NOR3X1 _17438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6724_),
    .B(_6726_),
    .C(_6723_),
    .Y(_7150_)
);

NOR2X1 _17018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6683_),
    .B(_6684_),
    .Y(_6689_)
);

OAI21X1 _12993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_2287__bF$buf3),
    .C(_582_),
    .Y(_2288_)
);

NAND3X1 _12573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8511_),
    .B(_9609_),
    .C(_9620_),
    .Y(_9631_)
);

INVX2 _12153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5014_),
    .Y(_5025_)
);

NAND2X1 _22671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(_970_),
    .Y(_977_)
);

OR2X2 _22251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_512_),
    .Y(_517_)
);

FILL SFILL64280x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3134_),
    .B(_3138_),
    .Y(_3139_)
);

XNOR2X1 _13358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2653_),
    .Y(_2680_)
);

NAND2X1 _23876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2285_),
    .B(_2283_),
    .Y(_0_[63])
);

OAI21X1 _23456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(_1831_),
    .C(_1830_),
    .Y(_1833_)
);

AOI21X1 _23036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1370_),
    .B(_1374_),
    .C(_1267_),
    .Y(_1375_)
);

NAND3X1 _17191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6876_),
    .B(_6877_),
    .C(_6875_),
    .Y(_6879_)
);

FILL SFILL33720x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5488_),
    .B(_5489_),
    .C(_5487_),
    .Y(_5490_)
);

AOI21X1 _15504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5028_),
    .B(_5027_),
    .C(_5026_),
    .Y(_5029_)
);

AND2X2 _18396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_8200_)
);

NOR3X1 _16709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5957_),
    .B(_5959_),
    .C(_5956_),
    .Y(_6350_)
);

OAI22X1 _21942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11229_),
    .B(_8773_),
    .C(_2379_),
    .D(_8759_),
    .Y(_179_)
);

OAI21X1 _21522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf4),
    .B(_6050__bF$buf3),
    .C(_11615_),
    .Y(_11627_)
);

NOR2X1 _21102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11166_),
    .B(_11160_),
    .Y(_11167_)
);

FILL SFILL13560x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10233_),
    .B(_10068_),
    .C(_10189_),
    .Y(_10244_)
);

AND2X2 _12209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5596_),
    .B(_5629_),
    .Y(_5640_)
);

NAND2X1 _22727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_27_bF$buf5),
    .Y(_1038_)
);

OAI21X1 _22307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_576_),
    .C(_577_),
    .Y(_578_)
);

INVX2 _16882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6513_),
    .Y(_6540_)
);

OAI21X1 _16462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf3),
    .B(_3781__bF$buf0),
    .C(_5688_),
    .Y(_6078_)
);

NAND3X1 _16042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5617_),
    .B(_5619_),
    .C(_5616_),
    .Y(_5620_)
);

OAI21X1 _17667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7396_),
    .B(_7397_),
    .C(_7399_),
    .Y(_7400_)
);

NOR3X1 _17247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6934_),
    .B(_6936_),
    .C(_6939_),
    .Y(_6940_)
);

NAND3X1 _12382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7503_),
    .B(_7514_),
    .C(_7525_),
    .Y(_7536_)
);

NAND3X1 _22480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_760_),
    .C(_737_),
    .Y(_767_)
);

OR2X2 _22060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_303_),
    .Y(_307_)
);

FILL SFILL13720x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2921_),
    .C(_2841_),
    .Y(_2931_)
);

NOR3X1 _13167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_2462_),
    .C(_2468_),
    .Y(_2471_)
);

XNOR2X1 _23685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2067_),
    .B(_2081_),
    .Y(_2082_)
);

INVX1 _23265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1621_),
    .Y(_1625_)
);

NAND2X1 _19813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9748_),
    .B(_9753_),
    .Y(_9754_)
);

FILL SFILL74280x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5275_),
    .B(_5276_),
    .C(_5272_),
    .Y(_5281_)
);

AND2X2 _15313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_18_bF$buf4),
    .Y(_4821_)
);

BUFX2 BUFX2_insert50 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf1)
);

BUFX2 BUFX2_insert51 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf0)
);

BUFX2 BUFX2_insert52 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf5)
);

BUFX2 BUFX2_insert53 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf4)
);

BUFX2 BUFX2_insert54 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf3)
);

BUFX2 BUFX2_insert55 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf2)
);

BUFX2 BUFX2_insert56 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf1)
);

BUFX2 BUFX2_insert57 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[28]),
    .Y(breg_28_bF$buf0)
);

BUFX2 BUFX2_insert58 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf4)
);

BUFX2 BUFX2_insert59 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf3)
);

AOI21X1 _16938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6342_),
    .B(_6348_),
    .C(_6265_),
    .Y(_6601_)
);

NOR2X1 _16518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5768_),
    .B(_6139_),
    .Y(_6140_)
);

INVX1 _21751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11875_),
    .Y(_11877_)
);

OAI21X1 _21331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11416_),
    .B(_11415_),
    .C(_11412_),
    .Y(_11418_)
);

FILL SFILL64280x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_823_),
    .B(_834_),
    .C(_812_),
    .Y(_845_)
);

AOI21X1 _12438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8095_),
    .B(_8106_),
    .C(_7272_),
    .Y(_8150_)
);

NAND2X1 _22956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1286_),
    .B(_1287_),
    .Y(_1288_)
);

XNOR2X1 _12018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3536_),
    .B(_3503_),
    .Y(_3547_)
);

INVX1 _22536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .Y(_829_)
);

NAND2X1 _22116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf2),
    .B(areg_24_bF$buf0),
    .Y(_368_)
);

FILL SFILL64200x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6305_),
    .B(_6302_),
    .Y(_6331_)
);

NAND3X1 _16271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5868_),
    .B(_5869_),
    .C(_5867_),
    .Y(_5871_)
);

AOI21X1 _17896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7650_),
    .B(_4648_),
    .C(_7649_),
    .Y(_7651_)
);

NAND3X1 _17476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7183_),
    .B(_7190_),
    .C(_6813_),
    .Y(_7191_)
);

NAND2X1 _17056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6729_),
    .B(_6730_),
    .Y(_6731_)
);

NAND2X1 _12191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_7_bF$buf5),
    .Y(_5442_)
);

NAND3X1 _20602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10602_),
    .B(_10607_),
    .C(_10614_),
    .Y(_10619_)
);

FILL SFILL54200x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2721_),
    .B(_2556_),
    .C(_2718_),
    .Y(_2722_)
);

INVX1 _23494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .Y(_1874_)
);

NAND2X1 _23074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf4),
    .B(breg_27_bF$buf1),
    .Y(_1416_)
);

NAND3X1 _19622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9531_),
    .B(_9544_),
    .C(_9539_),
    .Y(_9545_)
);

AOI21X1 _19202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8695_),
    .B(_8729_),
    .C(_8738_),
    .Y(_9083_)
);

NAND2X1 _21807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf1),
    .B(breg_25_bF$buf2),
    .Y(_30_)
);

AOI21X1 _15962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5521_),
    .B(_5520_),
    .C(_5516_),
    .Y(_5532_)
);

OAI21X1 _15542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5068_),
    .B(_5070_),
    .C(_5067_),
    .Y(_5071_)
);

OAI21X1 _15122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4609_),
    .B(_4611_),
    .C(_4608_),
    .Y(_4612_)
);

FILL SFILL48920x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10161_),
    .B(_10162_),
    .C(_10159_),
    .Y(_10176_)
);

NAND3X1 _16747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6391_),
    .B(_6047_),
    .C(_6384_),
    .Y(_6392_)
);

AND2X2 _16327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_27_bF$buf3),
    .Y(_5932_)
);

AOI21X1 _21980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11600_),
    .B(_11847_),
    .C(_219_),
    .Y(_220_)
);

NOR2X1 _21560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11135_),
    .B(_11661_),
    .Y(_11667_)
);

NAND3X1 _21140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11192_),
    .B(_11196_),
    .C(_11199_),
    .Y(_11208_)
);

FILL SFILL13720x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10496_),
    .B(_10540_),
    .C(_10617_),
    .Y(_10661_)
);

NOR2X1 _12247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf3),
    .B(_6044__bF$buf5),
    .Y(_6055_)
);

OAI21X1 _22765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1079_),
    .B(_1074_),
    .C(_948_),
    .Y(_1080_)
);

NOR2X1 _22345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_6686__bF$buf0),
    .Y(_620_)
);

INVX1 _16080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5659_),
    .Y(_5660_)
);

NAND3X1 _14813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4233_),
    .B(_4266_),
    .C(_4272_),
    .Y(_4273_)
);

AOI21X1 _17285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6605_),
    .B(_6607_),
    .C(_6981_),
    .Y(_6982_)
);

NOR3X1 _20831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10853_),
    .B(_10862_),
    .C(_10863_),
    .Y(_10870_)
);

OAI22X1 _20411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9759_),
    .B(_10406_),
    .C(_10407_),
    .D(_10111_),
    .Y(_10409_)
);

FILL SFILL38840x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _19851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9794_),
    .Y(_9796_)
);

OAI22X1 _19431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8605_),
    .B(_9333_),
    .C(_9008_),
    .D(_9011_),
    .Y(_9335_)
);

NAND3X1 _19011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8872_),
    .B(_8873_),
    .C(_8871_),
    .Y(_8875_)
);

OAI22X1 _11938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_2661_),
    .C(_2650_),
    .D(_2376__bF$buf0),
    .Y(_2672_)
);

NAND2X1 _21616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_25_bF$buf2),
    .Y(_11729_)
);

FILL SFILL28840x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3480x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5309_),
    .B(_5319_),
    .C(_5320_),
    .Y(_5322_)
);

NAND2X1 _15351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_4863_)
);

OAI21X1 _16976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6642_),
    .B(_6638_),
    .C(_6603_),
    .Y(_6643_)
);

AOI21X1 _16556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6171_),
    .B(_6170_),
    .C(_6167_),
    .Y(_6182_)
);

AOI21X1 _16136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5714_),
    .B(_5715_),
    .C(_5713_),
    .Y(_5722_)
);

FILL SFILL18840x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9915_),
    .B(_9904_),
    .C(_8402_),
    .Y(_1260_)
);

NOR2X1 _12476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf3),
    .B(_8555_),
    .Y(_8566_)
);

OAI21X1 _22994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1327_),
    .B(_1328_),
    .C(_1326_),
    .Y(_1329_)
);

INVX1 _12056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3953_),
    .Y(_3964_)
);

NAND2X1 _22574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .B(_865_),
    .Y(_871_)
);

INVX1 _22154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .Y(_411_)
);

AND2X2 _18702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8531_),
    .B(_8532_),
    .Y(_8535_)
);

XNOR2X1 _23779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .B(_2182_),
    .Y(_2183_)
);

NAND3X1 _23359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1722_),
    .B(_1726_),
    .C(_1664_),
    .Y(_1727_)
);

NAND2X1 _19907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_23_bF$buf1),
    .Y(_9857_)
);

XOR2X1 _14622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4062_),
    .B(_4060_),
    .Y(_4063_)
);

OAI21X1 _14202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf1),
    .B(_7217__bF$buf0),
    .C(_3602_),
    .Y(_3603_)
);

OAI21X1 _17094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6498_),
    .B(_6502_),
    .C(_6504_),
    .Y(_6773_)
);

FILL SFILL48920x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_18_bF$buf0),
    .Y(_5383_)
);

NOR3X1 _15407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4595_),
    .B(_4596_),
    .C(_4594_),
    .Y(_4924_)
);

NAND2X1 _20640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10659_),
    .B(_10654_),
    .Y(_10660_)
);

OAI21X1 _20220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10198_),
    .B(_10193_),
    .C(_10110_),
    .Y(_10199_)
);

NAND3X1 _18299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8088_),
    .B(_8092_),
    .C(_8091_),
    .Y(_8093_)
);

AOI21X1 _19660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9210_),
    .B(_9208_),
    .C(_9585_),
    .Y(_9586_)
);

NAND3X1 _19240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9120_),
    .B(_9105_),
    .C(_9121_),
    .Y(_9125_)
);

AOI21X1 _21845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_65_),
    .C(_64_),
    .Y(_72_)
);

OAI21X1 _21425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11507_),
    .B(_11511_),
    .C(_11251_),
    .Y(_11521_)
);

OAI21X1 _21005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10749_),
    .B(_10744_),
    .C(_10752_),
    .Y(_11060_)
);

AND2X2 _15580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_15_bF$buf4),
    .Y(_5112_)
);

NAND2X1 _15160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4356_),
    .B(_4358_),
    .Y(_4652_)
);

FILL SFILL38920x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _16785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6432_),
    .B(_6429_),
    .Y(_6433_)
);

OAI21X1 _16365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5972_),
    .B(_5973_),
    .C(_5971_),
    .Y(_5974_)
);

FILL SFILL3560x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert490 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(breg_2_bF$buf0)
);

BUFX2 BUFX2_insert491 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .Y(_6686__bF$buf3)
);

BUFX2 BUFX2_insert492 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .Y(_6686__bF$buf2)
);

BUFX2 BUFX2_insert493 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .Y(_6686__bF$buf1)
);

BUFX2 BUFX2_insert494 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686_),
    .Y(_6686__bF$buf0)
);

BUFX2 BUFX2_insert495 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf4)
);

BUFX2 BUFX2_insert496 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf3)
);

BUFX2 BUFX2_insert497 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf2)
);

FILL SFILL69240x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert498 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf1)
);

BUFX2 BUFX2_insert499 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(breg_11_bF$buf0)
);

FILL SFILL43960x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_4434__bF$buf2),
    .Y(_6472_)
);

NAND3X1 _22383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_655_),
    .B(_661_),
    .C(_608_),
    .Y(_662_)
);

FILL SFILL28920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8770_),
    .B(_7968_),
    .C(_8781_),
    .Y(_8787_)
);

AOI21X1 _18511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8319_),
    .B(_8320_),
    .C(_8322_),
    .Y(_8327_)
);

FILL SFILL3880x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28840x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _23588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(_725_),
    .Y(_1976_)
);

NOR3X1 _23168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1517_),
    .B(_1516_),
    .C(_1518_),
    .Y(_1519_)
);

INVX1 _19716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9646_),
    .Y(_9647_)
);

OAI21X1 _14851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4312_),
    .B(_4313_),
    .C(_4311_),
    .Y(_4315_)
);

NAND3X1 _14431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3852_),
    .B(_3853_),
    .C(_3848_),
    .Y(_3855_)
);

XNOR2X1 _14011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3393_),
    .B(_3388_),
    .Y(_3395_)
);

AND2X2 _15636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4824_),
    .B(_4822_),
    .Y(_5174_)
);

AND2X2 _15216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_16_bF$buf2),
    .Y(_4714_)
);

FILL SFILL18840x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3077_),
    .B(_3066_),
    .Y(_3088_)
);

INVX1 _21654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11757_),
    .Y(_11771_)
);

OAI21X1 _21234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11001_),
    .B(_10994_),
    .C(_11310_),
    .Y(_11311_)
);

OAI21X1 _22859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1181_),
    .B(_1180_),
    .C(_1060_),
    .Y(_1182_)
);

OAI21X1 _22439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_721_),
    .B(_718_),
    .C(_711_),
    .Y(_722_)
);

NAND2X1 _22019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_261_),
    .Y(_262_)
);

NOR2X1 _13702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3054_),
    .B(_3056_),
    .Y(_3057_)
);

NAND3X1 _23800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(_2202_),
    .C(_2205_),
    .Y(_2206_)
);

XOR2X1 _16594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5842_),
    .B(_6223_),
    .Y(_6224_)
);

AOI21X1 _16174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5763_),
    .B(_5762_),
    .C(_5761_),
    .Y(_5764_)
);

INVX2 _14907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4370_),
    .Y(_4375_)
);

OAI21X1 _17799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7544_),
    .B(_7543_),
    .C(_7542_),
    .Y(_7545_)
);

INVX1 _17379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6655_),
    .Y(_7085_)
);

NOR2X1 _12094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf1),
    .B(_2508_),
    .Y(_4379_)
);

AOI21X1 _22192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_363_),
    .C(_361_),
    .Y(_453_)
);

OAI21X1 _18740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8562_),
    .B(_8561_),
    .C(_8559_),
    .Y(_8576_)
);

OAI21X1 _18320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8115_),
    .B(_8111_),
    .C(_8081_),
    .Y(_8116_)
);

NOR3X1 _20925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10609_),
    .B(_10615_),
    .C(_10618_),
    .Y(_10973_)
);

AND2X2 _20505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10157_),
    .B(_10212_),
    .Y(_10512_)
);

AOI21X1 _13299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2600_),
    .B(_2603_),
    .C(_2590_),
    .Y(_2614_)
);

XNOR2X1 _23397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1656_),
    .B(_1768_),
    .Y(_0_[53])
);

NAND3X1 _19945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9894_),
    .B(_9884_),
    .C(_9889_),
    .Y(_9898_)
);

NAND3X1 _19525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9428_),
    .B(_9436_),
    .C(_9437_),
    .Y(_9438_)
);

OAI21X1 _19105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8969_),
    .B(_8968_),
    .C(_8966_),
    .Y(_8977_)
);

FILL SFILL59080x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf2),
    .B(_2362__bF$buf0),
    .C(_3817_),
    .Y(_4104_)
);

NAND2X1 _14240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3643_),
    .B(_3644_),
    .Y(_3645_)
);

FILL SFILL38920x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5414_),
    .B(_5413_),
    .C(_5410_),
    .Y(_5425_)
);

NOR3X1 _15445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4954_),
    .B(_4955_),
    .C(_4951_),
    .Y(_4964_)
);

NAND2X1 _15025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4503_),
    .B(_4504_),
    .Y(_4505_)
);

FILL SFILL3560x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_113_),
    .B(_112_),
    .C(_109_),
    .Y(_114_)
);

AOI21X1 _21463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11541_),
    .B(_11544_),
    .C(_11546_),
    .Y(_11563_)
);

OAI21X1 _21043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11100_),
    .B(_11101_),
    .C(_11098_),
    .Y(_11102_)
);

FILL SFILL28920x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_972_),
    .Y(_973_)
);

AND2X2 _22248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_267_),
    .B(_512_),
    .Y(_513_)
);

NAND3X1 _13931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3249_),
    .B(_3305_),
    .C(_3306_),
    .Y(_3308_)
);

NAND2X1 _13511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2844_),
    .B(_2846_),
    .Y(_2848_)
);

FILL SFILL39080x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf5),
    .B(areg_12_bF$buf0),
    .Y(_4166_)
);

INVX1 _17188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6850_),
    .Y(_6875_)
);

FILL SFILL18760x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf3),
    .B(_3781__bF$buf1),
    .C(_10406_),
    .Y(_10763_)
);

AOI21X1 _20314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10283_),
    .B(_10290_),
    .C(_10108_),
    .Y(_10303_)
);

NAND2X1 _19754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9336_),
    .B(_9342_),
    .Y(_9689_)
);

AOI21X1 _19334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8842_),
    .B(_8844_),
    .C(_9228_),
    .Y(_9229_)
);

NAND3X1 _21939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_173_),
    .C(_174_),
    .Y(_175_)
);

OAI21X1 _21519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11622_),
    .B(_11621_),
    .C(_11611_),
    .Y(_11623_)
);

NAND3X1 _15674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5213_),
    .B(_5215_),
    .C(_5214_),
    .Y(_5216_)
);

AOI21X1 _15254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4739_),
    .B(_4746_),
    .C(_4709_),
    .Y(_4756_)
);

OAI21X1 _16879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6535_),
    .B(_6534_),
    .C(_6520_),
    .Y(_6536_)
);

AOI21X1 _16459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6067_),
    .B(_6068_),
    .C(_6060_),
    .Y(_6074_)
);

NAND2X1 _16039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5614_),
    .B(_5615_),
    .Y(_5616_)
);

NAND2X1 _21692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_31_bF$buf3),
    .Y(_11813_)
);

NOR3X1 _21272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11351_),
    .B(_11346_),
    .C(_11349_),
    .Y(_11352_)
);

AOI21X1 _17820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7091_),
    .B(_7140_),
    .C(_7567_),
    .Y(_7568_)
);

NAND2X1 _17400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf4),
    .B(areg_28_bF$buf3),
    .Y(_7108_)
);

OAI21X1 _12799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10463_),
    .B(_177_),
    .C(_188_),
    .Y(_199_)
);

OR2X2 _12379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6253_),
    .B(_7305_),
    .Y(_7503_)
);

OAI21X1 _22897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .B(_1222_),
    .C(_1223_),
    .Y(_1224_)
);

AOI21X1 _22477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_762_),
    .B(_763_),
    .C(_736_),
    .Y(_764_)
);

FILL SFILL3560x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _22057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_302_),
    .B(_303_),
    .Y(_304_)
);

AOI21X1 _18605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8422_),
    .B(_8428_),
    .C(_8185_),
    .Y(_8429_)
);

FILL SFILL59080x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3097_),
    .B(_2859_),
    .Y(_3098_)
);

NAND2X1 _13320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf3),
    .B(areg_10_bF$buf4),
    .Y(_2638_)
);

FILL SFILL3640x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4399_),
    .B(_4404_),
    .C(_4408_),
    .Y(_4417_)
);

INVX8 _14525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf2),
    .Y(_3958_)
);

NAND2X1 _14105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(_3491_),
    .Y(_3498_)
);

OAI21X1 _20963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10811_),
    .B(_11013_),
    .C(_10969_),
    .Y(_11014_)
);

OAI21X1 _20543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10552_),
    .B(_10553_),
    .C(_10550_),
    .Y(_10554_)
);

OAI21X1 _20123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10087_),
    .B(_10088_),
    .C(_10042_),
    .Y(_10093_)
);

AOI21X1 _19983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9582_),
    .B(_9580_),
    .C(_9939_),
    .Y(_9940_)
);

OAI21X1 _19563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9479_),
    .B(_9478_),
    .C(_9476_),
    .Y(_9480_)
);

AND2X2 _19143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf3),
    .B(breg_18_bF$buf1),
    .Y(_9019_)
);

FILL SFILL33880x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11868_),
    .B(_11867_),
    .C(_11872_),
    .Y(_11873_)
);

OAI21X1 _21328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11402_),
    .B(_11401_),
    .C(_11399_),
    .Y(_11414_)
);

NAND3X1 _15483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4669_),
    .B(_5005_),
    .C(_5004_),
    .Y(_5006_)
);

NOR2X1 _15063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4245_),
    .B(_4539_),
    .Y(_4547_)
);

AOI21X1 _16688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6315_),
    .B(_6313_),
    .C(_6310_),
    .Y(_6327_)
);

XNOR2X1 _16268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5844_),
    .B(_5840_),
    .Y(_5867_)
);

AND2X2 _21081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_22_bF$buf1),
    .Y(_11144_)
);

FILL SFILL39000x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5387_),
    .B(_5398_),
    .C(_5354_),
    .Y(_5409_)
);

OAI21X1 _22286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf1),
    .B(_5676_),
    .C(_554_),
    .Y(_555_)
);

AOI21X1 _18834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8283_),
    .B(_8318_),
    .C(_8328_),
    .Y(_8680_)
);

OAI21X1 _18414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8202_),
    .B(_8207_),
    .C(_8209_),
    .Y(_8220_)
);

FILL SFILL29080x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_30_bF$buf3),
    .Y(_9541_)
);

INVX1 _14754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4207_),
    .Y(_4208_)
);

AOI21X1 _14334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3743_),
    .B(_3748_),
    .C(_3521_),
    .Y(_3749_)
);

DFFPOSX1 _24012_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[2]),
    .CLK(clk_bF$buf0),
    .D(a[2])
);

FILL SFILL29000x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5527_),
    .Y(_5528_)
);

AOI21X1 _15539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4395_),
    .B(_5046_),
    .C(_4727_),
    .Y(_5067_)
);

AOI21X1 _15119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4300_),
    .B(_4152_),
    .C(_4607_),
    .Y(_4608_)
);

OAI21X1 _20772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10802_),
    .B(_10801_),
    .C(_10804_),
    .Y(_10805_)
);

OAI21X1 _20352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10343_),
    .B(_10306_),
    .C(_10298_),
    .Y(_10344_)
);

NAND3X1 _16900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6550_),
    .B(_6557_),
    .C(_6558_),
    .Y(_6559_)
);

NAND3X1 _19792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9711_),
    .B(_9715_),
    .C(_9721_),
    .Y(_9731_)
);

INVX2 _19372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9269_),
    .Y(_9270_)
);

AOI21X1 _21977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_216_),
    .C(_11885_),
    .Y(_217_)
);

NAND3X1 _21557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11655_),
    .B(_11660_),
    .C(_11663_),
    .Y(_11664_)
);

NAND3X1 _21137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11197_),
    .B(_11204_),
    .C(_11167_),
    .Y(_11205_)
);

FILL SFILL43960x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_10_bF$buf4),
    .Y(_429_)
);

NAND3X1 _12400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7678_),
    .B(_7722_),
    .C(_7700_),
    .Y(_7733_)
);

NAND3X1 _15292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4789_),
    .B(_4782_),
    .C(_4787_),
    .Y(_4798_)
);

FILL SFILL43880x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2934_),
    .B(_2940_),
    .C(_2790_),
    .Y(_2951_)
);

XOR2X1 _23703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2101_),
    .B(_2058_),
    .Y(_2102_)
);

AOI21X1 _16497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6112_),
    .B(_6113_),
    .C(_6053_),
    .Y(_6117_)
);

NAND2X1 _16077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5654_),
    .B(_5657_),
    .Y(_5658_)
);

AOI21X1 _22095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_334_),
    .B(_327_),
    .C(_296_),
    .Y(_346_)
);

AOI22X1 _18643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8458_),
    .B(_8462_),
    .C(_8058_),
    .D(_8066_),
    .Y(_8470_)
);

NAND3X1 _18223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8009_),
    .B(_8010_),
    .C(_8007_),
    .Y(_8011_)
);

FILL SFILL33880x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54360x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10511_),
    .B(_10558_),
    .Y(_10866_)
);

NAND3X1 _20408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10402_),
    .B(_10404_),
    .C(_10403_),
    .Y(_10405_)
);

AND2X2 _19848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_21_bF$buf3),
    .Y(_9792_)
);

OAI21X1 _19428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf1),
    .B(_5315__bF$buf4),
    .C(_9324_),
    .Y(_9331_)
);

AOI21X1 _19008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8071_),
    .B(_8455_),
    .C(_8870_),
    .Y(_8871_)
);

AND2X2 _14983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_14_bF$buf0),
    .Y(_4458_)
);

AOI21X1 _14563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3710_),
    .B(_3713_),
    .C(_3999_),
    .Y(_4000_)
);

OAI21X1 _14143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2993_),
    .B(_3266_),
    .C(_3265_),
    .Y(_3539_)
);

INVX4 _15768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .Y(_5318_)
);

AOI22X1 _15348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_24_bF$buf4),
    .C(breg_1_bF$buf4),
    .D(areg_23_bF$buf3),
    .Y(_4859_)
);

NOR2X1 _20581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10257_),
    .B(_9535_),
    .Y(_10596_)
);

FILL SFILL23880x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10131_),
    .B(_10132_),
    .C(_10133_),
    .Y(_10135_)
);

FILL SFILL39000x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8657_),
    .B(_8699_),
    .Y(_9061_)
);

AOI21X1 _21786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11903_),
    .B(_11901_),
    .C(_11897_),
    .Y(_7_)
);

FILL SFILL23800x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11451_),
    .B(_11452_),
    .Y(_11456_)
);

OAI21X1 _17914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7245_),
    .B(_7235_),
    .C(_7240_),
    .Y(_7671_)
);

FILL SFILL8840x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3200_),
    .B(_3201_),
    .C(_3095_),
    .Y(_3202_)
);

NAND3X1 _13414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2729_),
    .B(_2732_),
    .C(_2735_),
    .Y(_2742_)
);

BUFX2 _23932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[50]),
    .Y(y[50])
);

OAI21X1 _23512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf0),
    .B(_7225__bF$buf2),
    .C(_1892_),
    .Y(_1893_)
);

FILL SFILL29000x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4029_),
    .B(_3778_),
    .C(_4033_),
    .Y(_4059_)
);

NAND3X1 _18872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8715_),
    .B(_8716_),
    .C(_8721_),
    .Y(_8722_)
);

AOI21X1 _18452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8254_),
    .B(_8261_),
    .C(_8222_),
    .Y(_8262_)
);

NAND3X1 _18032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7795_),
    .B(_7800_),
    .C(_7798_),
    .Y(_7801_)
);

NAND3X1 _20637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10340_),
    .B(_10652_),
    .C(_10651_),
    .Y(_10657_)
);

NOR3X1 _20217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9893_),
    .B(_9894_),
    .C(_9892_),
    .Y(_10196_)
);

FILL SFILL43960x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9582_),
    .B(_9581_),
    .C(_9580_),
    .Y(_9583_)
);

NAND3X1 _19237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9119_),
    .B(_9120_),
    .C(_9121_),
    .Y(_9122_)
);

NAND3X1 _14792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4244_),
    .B(_4248_),
    .C(_4246_),
    .Y(_4249_)
);

NAND2X1 _14372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf4),
    .B(breg_18_bF$buf5),
    .Y(_3790_)
);

DFFPOSX1 _24050_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[8]),
    .CLK(clk_bF$buf8),
    .D(b[8])
);

AOI21X1 _15997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5561_),
    .B(_5559_),
    .C(_5557_),
    .Y(_5570_)
);

OAI21X1 _15577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4786_),
    .B(_4776_),
    .C(_4780_),
    .Y(_5109_)
);

NOR3X1 _15157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4633_),
    .B(_4634_),
    .C(_4631_),
    .Y(_4649_)
);

NOR3X1 _20390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10382_),
    .B(_10383_),
    .C(_10384_),
    .Y(_10385_)
);

AOI21X1 _21595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11519_),
    .B(_11521_),
    .C(_11512_),
    .Y(_11706_)
);

NOR2X1 _21175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11235_),
    .B(_11246_),
    .Y(_11247_)
);

AOI21X1 _17723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7450_),
    .B(_7449_),
    .C(_7445_),
    .Y(_7462_)
);

NAND3X1 _17303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7000_),
    .B(_6998_),
    .C(_7001_),
    .Y(_7002_)
);

AOI22X1 _18928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8778_),
    .B(_8782_),
    .C(_8769_),
    .D(_8763_),
    .Y(_8783_)
);

NAND3X1 _18508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8322_),
    .B(_8319_),
    .C(_8320_),
    .Y(_8323_)
);

NOR2X1 _13643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2763_),
    .Y(_2992_)
);

OAI21X1 _13223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2351_),
    .B(_2346_),
    .C(_2341_),
    .Y(_2533_)
);

XNOR2X1 _23741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2137_),
    .Y(_2143_)
);

NOR2X1 _23321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1684_),
    .B(_1671_),
    .Y(_1686_)
);

FILL SFILL8920x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4021_),
    .B(_4023_),
    .C(_4310_),
    .Y(_4311_)
);

NAND3X1 _14428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3833_),
    .B(_3837_),
    .C(_3841_),
    .Y(_3851_)
);

INVX2 _14008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3390_),
    .Y(_3391_)
);

FILL SFILL23880x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8507_),
    .B(_8508_),
    .C(_8504_),
    .Y(_8512_)
);

NAND3X1 _18261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8047_),
    .B(_8048_),
    .C(_8051_),
    .Y(_8053_)
);

FILL SFILL23800x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10905_),
    .B(_10906_),
    .C(_10907_),
    .Y(_10908_)
);

NAND3X1 _20446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10444_),
    .B(_10445_),
    .C(_10446_),
    .Y(_10447_)
);

OAI21X1 _20026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9983_),
    .B(_9984_),
    .C(_9985_),
    .Y(_9986_)
);

AOI21X1 _19886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9782_),
    .B(_9778_),
    .C(_9764_),
    .Y(_9834_)
);

NAND3X1 _19466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9354_),
    .B(_9359_),
    .C(_9363_),
    .Y(_9373_)
);

AOI21X1 _19046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8492_),
    .B(_8496_),
    .C(_8499_),
    .Y(_8912_)
);

AOI21X1 _14181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3566_),
    .B(_3571_),
    .C(_3537_),
    .Y(_3581_)
);

FILL SFILL13880x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1445_),
    .B(_11723_),
    .Y(_1456_)
);

OAI21X1 _15386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4805_),
    .B(_4801_),
    .C(_4808_),
    .Y(_4901_)
);

FILL SFILL13800x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert110 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434_),
    .Y(_4434__bF$buf0)
);

BUFX2 BUFX2_insert111 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .Y(_3781__bF$buf3)
);

BUFX2 BUFX2_insert112 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .Y(_3781__bF$buf2)
);

BUFX2 BUFX2_insert113 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .Y(_3781__bF$buf1)
);

NAND2X1 _17952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_24_bF$buf4),
    .Y(_7713_)
);

BUFX2 BUFX2_insert114 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781_),
    .Y(_3781__bF$buf0)
);

AOI21X1 _17532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7249_),
    .B(_7251_),
    .C(_7235_),
    .Y(_7252_)
);

BUFX2 BUFX2_insert115 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf5)
);

BUFX2 BUFX2_insert116 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf4)
);

NAND3X1 _17112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6787_),
    .B(_6420_),
    .C(_6792_),
    .Y(_6793_)
);

BUFX2 BUFX2_insert117 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf3)
);

BUFX2 BUFX2_insert118 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf2)
);

BUFX2 BUFX2_insert119 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[16]),
    .Y(breg_16_bF$buf1)
);

FILL SFILL23640x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _22189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_364_),
    .C(_448_),
    .D(_447_),
    .Y(_449_)
);

NOR3X1 _18737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8153_),
    .B(_8152_),
    .C(_8154_),
    .Y(_8573_)
);

AOI21X1 _18317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8108_),
    .B(_8109_),
    .C(_8083_),
    .Y(_8113_)
);

NOR3X1 _13872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3218_),
    .B(_3222_),
    .C(_3225_),
    .Y(_3243_)
);

AOI21X1 _13452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2619_),
    .C(_2622_),
    .Y(_2783_)
);

DFFPOSX1 _23970_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[24]),
    .CLK(clk_bF$buf7),
    .D(_0_[24])
);

NAND3X1 _13032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2326_),
    .C(_1478_),
    .Y(_2327_)
);

INVX1 _23550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1929_),
    .Y(_1935_)
);

NAND3X1 _23130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1470_),
    .B(_1476_),
    .C(_1436_),
    .Y(_1477_)
);

FILL SFILL64040x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_16_bF$buf2),
    .Y(_4101_)
);

NOR2X1 _14237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf1),
    .B(_10869__bF$buf3),
    .Y(_3642_)
);

NAND3X1 _18490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8297_),
    .B(_8299_),
    .C(_8298_),
    .Y(_8303_)
);

AOI21X1 _18070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7835_),
    .B(_7841_),
    .C(_7819_),
    .Y(_7842_)
);

NAND2X1 _20675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10435_),
    .B(_10443_),
    .Y(_10698_)
);

NAND3X1 _20255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10229_),
    .B(_10237_),
    .C(_10214_),
    .Y(_10238_)
);

OAI21X1 _16803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf0),
    .B(_5315__bF$buf3),
    .C(_6446_),
    .Y(_6453_)
);

AOI21X1 _19695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8882_),
    .B(_9246_),
    .C(_9624_),
    .Y(_9625_)
);

FILL SFILL54040x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _19275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8364_),
    .B(_8772_),
    .C(_9163_),
    .D(_8771_),
    .Y(_9164_)
);

FILL SFILL59240x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10430_),
    .B(_11132_),
    .C(_11176_),
    .Y(_11275_)
);

NOR3X1 _12303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6615_),
    .B(_6450_),
    .C(_6626_),
    .Y(_6670_)
);

OAI21X1 _22821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_989_),
    .B(_1139_),
    .C(_1138_),
    .Y(_1141_)
);

OAI21X1 _22401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_675_),
    .C(_677_),
    .Y(_681_)
);

INVX1 _15195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4690_),
    .Y(_4691_)
);

NAND3X1 _13928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3298_),
    .B(_3250_),
    .C(_3303_),
    .Y(_3304_)
);

NOR2X1 _13508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf2),
    .B(_6582__bF$buf3),
    .Y(_2844_)
);

OAI21X1 _23606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(_1877_),
    .C(_1891_),
    .Y(_1996_)
);

FILL SFILL44040x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7095_),
    .B(_7101_),
    .C(_7103_),
    .Y(_7504_)
);

NAND3X1 _17341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7038_),
    .B(_7042_),
    .C(_7023_),
    .Y(_7044_)
);

AOI21X1 _18966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8824_),
    .B(_8802_),
    .C(_8692_),
    .Y(_8825_)
);

NOR2X1 _18546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8364_),
    .B(_7961_),
    .Y(_8365_)
);

NOR2X1 _18126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7452_),
    .B(_7903_),
    .Y(_7904_)
);

NAND3X1 _13681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3030_),
    .B(_3032_),
    .C(_3031_),
    .Y(_3034_)
);

NAND2X1 _13261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2414_),
    .B(_2409_),
    .Y(_2574_)
);

FILL SFILL69160x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4351_),
    .B(_4317_),
    .C(_4309_),
    .Y(_4352_)
);

NAND3X1 _14466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3888_),
    .B(_3889_),
    .C(_3892_),
    .Y(_3893_)
);

AOI21X1 _14046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3423_),
    .B(_3419_),
    .C(_3386_),
    .Y(_3433_)
);

FILL SFILL28920x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28840x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10482_),
    .B(_10483_),
    .C(_10488_),
    .Y(_10489_)
);

OAI21X1 _20064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10023_),
    .B(_10025_),
    .C(_10020_),
    .Y(_10028_)
);

NAND3X1 _16612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6238_),
    .B(_6243_),
    .C(_6225_),
    .Y(_6244_)
);

NOR3X1 _19084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8937_),
    .B(_8941_),
    .C(_8942_),
    .Y(_8954_)
);

NOR2X1 _21689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11533_),
    .B(_11531_),
    .Y(_11809_)
);

OAI21X1 _21269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf4),
    .B(_5668__bF$buf5),
    .C(_11336_),
    .Y(_11348_)
);

NAND3X1 _17817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7564_),
    .B(_7562_),
    .C(_7563_),
    .Y(_7565_)
);

NAND3X1 _12952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1838_),
    .B(_1860_),
    .C(_1849_),
    .Y(_1870_)
);

NAND3X1 _12532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9038_),
    .B(_9126_),
    .C(_9170_),
    .Y(_9181_)
);

OAI21X1 _22630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9992_),
    .B(_10336_),
    .C(_930_),
    .Y(_931_)
);

OAI21X1 _12112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4555_),
    .B(_4566_),
    .C(_4544_),
    .Y(_4577_)
);

AOI21X1 _22210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_465_),
    .B(_471_),
    .C(_244_),
    .Y(_472_)
);

FILL SFILL64040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3090_),
    .B(_3094_),
    .Y(_3095_)
);

NAND2X1 _23835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2225_),
    .B(_2222_),
    .Y(_2243_)
);

NAND2X1 _13317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_12_bF$buf1),
    .Y(_2635_)
);

NOR2X1 _23415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf0),
    .B(_6815__bF$buf3),
    .Y(_1788_)
);

NAND3X1 _17990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7730_),
    .B(_7735_),
    .C(_7742_),
    .Y(_7754_)
);

OAI21X1 _17570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7289_),
    .B(_7290_),
    .C(_7292_),
    .Y(_7293_)
);

INVX1 _17150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6819_),
    .Y(_6833_)
);

FILL SFILL54120x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf1),
    .B(_3529__bF$buf4),
    .C(_8614_),
    .Y(_8615_)
);

OAI21X1 _18355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8153_),
    .B(_8152_),
    .C(_8154_),
    .Y(_8155_)
);

NAND3X1 _13490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2821_),
    .B(_2822_),
    .C(_2823_),
    .Y(_2824_)
);

NAND3X1 _13070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_14_bF$buf2),
    .C(_1522_),
    .Y(_2364_)
);

NOR2X1 _21901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11764_),
    .B(_131_),
    .Y(_134_)
);

AOI21X1 _14695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4126_),
    .B(_4133_),
    .C(_4097_),
    .Y(_4143_)
);

INVX2 _14275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3678_),
    .Y(_3684_)
);

FILL SFILL44040x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10273_),
    .B(_10272_),
    .Y(_10280_)
);

OAI21X1 _16841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6480_),
    .B(_6485_),
    .C(_6487_),
    .Y(_6495_)
);

XNOR2X1 _16421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5663_),
    .B(_6033_),
    .Y(_0_[27])
);

OAI21X1 _16001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5570_),
    .B(_5569_),
    .C(_5555_),
    .Y(_5575_)
);

NAND2X1 _21498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11426_),
    .B(_11433_),
    .Y(_11600_)
);

NAND2X1 _21078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf2),
    .B(areg_21_bF$buf0),
    .Y(_11140_)
);

NAND2X1 _17626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_18_bF$buf1),
    .Y(_7355_)
);

NAND2X1 _17206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6466_),
    .B(_6470_),
    .Y(_6895_)
);

OAI21X1 _12761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10178_),
    .B(_10035_),
    .C(_10288_),
    .Y(_11690_)
);

AOI22X1 _12341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6955_),
    .B(_6999_),
    .C(_7076_),
    .D(_4981_),
    .Y(_7087_)
);

FILL SFILL69160x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3343_),
    .B(_3339_),
    .C(_3344_),
    .Y(_3345_)
);

NAND3X1 _13546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2879_),
    .B(_2885_),
    .C(_2883_),
    .Y(_2886_)
);

NOR2X1 _13126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf3),
    .B(_5420__bF$buf0),
    .Y(_2426_)
);

NOR2X1 _23644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .B(_2036_),
    .Y(_2038_)
);

OAI21X1 _23224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315__bF$buf0),
    .B(_7520__bF$buf2),
    .C(_1443_),
    .Y(_1579_)
);

DFFPOSX1 _24009_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[63]),
    .CLK(clk_bF$buf3),
    .D(_0_[63])
);

OAI21X1 _18584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8384_),
    .B(_8390_),
    .C(_8394_),
    .Y(_8406_)
);

AOI21X1 _18164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7937_),
    .B(_7936_),
    .C(_7933_),
    .Y(_7946_)
);

FILL SFILL59160x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10796_),
    .B(_10797_),
    .C(_10795_),
    .Y(_10801_)
);

OAI21X1 _20349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10031_),
    .B(_10001_),
    .C(_10039_),
    .Y(_10340_)
);

AOI21X1 _21710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11711_),
    .B(_11713_),
    .C(_11710_),
    .Y(_11832_)
);

OAI21X1 _19789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9725_),
    .B(_9726_),
    .C(_9724_),
    .Y(_9727_)
);

AOI21X1 _19369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9241_),
    .B(_9242_),
    .C(_8886_),
    .Y(_9266_)
);

NAND3X1 _14084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3246_),
    .B(_3474_),
    .C(_3466_),
    .Y(_3475_)
);

OAI21X1 _12817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11011_),
    .B(_11043_),
    .C(_10946_),
    .Y(_396_)
);

OAI21X1 _22915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .B(_1243_),
    .C(_1098_),
    .Y(_1244_)
);

INVX2 _15289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4770_),
    .Y(_4794_)
);

OAI21X1 _16650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6281_),
    .B(_6284_),
    .C(_6267_),
    .Y(_6285_)
);

AOI21X1 _16230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5821_),
    .B(_5820_),
    .C(_5819_),
    .Y(_5825_)
);

NAND2X1 _17855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7605_),
    .B(_7606_),
    .Y(_7607_)
);

NAND3X1 _17435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7129_),
    .B(_7134_),
    .C(_7137_),
    .Y(_7147_)
);

INVX8 _17015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_26_bF$buf1),
    .Y(_6686_)
);

NAND2X1 _12990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_14_bF$buf4),
    .Y(_2280_)
);

NAND3X1 _12570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8522_),
    .B(_9587_),
    .C(_9532_),
    .Y(_9598_)
);

OAI21X1 _12150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4653_),
    .B(_4675_),
    .C(_4588_),
    .Y(_4992_)
);

NOR2X1 _13775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3111_),
    .B(_3130_),
    .Y(_3136_)
);

OAI21X1 _23873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2282_),
    .B(_2276_),
    .C(_2271_),
    .Y(_2283_)
);

AOI21X1 _13355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2670_),
    .B(_2668_),
    .C(_2664_),
    .Y(_2677_)
);

AOI21X1 _23453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1693_),
    .B(_1721_),
    .C(_1725_),
    .Y(_1830_)
);

NAND3X1 _23033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1340_),
    .C(_1344_),
    .Y(_1372_)
);

AOI21X1 _15921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5111_),
    .B(_5116_),
    .C(_5118_),
    .Y(_5487_)
);

INVX2 _15501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5020_),
    .Y(_5026_)
);

NAND2X1 _18393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_20_bF$buf0),
    .Y(_8197_)
);

OAI21X1 _20998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11051_),
    .B(_11047_),
    .C(_11017_),
    .Y(_11052_)
);

NAND3X1 _20578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10262_),
    .B(_10579_),
    .C(_10585_),
    .Y(_10592_)
);

AOI21X1 _20158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9767_),
    .B(_9771_),
    .C(_9775_),
    .Y(_10131_)
);

NAND3X1 _16706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6329_),
    .B(_6334_),
    .C(_6337_),
    .Y(_6347_)
);

AOI21X1 _19598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9513_),
    .B(_9514_),
    .C(_9512_),
    .Y(_9518_)
);

AOI21X1 _19178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9050_),
    .B(_9051_),
    .C(_9043_),
    .Y(_9057_)
);

FILL SFILL59320x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf3),
    .B(_7217__bF$buf0),
    .C(_10112_),
    .Y(_10221_)
);

NAND2X1 _12206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5574_),
    .B(_5486_),
    .Y(_5607_)
);

NOR2X1 _22724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_863_),
    .Y(_1035_)
);

AOI21X1 _22304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_569_),
    .B(_570_),
    .C(_568_),
    .Y(_575_)
);

NAND3X1 _15098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4448_),
    .B(_4492_),
    .C(_4493_),
    .Y(_4585_)
);

BUFX2 _23929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[47]),
    .Y(y[47])
);

XNOR2X1 _23509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1889_),
    .Y(_1890_)
);

FILL SFILL59240x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7387_),
    .B(_7386_),
    .C(_7383_),
    .Y(_7397_)
);

AND2X2 _17244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_19_bF$buf1),
    .Y(_6937_)
);

FILL SFILL59160x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8305_),
    .B(_8717_),
    .Y(_8718_)
);

AOI21X1 _18449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8232_),
    .B(_8235_),
    .C(_8245_),
    .Y(_8258_)
);

AND2X2 _18029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_18_bF$buf1),
    .Y(_7797_)
);

AOI21X1 _13584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2927_),
    .B(_2926_),
    .C(_2835_),
    .Y(_2928_)
);

AND2X2 _13164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2294_),
    .B(_2461_),
    .Y(_2468_)
);

NAND2X1 _23682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2078_),
    .Y(_2079_)
);

NAND3X1 _23262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1621_),
    .B(_1612_),
    .C(_1616_),
    .Y(_1622_)
);

NAND3X1 _19810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9741_),
    .B(_9746_),
    .C(_9736_),
    .Y(_9750_)
);

FILL SFILL33960x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3959_),
    .B(_4245_),
    .Y(_4246_)
);

AOI21X1 _14369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3527_),
    .B(_3530_),
    .C(_3784_),
    .Y(_3785_)
);

DFFPOSX1 _24047_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[5]),
    .CLK(clk_bF$buf1),
    .D(b[5])
);

FILL SFILL18760x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5275_),
    .B(_5276_),
    .C(_5272_),
    .Y(_5277_)
);

INVX2 _15310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4816_),
    .Y(_4817_)
);

BUFX2 BUFX2_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .Y(_3529__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .Y(_3529__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .Y(_3529__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .Y(_3529__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529_),
    .Y(_3529__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf5)
);

BUFX2 BUFX2_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf4)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf3)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf2)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .Y(_2362__bF$buf1)
);

AOI21X1 _20387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10004_),
    .B(_10028_),
    .C(_10026_),
    .Y(_10382_)
);

NAND3X1 _16935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6583_),
    .B(_6588_),
    .C(_6587_),
    .Y(_6598_)
);

OAI21X1 _16515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5770_),
    .B(_5754_),
    .C(_5762_),
    .Y(_6137_)
);

FILL SFILL23960x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_374_),
    .Y(_812_)
);

NAND3X1 _12435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7272_),
    .B(_8095_),
    .C(_8106_),
    .Y(_8117_)
);

NAND2X1 _22953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1272_),
    .B(_1284_),
    .Y(_1285_)
);

NAND2X1 _12015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_4_bF$buf5),
    .Y(_3514_)
);

NAND3X1 _22533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_810_),
    .B(_815_),
    .C(_818_),
    .Y(_826_)
);

NAND2X1 _22113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_364_),
    .Y(_365_)
);

NAND2X1 _23738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_28_bF$buf5),
    .B(areg_31_bF$buf1),
    .Y(_2139_)
);

XOR2X1 _23318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1681_),
    .B(_1678_),
    .Y(_1682_)
);

AOI21X1 _17893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6804_),
    .B(_7646_),
    .C(_7647_),
    .Y(_7648_)
);

OAI21X1 _17473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7180_),
    .B(_7181_),
    .C(_6921_),
    .Y(_7188_)
);

NAND3X1 _17053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6721_),
    .B(_6727_),
    .C(_6677_),
    .Y(_6728_)
);

AOI21X1 _18678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8496_),
    .B(_8495_),
    .C(_8492_),
    .Y(_8508_)
);

NOR3X1 _18258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8025_),
    .B(_8032_),
    .C(_8035_),
    .Y(_8049_)
);

OAI21X1 _13393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_2715_),
    .C(_2579_),
    .Y(_2719_)
);

NAND2X1 _23491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1782_),
    .B(_1801_),
    .Y(_1871_)
);

AOI21X1 _23071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1273_),
    .B(_1283_),
    .C(_1411_),
    .Y(_1413_)
);

NAND2X1 _21804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11664_),
    .B(_11671_),
    .Y(_27_)
);

NAND3X1 _14598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4032_),
    .B(_4034_),
    .C(_4033_),
    .Y(_4038_)
);

OAI21X1 _14178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3345_),
    .B(_3353_),
    .C(_3355_),
    .Y(_3577_)
);

FILL SFILL64120x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10142_),
    .B(_10168_),
    .C(_10172_),
    .Y(_10173_)
);

OAI21X1 _16744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6381_),
    .B(_6382_),
    .C(_6129_),
    .Y(_6389_)
);

OAI21X1 _16324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5556_),
    .B(_5560_),
    .C(_5559_),
    .Y(_5929_)
);

NAND2X1 _17949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7288_),
    .B(_7295_),
    .Y(_7709_)
);

AOI21X1 _17529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6828_),
    .B(_6830_),
    .C(_6822_),
    .Y(_7248_)
);

OAI21X1 _17109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6784_),
    .B(_6785_),
    .C(_6423_),
    .Y(_6789_)
);

OAI21X1 _12664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10595_),
    .B(_10584_),
    .C(_10617_),
    .Y(_10628_)
);

NOR3X1 _12244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5815_),
    .B(_5826_),
    .C(_5837_),
    .Y(_6023_)
);

AOI21X1 _22762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .B(_1071_),
    .C(_1070_),
    .Y(_1077_)
);

NOR2X1 _22342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(_383_),
    .Y(_617_)
);

OAI21X1 _13869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3229_),
    .B(_3233_),
    .C(_2970_),
    .Y(_3239_)
);

OAI21X1 _13449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2557_),
    .B(_2558_),
    .C(_2566_),
    .Y(_2779_)
);

DFFPOSX1 _23967_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[21]),
    .CLK(clk_bF$buf10),
    .D(_0_[21])
);

OAI21X1 _13029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_2319_),
    .C(_1902_),
    .Y(_2324_)
);

AND2X2 _23547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1924_),
    .Y(_1932_)
);

AOI21X1 _23127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1472_),
    .C(_1465_),
    .Y(_1474_)
);

AOI21X1 _14810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4264_),
    .B(_4263_),
    .C(_4262_),
    .Y(_4269_)
);

NOR3X1 _17282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6961_),
    .B(_6971_),
    .C(_6972_),
    .Y(_6979_)
);

FILL SFILL34120x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8299_),
    .B(_8298_),
    .C(_8297_),
    .Y(_8300_)
);

AND2X2 _18067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7392_),
    .B(_7440_),
    .Y(_7839_)
);

FILL SFILL23960x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _11935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_2616_),
    .Y(_2639_)
);

XNOR2X1 _21613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11725_),
    .B(_11720_),
    .Y(_11726_)
);

OAI21X1 _22818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_777_),
    .B(_989_),
    .C(_991_),
    .Y(_1137_)
);

AOI21X1 _16973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6629_),
    .B(_6622_),
    .C(_6609_),
    .Y(_6640_)
);

OAI22X1 _16553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5795_),
    .B(_5842_),
    .C(_6178_),
    .D(_5840_),
    .Y(_6179_)
);

NAND2X1 _16133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5331_),
    .B(_5336_),
    .Y(_5719_)
);

NAND3X1 _17758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7495_),
    .B(_7498_),
    .C(_7499_),
    .Y(_7500_)
);

NOR3X1 _17338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7025_),
    .B(_7035_),
    .C(_7036_),
    .Y(_7040_)
);

XNOR2X1 _12893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1217_),
    .B(_1206_),
    .Y(_1228_)
);

AOI21X1 _12473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7931_),
    .B(_7997_),
    .C(_7294_),
    .Y(_8533_)
);

AOI21X1 _22991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .B(_1159_),
    .C(_1163_),
    .Y(_1326_)
);

INVX1 _12053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3854_),
    .Y(_3931_)
);

NOR2X1 _22571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_866_),
    .Y(_868_)
);

AOI22X1 _22151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_30_bF$buf1),
    .C(breg_16_bF$buf0),
    .D(areg_29_bF$buf1),
    .Y(_408_)
);

INVX1 _13678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2990_),
    .Y(_3030_)
);

NOR2X1 _13258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2568_),
    .B(_2567_),
    .Y(_2570_)
);

XOR2X1 _23776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2139_),
    .B(_2179_),
    .Y(_2180_)
);

NOR2X1 _23356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1694_),
    .B(_1723_),
    .Y(_1724_)
);

NAND2X1 _19904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9848_),
    .B(_9853_),
    .Y(_9854_)
);

OAI21X1 _17091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6767_),
    .B(_6768_),
    .C(_6766_),
    .Y(_6770_)
);

FILL SFILL33720x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg_20_bF$buf3),
    .Y(_5380_)
);

AOI21X1 _15404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4899_),
    .B(_4905_),
    .C(_4768_),
    .Y(_4921_)
);

AND2X2 _18296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg_27_bF$buf3),
    .Y(_8090_)
);

NOR3X1 _16609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6227_),
    .B(_6235_),
    .C(_6236_),
    .Y(_6240_)
);

NAND3X1 _21842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_63_),
    .B(_68_),
    .C(_26_),
    .Y(_69_)
);

OAI21X1 _21422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11512_),
    .B(_11517_),
    .C(_11440_),
    .Y(_11518_)
);

AND2X2 _21002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11052_),
    .B(_11056_),
    .Y(_11057_)
);

FILL SFILL13640x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11822_),
    .B(_11844_),
    .C(_11866_),
    .Y(_1838_)
);

NOR2X1 _12529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7689_),
    .B(_9137_),
    .Y(_9148_)
);

AOI21X1 _22627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9633_),
    .B(_926_),
    .C(_927_),
    .Y(_928_)
);

XNOR2X1 _12109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4314_),
    .B(_4259_),
    .Y(_4544_)
);

NAND3X1 _22207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_461_),
    .C(_463_),
    .Y(_469_)
);

NAND2X1 _16782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_28_bF$buf4),
    .Y(_6430_)
);

AOI21X1 _16362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5539_),
    .B(_5583_),
    .C(_5970_),
    .Y(_5971_)
);

BUFX2 BUFX2_insert460 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[23]),
    .Y(breg_23_bF$buf2)
);

BUFX2 BUFX2_insert461 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[23]),
    .Y(breg_23_bF$buf1)
);

BUFX2 BUFX2_insert462 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[23]),
    .Y(breg_23_bF$buf0)
);

BUFX2 BUFX2_insert463 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf4)
);

BUFX2 BUFX2_insert464 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf3)
);

NAND2X1 _17987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7295_),
    .B(_7299_),
    .Y(_7751_)
);

BUFX2 BUFX2_insert465 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf2)
);

NOR3X1 _17567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7276_),
    .B(_7277_),
    .C(_7279_),
    .Y(_7290_)
);

OAI21X1 _17147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5668__bF$buf0),
    .C(_6430_),
    .Y(_6830_)
);

BUFX2 BUFX2_insert466 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf1)
);

BUFX2 BUFX2_insert467 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[10]),
    .Y(areg_10_bF$buf0)
);

BUFX2 BUFX2_insert468 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[20]),
    .Y(breg_20_bF$buf4)
);

FILL SFILL23640x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert469 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[20]),
    .Y(breg_20_bF$buf3)
);

NOR2X1 _12282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4423_),
    .B(_5146_),
    .Y(_6439_)
);

OAI21X1 _22380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_420_),
    .B(_417_),
    .C(_412_),
    .Y(_658_)
);

FILL SFILL8680x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .Y(_2821_)
);

OAI21X1 _13067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2334_),
    .B(_1456_),
    .C(_2327_),
    .Y(_2361_)
);

INVX1 _23585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .Y(_1973_)
);

INVX2 _23165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .Y(_1516_)
);

FILL SFILL69000x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9387_),
    .B(_9643_),
    .C(_9595_),
    .Y(_9644_)
);

FILL SFILL8600x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _15633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4831_),
    .B(_4849_),
    .C(_5170_),
    .D(_4872_),
    .Y(_5171_)
);

OAI21X1 _15213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4403_),
    .B(_4392_),
    .C(_4396_),
    .Y(_4711_)
);

FILL SFILL74200x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6490_),
    .B(_6486_),
    .C(_6438_),
    .Y(_6491_)
);

AOI21X1 _16418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6016_),
    .B(_6020_),
    .C(_5665_),
    .Y(_6031_)
);

NAND2X1 _11973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_1_bF$buf3),
    .Y(_3055_)
);

AOI22X1 _21651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_30_bF$buf1),
    .C(breg_13_bF$buf2),
    .D(areg_29_bF$buf2),
    .Y(_11768_)
);

XNOR2X1 _21231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11003_),
    .B(_11307_),
    .Y(_0_[41])
);

FILL SFILL64280x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11297_),
    .B(_10002_),
    .C(_11395_),
    .Y(_11657_)
);

NAND3X1 _12338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7043_),
    .B(_6012_),
    .C(_7020_),
    .Y(_7054_)
);

NAND3X1 _22856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1059_),
    .B(_1178_),
    .C(_1174_),
    .Y(_1179_)
);

AOI22X1 _22436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11869_),
    .B(_11871_),
    .C(_11312_),
    .D(_11874_),
    .Y(_719_)
);

INVX2 _22016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .Y(_259_)
);

FILL SFILL64200x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5858_),
    .B(_5866_),
    .Y(_6221_)
);

INVX2 _16171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5754_),
    .Y(_5761_)
);

NOR2X1 _14904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4076_),
    .B(_4371_),
    .Y(_4372_)
);

AOI21X1 _17796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7110_),
    .B(_7114_),
    .C(_7117_),
    .Y(_7542_)
);

AOI21X1 _17376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6682_),
    .B(_6687_),
    .C(_6689_),
    .Y(_7082_)
);

NOR2X1 _12091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2814_),
    .B(_4336_),
    .Y(_4346_)
);

OAI21X1 _20922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10956_),
    .B(_10952_),
    .C(_10960_),
    .Y(_10970_)
);

OAI21X1 _20502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf3),
    .B(_5921__bF$buf2),
    .C(_10502_),
    .Y(_10509_)
);

OAI21X1 _13296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2443_),
    .C(_2434_),
    .Y(_2611_)
);

NAND3X1 _23394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1753_),
    .C(_1757_),
    .Y(_1766_)
);

OAI21X1 _19942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9892_),
    .B(_9893_),
    .C(_9894_),
    .Y(_9895_)
);

NAND3X1 _19522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9429_),
    .B(_9434_),
    .C(_9431_),
    .Y(_9435_)
);

NAND3X1 _19102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8935_),
    .B(_8973_),
    .C(_8967_),
    .Y(_8974_)
);

NOR3X1 _21707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11804_),
    .B(_11820_),
    .C(_11808_),
    .Y(_11829_)
);

OAI22X1 _15862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4771_),
    .B(_5419_),
    .C(_5421_),
    .D(_5105_),
    .Y(_5422_)
);

XNOR2X1 _15442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4648_),
    .B(_4961_),
    .Y(_0_[24])
);

NOR2X1 _15022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf1),
    .B(_2465__bF$buf2),
    .Y(_4502_)
);

INVX1 _20099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10044_),
    .Y(_10066_)
);

AOI21X1 _16647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6276_),
    .B(_6277_),
    .C(_6274_),
    .Y(_6282_)
);

NAND3X1 _16227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5820_),
    .B(_5821_),
    .C(_5819_),
    .Y(_5822_)
);

AND2X2 _21880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_26_bF$buf2),
    .Y(_110_)
);

AOI21X1 _21460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11273_),
    .B(_11269_),
    .C(_11281_),
    .Y(_11559_)
);

AND2X2 _21040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10766_),
    .B(_10758_),
    .Y(_11098_)
);

FILL SFILL13720x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .Y(_2249_)
);

AOI21X1 _12567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9510_),
    .B(_9499_),
    .C(_9488_),
    .Y(_9565_)
);

NOR2X1 _12147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4928_),
    .B(_4950_),
    .Y(_0_[7])
);

XNOR2X1 _22665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_957_),
    .Y(_970_)
);

NAND2X1 _22245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf3),
    .B(breg_28_bF$buf3),
    .Y(_510_)
);

OAI21X1 _14713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3891_),
    .B(_3875_),
    .C(_3883_),
    .Y(_4163_)
);

AOI21X1 _17185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6513_),
    .B(_6871_),
    .C(_6870_),
    .Y(_6872_)
);

FILL SFILL74200x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .B(_5481_),
    .Y(_5483_)
);

AOI21X1 _20731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10753_),
    .B(_10752_),
    .C(_10751_),
    .Y(_10760_)
);

NOR3X1 _20311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9930_),
    .B(_9936_),
    .C(_9940_),
    .Y(_10300_)
);

NAND3X1 _19751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9646_),
    .B(_9684_),
    .C(_9683_),
    .Y(_9686_)
);

AOI21X1 _19331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9223_),
    .B(_9224_),
    .C(_9222_),
    .Y(_9226_)
);

NAND2X1 _21936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11785_),
    .B(_11794_),
    .Y(_172_)
);

NAND2X1 _21516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_27_bF$buf4),
    .Y(_11620_)
);

FILL SFILL28840x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5187_),
    .B(_5192_),
    .Y(_5213_)
);

OAI21X1 _15251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4484_),
    .B(_4491_),
    .C(_4493_),
    .Y(_4753_)
);

NAND2X1 _16876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_19_bF$buf1),
    .Y(_6533_)
);

AND2X2 _16456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5688_),
    .B(_5750_),
    .Y(_6071_)
);

NAND3X1 _16036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5606_),
    .B(_5612_),
    .C(_5461_),
    .Y(_5613_)
);

FILL SFILL58920x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf3),
    .B(_5420__bF$buf0),
    .Y(_166_)
);

INVX2 _12376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7393_),
    .Y(_7470_)
);

AOI21X1 _22894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1186_),
    .B(_1187_),
    .C(_1185_),
    .Y(_1221_)
);

AOI21X1 _22474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_756_),
    .B(_760_),
    .C(_737_),
    .Y(_761_)
);

NOR2X1 _22054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_31_),
    .B(_300_),
    .Y(_301_)
);

NAND3X1 _18602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8419_),
    .B(_8420_),
    .C(_8418_),
    .Y(_8426_)
);

OAI21X1 _23679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2074_),
    .C(_2071_),
    .Y(_2075_)
);

NAND2X1 _23259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_31_bF$buf4),
    .Y(_1618_)
);

OAI21X1 _19807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9745_),
    .B(_9744_),
    .C(_9746_),
    .Y(_9747_)
);

NAND3X1 _14942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4391_),
    .B(_4413_),
    .C(_4409_),
    .Y(_4414_)
);

XNOR2X1 _14522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .B(_3949_),
    .Y(_3955_)
);

NOR2X1 _14102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3222_),
    .B(_3218_),
    .Y(_3495_)
);

FILL SFILL48920x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5258_),
    .B(_5249_),
    .C(_5255_),
    .Y(_5274_)
);

OAI21X1 _15307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4573_),
    .B(_4813_),
    .C(_4563_),
    .Y(_4814_)
);

NAND2X1 _20960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10800_),
    .B(_10806_),
    .Y(_11010_)
);

AND2X2 _20540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10181_),
    .B(_10173_),
    .Y(_10550_)
);

OAI21X1 _20120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10087_),
    .B(_10088_),
    .C(_10084_),
    .Y(_10089_)
);

NAND3X1 _18199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7982_),
    .B(_7983_),
    .C(_7981_),
    .Y(_7984_)
);

FILL SFILL13720x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9934_),
    .B(_9935_),
    .C(_9933_),
    .Y(_9936_)
);

AND2X2 _19560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9085_),
    .B(_9080_),
    .Y(_9476_)
);

NAND2X1 _19140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_20_bF$buf0),
    .Y(_9015_)
);

NAND3X1 _21745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11862_),
    .B(_11863_),
    .C(_11596_),
    .Y(_11870_)
);

NAND3X1 _21325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11369_),
    .B(_11405_),
    .C(_11410_),
    .Y(_11411_)
);

NAND3X1 _15480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4670_),
    .B(_5001_),
    .C(_4999_),
    .Y(_5002_)
);

NAND3X1 _15060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4538_),
    .B(_4542_),
    .C(_4540_),
    .Y(_4543_)
);

NAND2X1 _16685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6317_),
    .B(_6312_),
    .Y(_6324_)
);

AOI21X1 _16265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5852_),
    .B(_5851_),
    .C(_5849_),
    .Y(_5864_)
);

NAND3X1 _12185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5113_),
    .B(_5233_),
    .C(_5168_),
    .Y(_5376_)
);

NAND3X1 _22283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .B(_551_),
    .C(_550_),
    .Y(_552_)
);

FILL SFILL28920x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8636_),
    .B(_8669_),
    .C(_8672_),
    .Y(_8677_)
);

AOI21X1 _18411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8208_),
    .B(_8215_),
    .C(_8195_),
    .Y(_8217_)
);

AOI21X1 _23488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .B(_1854_),
    .C(_1857_),
    .Y(_1867_)
);

NOR2X1 _23068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf0),
    .B(_7225__bF$buf0),
    .Y(_1409_)
);

OAI21X1 _19616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_8759_),
    .C(_9537_),
    .Y(_9538_)
);

OAI21X1 _14751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3916_),
    .B(_4203_),
    .C(_3924_),
    .Y(_4205_)
);

NAND3X1 _14331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3741_),
    .B(_3739_),
    .C(_3740_),
    .Y(_3746_)
);

OAI21X1 _15956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3958__bF$buf2),
    .C(_5517_),
    .Y(_5525_)
);

AOI21X1 _15536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4794_),
    .B(_5063_),
    .C(_5062_),
    .Y(_5064_)
);

NAND3X1 _15116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4604_),
    .B(_4603_),
    .C(_4602_),
    .Y(_4605_)
);

FILL SFILL18840x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_213_),
    .C(_11886_),
    .Y(_214_)
);

NAND2X1 _21554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf0),
    .B(breg_21_bF$buf1),
    .Y(_11661_)
);

AOI21X1 _21134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11200_),
    .B(_11201_),
    .C(_11193_),
    .Y(_11202_)
);

FILL SFILL38920x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1070_),
    .B(_1072_),
    .C(_1071_),
    .Y(_1073_)
);

OAI21X1 _22339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4069_),
    .B(_5921__bF$buf3),
    .C(_611_),
    .Y(_613_)
);

NOR3X1 _13602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2714_),
    .B(_2715_),
    .C(_2713_),
    .Y(_2948_)
);

NAND2X1 _23700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2060_),
    .B(_2097_),
    .Y(_2098_)
);

NAND3X1 _16494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6053_),
    .B(_6112_),
    .C(_6113_),
    .Y(_6114_)
);

INVX1 _16074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5284_),
    .Y(_5655_)
);

NAND3X1 _14807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(_4265_),
    .C(_4235_),
    .Y(_4266_)
);

AOI21X1 _17699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7141_),
    .B(_7148_),
    .C(_7064_),
    .Y(_7435_)
);

AND2X2 _17279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6561_),
    .B(_6974_),
    .Y(_6975_)
);

NOR2X1 _22092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_342_),
    .Y(_343_)
);

OAI21X1 _18640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8453_),
    .B(_8456_),
    .C(_8459_),
    .Y(_8466_)
);

AOI21X1 _18220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7483_),
    .B(_7572_),
    .C(_8006_),
    .Y(_8007_)
);

NOR2X1 _20825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10855_),
    .B(_10856_),
    .Y(_10863_)
);

INVX1 _20405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10395_),
    .Y(_10402_)
);

NAND3X1 _13199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2501_),
    .B(_2505_),
    .C(_2377_),
    .Y(_2506_)
);

AND2X2 _23297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1571_),
    .B(_1556_),
    .Y(_1659_)
);

OAI21X1 _19845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9787_),
    .B(_9788_),
    .C(_9786_),
    .Y(_9789_)
);

OAI21X1 _19425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9327_),
    .B(_9326_),
    .C(_9322_),
    .Y(_9328_)
);

AOI21X1 _19005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8866_),
    .B(_8867_),
    .C(_8474_),
    .Y(_8868_)
);

FILL SFILL59080x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf4),
    .B(areg_12_bF$buf2),
    .Y(_4455_)
);

AOI21X1 _14560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3994_),
    .B(_3995_),
    .C(_3993_),
    .Y(_3996_)
);

INVX2 _14140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3534_),
    .Y(_3535_)
);

FILL SFILL3640x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _15765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf5),
    .Y(_5315_)
);

INVX2 _15345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4855_),
    .Y(_4856_)
);

FILL SFILL3560x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf3),
    .B(_6050__bF$buf3),
    .C(_11900_),
    .Y(_4_)
);

NOR2X1 _21363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11451_),
    .B(_11452_),
    .Y(_11453_)
);

FILL SFILL28920x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7247_),
    .B(_7233_),
    .C(_7257_),
    .Y(_7668_)
);

NOR2X1 _22988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1315_),
    .Y(_1322_)
);

OAI21X1 _22568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_406_),
    .B(_410_),
    .C(_649_),
    .Y(_864_)
);

NAND2X1 _22148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf2),
    .B(areg_28_bF$buf0),
    .Y(_404_)
);

NAND3X1 _13831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3192_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3199_)
);

OAI21X1 _13411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2737_),
    .C(_2735_),
    .Y(_2739_)
);

FILL SFILL18920x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .Y(_4056_)
);

AOI21X1 _17088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6217_),
    .B(_6369_),
    .C(_6765_),
    .Y(_6766_)
);

FILL SFILL18760x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10649_),
    .B(_10653_),
    .C(_10339_),
    .Y(_10654_)
);

AOI21X1 _20214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10190_),
    .B(_10181_),
    .C(_10192_),
    .Y(_10193_)
);

FILL SFILL63880x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9579_),
    .B(_9578_),
    .Y(_9580_)
);

AOI21X1 _19234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8710_),
    .B(_8712_),
    .C(_8718_),
    .Y(_9119_)
);

NAND3X1 _21839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .C(_61_),
    .Y(_65_)
);

NAND3X1 _21419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11509_),
    .B(_11510_),
    .C(_11508_),
    .Y(_11514_)
);

NAND3X1 _15994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5555_),
    .B(_5566_),
    .C(_5562_),
    .Y(_5567_)
);

NAND2X1 _15574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_13_bF$buf3),
    .Y(_5106_)
);

AOI21X1 _15154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4052_),
    .B(_4644_),
    .C(_4645_),
    .Y(_4646_)
);

NAND2X1 _16779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6425_),
    .B(_5669_),
    .Y(_6426_)
);

NAND3X1 _16359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5964_),
    .B(_5966_),
    .C(_5965_),
    .Y(_5967_)
);

NAND3X1 _21592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11700_),
    .B(_11702_),
    .C(_11696_),
    .Y(_11703_)
);

OAI21X1 _21172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11243_),
    .B(_11241_),
    .C(_11235_),
    .Y(_11244_)
);

OAI21X1 _17720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf1),
    .B(_3961__bF$buf2),
    .C(_7447_),
    .Y(_7458_)
);

OR2X2 _17300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6951_),
    .B(_6956_),
    .Y(_6998_)
);

XNOR2X1 _12699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10781_),
    .B(_10715_),
    .Y(_11011_)
);

AND2X2 _12279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6187_),
    .B(_6385_),
    .Y(_6407_)
);

OAI21X1 _22797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf2),
    .B(_5668__bF$buf1),
    .C(_959_),
    .Y(_1114_)
);

NAND3X1 _22377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_641_),
    .B(_654_),
    .C(_651_),
    .Y(_655_)
);

INVX2 _18925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8771_),
    .Y(_8780_)
);

NAND3X1 _18505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8301_),
    .B(_8309_),
    .C(_8288_),
    .Y(_8320_)
);

FILL SFILL59080x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2566_),
    .B(_2778_),
    .Y(_2988_)
);

NAND3X1 _13220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2529_)
);

FILL SFILL3640x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4307_),
    .B(_4306_),
    .C(_4305_),
    .Y(_4308_)
);

NAND3X1 _14425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3838_),
    .B(_3847_),
    .C(_3806_),
    .Y(_3848_)
);

INVX2 _14005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3387_),
    .Y(_3388_)
);

AND2X2 _20863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10535_),
    .B(_10527_),
    .Y(_10905_)
);

NAND2X1 _20443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10390_),
    .B(_10387_),
    .Y(_10444_)
);

NOR3X1 _20023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9618_),
    .B(_9622_),
    .C(_9625_),
    .Y(_9983_)
);

OAI21X1 _19883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9780_),
    .B(_9781_),
    .C(_9765_),
    .Y(_9831_)
);

NAND3X1 _19463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9369_),
    .B(_9360_),
    .C(_9317_),
    .Y(_9370_)
);

NOR2X1 _19043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8901_),
    .B(_8902_),
    .Y(_8909_)
);

FILL SFILL33880x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18600x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_11764_)
);

NAND3X1 _21228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11007_),
    .B(_11295_),
    .C(_11290_),
    .Y(_11305_)
);

NAND2X1 _12911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_1042_),
    .Y(_1423_)
);

OAI21X1 _15383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4896_),
    .B(_4897_),
    .C(_4894_),
    .Y(_4898_)
);

FILL SFILL18920x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6216_),
    .B(_6212_),
    .Y(_6217_)
);

AND2X2 _16168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_19_bF$buf2),
    .Y(_5757_)
);

FILL SFILL39000x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4292_),
    .B(_4303_),
    .Y(_4314_)
);

NOR2X1 _22186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_445_),
    .Y(_446_)
);

AOI21X1 _18734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8552_),
    .B(_8557_),
    .C(_8559_),
    .Y(_8570_)
);

NAND3X1 _18314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8083_),
    .B(_8108_),
    .C(_8109_),
    .Y(_8110_)
);

NAND3X1 _20919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10698_),
    .B(_10808_),
    .C(_10809_),
    .Y(_10966_)
);

FILL SFILL8760x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9887_),
    .B(_9888_),
    .C(_9886_),
    .Y(_9892_)
);

NAND2X1 _19519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9426_),
    .B(_9430_),
    .Y(_9431_)
);

OAI21X1 _14654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3836_),
    .B(_3834_),
    .C(_3825_),
    .Y(_4098_)
);

OAI21X1 _14234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3433_),
    .B(_3431_),
    .C(_3424_),
    .Y(_3639_)
);

FILL SFILL53960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5408_),
    .B(_5416_),
    .C(_5417_),
    .Y(_5418_)
);

NAND3X1 _15439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4951_),
    .B(_4944_),
    .C(_4947_),
    .Y(_4959_)
);

NAND2X1 _15019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_16_bF$buf2),
    .Y(_4498_)
);

INVX2 _20672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10694_),
    .Y(_10695_)
);

AOI21X1 _20252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10231_),
    .B(_10234_),
    .C(_10216_),
    .Y(_10235_)
);

OAI22X1 _16800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf0),
    .B(_5315__bF$buf3),
    .C(_2562__bF$buf1),
    .D(_5318_),
    .Y(_6449_)
);

AOI21X1 _19692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9621_),
    .B(_9619_),
    .C(_9269_),
    .Y(_9622_)
);

AOI21X1 _19272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9152_),
    .B(_9154_),
    .C(_9144_),
    .Y(_9161_)
);

AND2X2 _21877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11729_),
    .B(_105_),
    .Y(_107_)
);

NAND3X1 _21457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11258_),
    .B(_11547_),
    .C(_11548_),
    .Y(_11556_)
);

FILL SFILL3720x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10846_),
    .B(_10844_),
    .C(_11094_),
    .Y(_11095_)
);

FILL SFILL43960x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11231_),
    .B(_11187_),
    .C(_10419_),
    .Y(_11242_)
);

OAI21X1 _12300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6626_),
    .B(_6615_),
    .C(_6450_),
    .Y(_6637_)
);

NAND2X1 _15192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_19_bF$buf2),
    .Y(_4688_)
);

FILL SFILL43880x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3086_),
    .B(_3087_),
    .C(_3085_),
    .Y(_3301_)
);

OAI21X1 _13505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2685_),
    .B(_2651_),
    .C(_2696_),
    .Y(_2841_)
);

AOI21X1 _23603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1987_),
    .B(_1545_),
    .C(_1992_),
    .Y(_1993_)
);

NAND3X1 _16397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5988_),
    .B(_5995_),
    .C(_5998_),
    .Y(_6008_)
);

NOR2X1 _18963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8741_),
    .B(_8792_),
    .Y(_8822_)
);

NAND2X1 _18543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_28_bF$buf5),
    .Y(_8362_)
);

AOI21X1 _18123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7445_),
    .B(_7450_),
    .C(_7453_),
    .Y(_7901_)
);

FILL SFILL33880x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18600x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10406_),
    .B(_10466_),
    .Y(_10756_)
);

NAND3X1 _20308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10282_),
    .B(_10275_),
    .C(_10284_),
    .Y(_10296_)
);

OAI21X1 _19748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9681_),
    .B(_9677_),
    .C(_9647_),
    .Y(_9682_)
);

NOR2X1 _19328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9220_),
    .B(_9221_),
    .Y(_9222_)
);

NAND2X1 _14883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4060_),
    .B(_4062_),
    .Y(_4349_)
);

AND2X2 _14463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3879_),
    .B(_3877_),
    .Y(_3890_)
);

NAND3X1 _14043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3424_),
    .B(_3429_),
    .C(_3385_),
    .Y(_3430_)
);

FILL SFILL39080x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5200_),
    .B(_5198_),
    .C(_5196_),
    .Y(_5209_)
);

OAI21X1 _15248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4744_),
    .B(_4745_),
    .C(_4710_),
    .Y(_4749_)
);

NOR2X1 _20481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10119_),
    .B(_10484_),
    .Y(_10486_)
);

AOI21X1 _20061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10012_),
    .B(_10011_),
    .C(_10008_),
    .Y(_10025_)
);

FILL SFILL63960x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _19081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8192_),
    .B(_8948_),
    .C(_8949_),
    .D(_8603_),
    .Y(_8951_)
);

NOR3X1 _21686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11802_),
    .B(_11537_),
    .C(_11801_),
    .Y(_11806_)
);

FILL SFILL23800x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11340_),
    .B(_11344_),
    .C(_11333_),
    .Y(_11345_)
);

NAND2X1 _17814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7560_),
    .B(_7561_),
    .Y(_7562_)
);

FILL SFILL29080x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3087_),
    .B(_3078_),
    .C(_3082_),
    .Y(_3092_)
);

OAI21X1 _13314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_7711__bF$buf3),
    .C(_2427_),
    .Y(_2632_)
);

OAI21X1 _23832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .B(_2235_),
    .C(_2239_),
    .Y(_2240_)
);

NAND2X1 _23412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1784_),
    .B(_1682_),
    .Y(_1785_)
);

FILL SFILL29000x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4392_),
    .B(_4402_),
    .C(_4403_),
    .Y(_4410_)
);

INVX1 _14519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3950_),
    .Y(_3951_)
);

FILL SFILL74040x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_18_bF$buf1),
    .Y(_8612_)
);

AOI21X1 _18352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8146_),
    .B(_8147_),
    .C(_8145_),
    .Y(_8152_)
);

INVX2 _20957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11006_),
    .Y(_11007_)
);

AOI21X1 _20537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10251_),
    .B(_10253_),
    .C(_10546_),
    .Y(_10547_)
);

OAI21X1 _20117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10073_),
    .B(_10074_),
    .C(_10071_),
    .Y(_10086_)
);

FILL SFILL43960x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9932_),
    .B(_9931_),
    .Y(_9933_)
);

OAI21X1 _19557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9138_),
    .B(_9136_),
    .C(_9134_),
    .Y(_9473_)
);

NOR2X1 _19137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9010_),
    .B(_9011_),
    .Y(_9012_)
);

OAI21X1 _14692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3908_),
    .B(_3910_),
    .C(_3906_),
    .Y(_4140_)
);

NOR2X1 _14272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3407_),
    .B(_3680_),
    .Y(_3681_)
);

FILL SFILL43800x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5459_),
    .B(_5458_),
    .C(_5457_),
    .Y(_5460_)
);

NAND2X1 _15477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4998_),
    .B(_4997_),
    .Y(_4999_)
);

NAND2X1 _15057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4245_),
    .B(_4539_),
    .Y(_4540_)
);

NAND3X1 _20290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10110_),
    .B(_10203_),
    .C(_10202_),
    .Y(_10276_)
);

OAI21X1 _21495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11357_),
    .B(_11328_),
    .C(_11366_),
    .Y(_11597_)
);

OAI21X1 _21075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10818_),
    .B(_11135_),
    .C(_11136_),
    .Y(_11137_)
);

OAI21X1 _17623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6939_),
    .B(_6934_),
    .C(_6942_),
    .Y(_7352_)
);

OAI21X1 _17203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6884_),
    .B(_6883_),
    .C(_6881_),
    .Y(_6892_)
);

NAND3X1 _18828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8668_),
    .B(_8669_),
    .C(_8672_),
    .Y(_8673_)
);

NOR2X1 _18408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8200_),
    .B(_8198_),
    .Y(_8213_)
);

NAND3X1 _13963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3321_),
    .B(_3330_),
    .C(_3334_),
    .Y(_3342_)
);

OR2X2 _13543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2881_),
    .B(_2882_),
    .Y(_2883_)
);

OAI21X1 _13123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2131_),
    .C(_2315_),
    .Y(_2423_)
);

NAND2X1 _23641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2033_),
    .B(_2030_),
    .Y(_2035_)
);

NAND2X1 _23221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .B(_1575_),
    .Y(_1576_)
);

AOI21X1 _14748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3988_),
    .B(_3987_),
    .C(_3948_),
    .Y(_4201_)
);

AOI21X1 _14328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3741_),
    .B(_3740_),
    .C(_3739_),
    .Y(_3742_)
);

DFFPOSX1 _24006_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[60]),
    .CLK(clk_bF$buf9),
    .D(_0_[60])
);

FILL SFILL54280x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8323_),
    .B(_8325_),
    .C(_8318_),
    .Y(_8403_)
);

OAI21X1 _18161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7524_),
    .B(_7515_),
    .C(_7519_),
    .Y(_7943_)
);

FILL SFILL23800x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10795_),
    .B(_10796_),
    .C(_10797_),
    .Y(_10798_)
);

OAI21X1 _20346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9992_),
    .B(_10336_),
    .C(_10329_),
    .Y(_10337_)
);

FILL SFILL8840x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9342_),
    .B(_9336_),
    .Y(_9724_)
);

AOI21X1 _19366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9256_),
    .B(_8469_),
    .C(_9262_),
    .Y(_9263_)
);

AOI21X1 _14081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3470_),
    .B(_3469_),
    .C(_3462_),
    .Y(_3472_)
);

OAI21X1 _12814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_275_),
    .C(_232_),
    .Y(_373_)
);

NAND3X1 _22912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1101_),
    .B(_1236_),
    .C(_1237_),
    .Y(_1241_)
);

AOI21X1 _15286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4781_),
    .B(_4780_),
    .C(_4777_),
    .Y(_4791_)
);

FILL SFILL74440x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7597_),
    .B(_7341_),
    .C(_7603_),
    .Y(_7604_)
);

OAI21X1 _17432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7088_),
    .B(_7089_),
    .C(_7066_),
    .Y(_7144_)
);

NAND2X1 _17012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_25_bF$buf0),
    .Y(_6683_)
);

FILL SFILL49000x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3960x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_336_),
    .C(_337_),
    .Y(_339_)
);

XNOR2X1 _18637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8069_),
    .B(_8463_),
    .Y(_0_[33])
);

AOI21X1 _18217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8002_),
    .B(_8003_),
    .C(_8001_),
    .Y(_8004_)
);

OAI21X1 _13772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_2465__bF$buf2),
    .C(_3111_),
    .Y(_3133_)
);

INVX1 _23870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2261_),
    .Y(_2279_)
);

OAI21X1 _13352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2673_),
    .B(_2667_),
    .C(_2663_),
    .Y(_2674_)
);

NAND2X1 _23450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1820_),
    .B(_1822_),
    .Y(_1826_)
);

OAI21X1 _23030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1366_),
    .C(_1367_),
    .Y(_1368_)
);

XOR2X1 _14977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4450_),
    .B(_4451_),
    .Y(_4452_)
);

NAND2X1 _14557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3991_),
    .B(_3992_),
    .Y(_3993_)
);

XNOR2X1 _14137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3531_),
    .B(_3527_),
    .Y(_3532_)
);

XOR2X1 _18390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8191_),
    .B(_8192_),
    .Y(_8193_)
);

AOI21X1 _20995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11042_),
    .B(_11045_),
    .C(_11019_),
    .Y(_11049_)
);

OAI21X1 _20575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10587_),
    .B(_10588_),
    .C(_10262_),
    .Y(_10589_)
);

OAI22X1 _20155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf0),
    .B(_3958__bF$buf3),
    .C(_3402__bF$buf1),
    .D(_3253__bF$buf2),
    .Y(_10128_)
);

OAI21X1 _16703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6281_),
    .B(_6284_),
    .C(_6287_),
    .Y(_6344_)
);

NAND3X1 _19595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9513_),
    .B(_9514_),
    .C(_9512_),
    .Y(_9515_)
);

FILL SFILL54040x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_4551__bF$buf0),
    .C(_8657_),
    .Y(_9054_)
);

NAND2X1 _17908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7314_),
    .B(_7321_),
    .Y(_7664_)
);

FILL SFILL59160x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10145_),
    .B(_10167_),
    .C(_10079_),
    .Y(_10178_)
);

FILL SFILL33880x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5497_),
    .Y(_5574_)
);

NAND3X1 _22721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1028_),
    .B(_1029_),
    .C(_1030_),
    .Y(_1032_)
);

NAND3X1 _22301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_568_),
    .B(_569_),
    .C(_570_),
    .Y(_572_)
);

AOI21X1 _15095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4563_),
    .B(_4569_),
    .C(_4526_),
    .Y(_4582_)
);

OAI21X1 _13828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(_3194_),
    .C(_3049_),
    .Y(_3195_)
);

AOI21X1 _13408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2522_),
    .C(_2734_),
    .Y(_2735_)
);

BUFX2 _23926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[44]),
    .Y(y[44])
);

OAI21X1 _23506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668__bF$buf0),
    .B(_7520__bF$buf2),
    .C(_1795_),
    .Y(_1887_)
);

OAI22X1 _17661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6974_),
    .B(_7392_),
    .C(_7021_),
    .D(_7017_),
    .Y(_7394_)
);

NAND2X1 _17241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_20_bF$buf0),
    .Y(_6934_)
);

FILL SFILL48680x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8297_),
    .B(_8299_),
    .C(_8306_),
    .Y(_8715_)
);

AOI21X1 _18446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7844_),
    .B(_7846_),
    .C(_7851_),
    .Y(_8255_)
);

NAND2X1 _18026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_20_bF$buf0),
    .Y(_7794_)
);

NAND3X1 _13581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .B(_2923_),
    .C(_2840_),
    .Y(_2925_)
);

INVX8 _13161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf1),
    .Y(_2465_)
);

FILL SFILL69160x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf1),
    .B(areg_20_bF$buf3),
    .Y(_4243_)
);

NOR2X1 _14366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf0),
    .B(_3781__bF$buf3),
    .Y(_3782_)
);

DFFPOSX1 _24044_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[2]),
    .CLK(clk_bF$buf1),
    .D(b[2])
);

FILL SFILL28840x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10363_),
    .B(_10356_),
    .C(_10368_),
    .Y(_10379_)
);

OAI21X1 _16932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6594_),
    .B(_6589_),
    .C(_6512_),
    .Y(_6595_)
);

NAND2X1 _16512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_21_bF$buf0),
    .Y(_6134_)
);

NAND3X1 _21589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11685_),
    .B(_11692_),
    .C(_11689_),
    .Y(_11699_)
);

NOR2X1 _21169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11239_),
    .B(_11238_),
    .Y(_11240_)
);

FILL SFILL64120x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7454_),
    .B(_7453_),
    .C(_7444_),
    .Y(_7455_)
);

AOI21X1 _12852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_659_),
    .C(_473_),
    .Y(_779_)
);

NAND3X1 _12432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8073_),
    .B(_7283_),
    .C(_8008_),
    .Y(_8084_)
);

NAND2X1 _22950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1278_),
    .B(_1280_),
    .Y(_1281_)
);

NAND2X1 _12012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2858_),
    .Y(_3482_)
);

NAND3X1 _22530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_821_),
    .C(_770_),
    .Y(_822_)
);

FILL SFILL28680x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_353_),
    .C(_358_),
    .Y(_362_)
);

FILL SFILL54120x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2984_),
    .Y(_2985_)
);

NAND3X1 _13217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .B(_2524_),
    .C(_2525_),
    .Y(_2526_)
);

OAI21X1 _23735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2013_),
    .B(_2072_),
    .C(_2078_),
    .Y(_2136_)
);

NAND2X1 _23315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_26_bF$buf1),
    .B(breg_28_bF$buf5),
    .Y(_1679_)
);

FILL FILL74040x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7213_),
    .B(_6805_),
    .C(_7643_),
    .Y(_7644_)
);

NAND3X1 _17470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6915_),
    .B(_6908_),
    .C(_6913_),
    .Y(_7184_)
);

AOI21X1 _17050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6719_),
    .B(_6718_),
    .C(_6717_),
    .Y(_6724_)
);

FILL SFILL38680x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54040x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf0),
    .B(_6050__bF$buf0),
    .C(_8494_),
    .Y(_8505_)
);

NOR3X1 _18255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7614_),
    .B(_7615_),
    .C(_7613_),
    .Y(_8046_)
);

AOI21X1 _13390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .B(_2702_),
    .C(_2625_),
    .Y(_2715_)
);

AND2X2 _21801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_19_),
    .B(_22_),
    .Y(_24_)
);

AOI21X1 _14595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4034_),
    .B(_4033_),
    .C(_4032_),
    .Y(_4035_)
);

OAI21X1 _14175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3570_),
    .C(_3538_),
    .Y(_3574_)
);

NOR2X1 _12908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11538_),
    .B(_1336_),
    .Y(_1391_)
);

NOR3X1 _20193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10162_),
    .B(_10165_),
    .C(_10161_),
    .Y(_10170_)
);

NAND3X1 _16741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6123_),
    .B(_6124_),
    .C(_6125_),
    .Y(_6386_)
);

AND2X2 _16321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5918_),
    .B(_5919_),
    .Y(_5926_)
);

AOI21X1 _21398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11481_),
    .B(_11479_),
    .C(_11477_),
    .Y(_11491_)
);

AND2X2 _17946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7702_),
    .B(_7705_),
    .Y(_7706_)
);

NOR2X1 _17526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7237_),
    .B(_7238_),
    .Y(_7245_)
);

OAI21X1 _17106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6784_),
    .B(_6785_),
    .C(_6781_),
    .Y(_6786_)
);

AND2X2 _12661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10529_),
    .B(_10507_),
    .Y(_10595_)
);

OAI21X1 _12241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5837_),
    .B(_5826_),
    .C(_4981_),
    .Y(_5990_)
);

FILL SFILL69160x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3236_),
    .B(_3235_),
    .C(_2970_),
    .Y(_3237_)
);

DFFPOSX1 _23964_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[18]),
    .CLK(clk_bF$buf10),
    .D(_0_[18])
);

AOI21X1 _13446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2772_),
    .B(_2767_),
    .C(_2774_),
    .Y(_2776_)
);

OAI21X1 _13026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_2319_),
    .C(_2318_),
    .Y(_2321_)
);

NOR2X1 _23544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1829_),
    .B(_1924_),
    .Y(_1929_)
);

AOI21X1 _23124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1298_),
    .B(_1318_),
    .C(_1321_),
    .Y(_1471_)
);

INVX2 _18484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8290_),
    .Y(_8297_)
);

AOI21X1 _18064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7828_),
    .B(_7829_),
    .C(_7820_),
    .Y(_7836_)
);

FILL FILL74120x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _20669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10690_),
    .Y(_10691_)
);

AOI21X1 _20249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9864_),
    .B(_9869_),
    .C(_9873_),
    .Y(_10230_)
);

XNOR2X1 _11932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2605_),
    .B(_2530_),
    .Y(_2616_)
);

NOR2X1 _21610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11442_),
    .B(_11721_),
    .Y(_11722_)
);

AOI21X1 _19689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9610_),
    .B(_9617_),
    .C(_9270_),
    .Y(_9618_)
);

NOR2X1 _19269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8369_),
    .B(_9156_),
    .Y(_9157_)
);

FILL SFILL54120x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11154_),
    .B(_11165_),
    .C(_11143_),
    .Y(_11209_)
);

NAND3X1 _22815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_991_),
    .C(_993_),
    .Y(_1134_)
);

FILL SFILL33960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4375_),
    .B(_4377_),
    .C(_4372_),
    .Y(_4684_)
);

FILL FILL74040x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18760x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6281_),
    .B(_6287_),
    .C(_6289_),
    .Y(_6636_)
);

NAND3X1 _16550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6166_),
    .B(_6173_),
    .C(_6174_),
    .Y(_6175_)
);

OAI21X1 _16130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5708_),
    .B(_5709_),
    .C(_5706_),
    .Y(_5715_)
);

FILL SFILL18680x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_6300__bF$buf1),
    .C(_7486_),
    .Y(_7497_)
);

OAI21X1 _17335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7036_),
    .B(_7035_),
    .C(_7025_),
    .Y(_7037_)
);

OAI21X1 _12890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1173_),
    .B(_1184_),
    .C(_1162_),
    .Y(_1195_)
);

OAI21X1 _12470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8489_),
    .B(_7185_),
    .C(_8128_),
    .Y(_8500_)
);

INVX1 _12050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3887_),
    .Y(_3898_)
);

OAI21X1 _13675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3026_),
    .B(_3024_),
    .C(_2777_),
    .Y(_3027_)
);

INVX1 _13255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2566_),
    .Y(_2567_)
);

NOR2X1 _23773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9153_),
    .B(_6815__bF$buf3),
    .Y(_2177_)
);

XNOR2X1 _23353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1720_),
    .B(_1694_),
    .Y(_1721_)
);

AOI21X1 _19901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9844_),
    .B(_9843_),
    .C(_9846_),
    .Y(_9851_)
);

FILL SFILL69320x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5374_),
    .B(_5375_),
    .Y(_5377_)
);

OAI21X1 _15401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4758_),
    .B(_4754_),
    .C(_4761_),
    .Y(_4918_)
);

NAND2X1 _18293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_29_bF$buf3),
    .Y(_8087_)
);

OAI21X1 _20898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10941_),
    .B(_10942_),
    .C(_10940_),
    .Y(_10943_)
);

AOI21X1 _20478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10126_),
    .B(_10128_),
    .C(_10120_),
    .Y(_10482_)
);

OAI21X1 _20058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf3),
    .B(_6050__bF$buf1),
    .C(_10010_),
    .Y(_10021_)
);

OAI21X1 _16606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6236_),
    .B(_6235_),
    .C(_6227_),
    .Y(_6237_)
);

FILL SFILL69240x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf5),
    .B(breg_19_bF$buf3),
    .Y(_9408_)
);

NAND3X1 _19078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8944_),
    .B(_8946_),
    .C(_8945_),
    .Y(_8947_)
);

FILL SFILL38760x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_308_),
    .C(_1794_),
    .Y(_1805_)
);

OAI22X1 _12526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf0),
    .B(_9104__bF$buf1),
    .C(_3220_),
    .D(_7711__bF$buf1),
    .Y(_9115_)
);

NOR2X1 _22624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9974_),
    .B(_9971_),
    .Y(_925_)
);

NOR2X1 _12106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_4401_),
    .Y(_4511_)
);

NAND2X1 _22204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_212_),
    .Y(_466_)
);

FILL SFILL3800x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _23829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1993_),
    .B(_1986_),
    .C(_2209_),
    .Y(_2236_)
);

OAI21X1 _23409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1692_),
    .C(_1780_),
    .Y(_1781_)
);

FILL SFILL59240x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert430 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2586__bF$buf3)
);

BUFX2 BUFX2_insert431 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2586__bF$buf2)
);

BUFX2 BUFX2_insert432 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2586__bF$buf1)
);

BUFX2 BUFX2_insert433 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2586__bF$buf0)
);

AOI21X1 _17984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7730_),
    .B(_7735_),
    .C(_7737_),
    .Y(_7748_)
);

BUFX2 BUFX2_insert434 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .Y(_4541__bF$buf4)
);

OAI22X1 _17564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6514_),
    .B(_7286_),
    .C(_6929_),
    .D(_6925_),
    .Y(_7287_)
);

BUFX2 BUFX2_insert435 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .Y(_4541__bF$buf3)
);

NOR3X1 _17144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6820_),
    .B(_6822_),
    .C(_6826_),
    .Y(_6827_)
);

BUFX2 BUFX2_insert436 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .Y(_4541__bF$buf2)
);

BUFX2 BUFX2_insert437 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .Y(_4541__bF$buf1)
);

BUFX2 BUFX2_insert438 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541_),
    .Y(_4541__bF$buf0)
);

BUFX2 BUFX2_insert439 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[16]),
    .Y(areg_16_bF$buf5)
);

FILL SFILL59160x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8213_),
    .B(_8197_),
    .C(_8204_),
    .Y(_8608_)
);

NAND3X1 _18349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8145_),
    .B(_8146_),
    .C(_8147_),
    .Y(_8148_)
);

AOI21X1 _13484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2808_),
    .B(_2817_),
    .C(_2806_),
    .Y(_2818_)
);

NOR2X1 _13064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2337_),
    .B(_2357_),
    .Y(_2358_)
);

NOR3X1 _23582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1969_),
    .B(_1965_),
    .C(_2545_),
    .Y(_1970_)
);

NAND3X1 _23162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1503_),
    .C(_1494_),
    .Y(_1513_)
);

NAND2X1 _19710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9376_),
    .B(_9382_),
    .Y(_9640_)
);

FILL SFILL33960x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4131_),
    .B(_4132_),
    .C(_4098_),
    .Y(_4136_)
);

OAI21X1 _14269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3409_),
    .B(_3397_),
    .C(_3401_),
    .Y(_3677_)
);

FILL SFILL49160x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5161_),
    .B(_5162_),
    .C(_5153_),
    .Y(_5167_)
);

NAND3X1 _15210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4704_),
    .B(_4706_),
    .C(_4705_),
    .Y(_4707_)
);

NAND2X1 _20287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10270_),
    .B(_10267_),
    .Y(_10273_)
);

NAND3X1 _16835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6481_),
    .B(_6484_),
    .C(_6482_),
    .Y(_6488_)
);

OAI21X1 _16415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6026_),
    .B(_6027_),
    .C(_6022_),
    .Y(_6028_)
);

AND2X2 _11970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2968_),
    .B(_2705_),
    .Y(_3022_)
);

FILL SFILL39160x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11603_),
    .B(_11614_),
    .C(_11592_),
    .Y(_11625_)
);

OAI21X1 _12335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6977_),
    .B(_6988_),
    .C(_6034_),
    .Y(_7031_)
);

OAI21X1 _22853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1170_),
    .B(_1171_),
    .C(_1133_),
    .Y(_1176_)
);

INVX1 _22433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .Y(_716_)
);

INVX2 _22013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .Y(_256_)
);

FILL SFILL69320x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5676_),
    .B(_8773_),
    .Y(_2031_)
);

AOI21X1 _23218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1463_),
    .C(_1466_),
    .Y(_1573_)
);

AOI21X1 _14901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4082_),
    .B(_4085_),
    .C(_4077_),
    .Y(_4369_)
);

NAND2X1 _17793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7538_),
    .B(_7111_),
    .Y(_7539_)
);

NAND3X1 _17373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7073_),
    .B(_7077_),
    .C(_7078_),
    .Y(_7079_)
);

AOI21X1 _18998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8075_),
    .B(_8445_),
    .C(_8859_),
    .Y(_8860_)
);

NAND3X1 _18578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8395_),
    .B(_8398_),
    .C(_8394_),
    .Y(_8399_)
);

OAI21X1 _18158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf2),
    .B(_6300__bF$buf0),
    .C(_7935_),
    .Y(_7939_)
);

NAND2X1 _13293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .B(_2599_),
    .Y(_2608_)
);

OAI21X1 _23391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1761_),
    .B(_1758_),
    .C(_1657_),
    .Y(_1763_)
);

NAND3X1 _21704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11824_),
    .B(_11825_),
    .C(_11823_),
    .Y(_11826_)
);

NAND3X1 _14498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3926_),
    .B(_3927_),
    .C(_3925_),
    .Y(_3928_)
);

AOI21X1 _14078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3207_),
    .B(_3210_),
    .C(_3467_),
    .Y(_3468_)
);

FILL SFILL64120x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1229_),
    .B(_1225_),
    .C(_1103_),
    .Y(_1237_)
);

FILL FILL74200x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9785_),
    .B(_10062_),
    .C(_9760_),
    .Y(_10063_)
);

AOI21X1 _16644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5917_),
    .B(_5922_),
    .C(_5924_),
    .Y(_6279_)
);

OR2X2 _16224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5774_),
    .B(_5778_),
    .Y(_5819_)
);

AOI21X1 _17849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7595_),
    .B(_7594_),
    .C(_7593_),
    .Y(_7600_)
);

OAI21X1 _17429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7138_),
    .B(_7139_),
    .C(_7137_),
    .Y(_7140_)
);

OAI21X1 _17009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6678_),
    .B(_6331_),
    .C(_6322_),
    .Y(_6679_)
);

XNOR2X1 _12984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2163_),
    .Y(_2217_)
);

NAND3X1 _12564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9477_),
    .B(_9521_),
    .C(_8544_),
    .Y(_9532_)
);

AOI21X1 _12144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4917_),
    .B(_4906_),
    .C(_4008_),
    .Y(_4928_)
);

NAND3X1 _22662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_963_),
    .B(_960_),
    .C(_966_),
    .Y(_967_)
);

INVX2 _22242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .Y(_507_)
);

NOR2X1 _13769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf2),
    .B(_549__bF$buf4),
    .Y(_3129_)
);

NOR2X1 _23867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2275_),
    .B(_2276_),
    .Y(_2277_)
);

OAI21X1 _13349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_2669__bF$buf0),
    .C(_2665_),
    .Y(_2670_)
);

AND2X2 _23447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .B(_1820_),
    .Y(_1823_)
);

AOI21X1 _23027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1343_),
    .C(_1341_),
    .Y(_1365_)
);

NAND2X1 _14710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_12_bF$buf4),
    .Y(_4159_)
);

AOI21X1 _17182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6858_),
    .B(_6855_),
    .C(_6852_),
    .Y(_6869_)
);

FILL SFILL34040x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .B(_5479_),
    .C(_5477_),
    .Y(_5480_)
);

INVX2 _18387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8189_),
    .Y(_8190_)
);

NAND3X1 _21933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .B(_154_),
    .C(_126_),
    .Y(_169_)
);

NAND2X1 _21513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_28_bF$buf1),
    .Y(_11617_)
);

INVX1 _22718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .Y(_1028_)
);

FILL SFILL74280x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6525_),
    .B(_6529_),
    .C(_6518_),
    .Y(_6530_)
);

OAI21X1 _16453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_5315__bF$buf0),
    .C(_6062_),
    .Y(_6068_)
);

FILL SFILL13960x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5604_),
    .B(_5603_),
    .C(_5602_),
    .Y(_5610_)
);

OAI21X1 _17658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_2669__bF$buf1),
    .C(_7384_),
    .Y(_7390_)
);

NOR2X1 _17238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6928_),
    .B(_6929_),
    .Y(_6930_)
);

NAND2X1 _12793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_89_),
    .B(_122_),
    .Y(_133_)
);

OR2X2 _12373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6143_),
    .B(_7426_),
    .Y(_7437_)
);

INVX2 _22891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1216_),
    .Y(_1218_)
);

OAI21X1 _22471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_754_),
    .C(_740_),
    .Y(_758_)
);

OAI21X1 _22051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_33_),
    .C(_37_),
    .Y(_298_)
);

INVX1 _13998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3360_),
    .Y(_3380_)
);

AOI21X1 _13578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2917_),
    .B(_2916_),
    .C(_2915_),
    .Y(_2921_)
);

NAND2X1 _13158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_15_bF$buf3),
    .Y(_2461_)
);

NAND2X1 _23676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_28_bF$buf5),
    .B(areg_30_bF$buf0),
    .Y(_2072_)
);

NAND3X1 _23256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1603_),
    .B(_1605_),
    .C(_1607_),
    .Y(_1615_)
);

AOI21X1 _19804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9738_),
    .B(_9739_),
    .C(_9737_),
    .Y(_9744_)
);

FILL SFILL33720x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4929_),
    .B(_4930_),
    .C(_4925_),
    .Y(_5271_)
);

NAND3X1 _15304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4808_),
    .B(_4810_),
    .C(_4809_),
    .Y(_4811_)
);

AOI21X1 _18196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7527_),
    .B(_7545_),
    .C(_7980_),
    .Y(_7981_)
);

AOI21X1 _16929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6577_),
    .B(_6581_),
    .C(_6545_),
    .Y(_6591_)
);

NAND2X1 _16509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5810_),
    .B(_5818_),
    .Y(_6130_)
);

NAND2X1 _21742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11309_),
    .B(_11311_),
    .Y(_11867_)
);

NOR3X1 _21322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11401_),
    .B(_11402_),
    .C(_11403_),
    .Y(_11408_)
);

OAI21X1 _12849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_648_),
    .C(_494_),
    .Y(_746_)
);

AOI21X1 _12429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8040_),
    .B(_8041_),
    .C(_7964_),
    .Y(_8052_)
);

OAI21X1 _22947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf3),
    .B(_6427_),
    .C(_1277_),
    .Y(_1278_)
);

NAND2X1 _12009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3405_),
    .B(_3427_),
    .Y(_3449_)
);

AOI21X1 _22527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_813_),
    .C(_811_),
    .Y(_819_)
);

OAI21X1 _22107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_356_),
    .B(_357_),
    .C(_358_),
    .Y(_359_)
);

OAI21X1 _16682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6320_),
    .B(_6314_),
    .C(_6309_),
    .Y(_6321_)
);

OAI21X1 _16262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf1),
    .B(_2884__bF$buf1),
    .C(_5850_),
    .Y(_5861_)
);

AOI21X1 _17887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7634_),
    .B(_7636_),
    .C(_7202_),
    .Y(_7641_)
);

AOI21X1 _17467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7163_),
    .B(_7169_),
    .C(_7013_),
    .Y(_7181_)
);

NAND3X1 _17047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6679_),
    .B(_6720_),
    .C(_6716_),
    .Y(_6721_)
);

AOI21X1 _12182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5289_),
    .B(_5332_),
    .C(_5003_),
    .Y(_5343_)
);

INVX1 _22280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .Y(_548_)
);

FILL SFILL69400x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2499_),
    .B(_2498_),
    .C(_2496_),
    .Y(_2712_)
);

XOR2X1 _23485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1774_),
    .B(_1864_),
    .Y(_0_[54])
);

AOI21X1 _23065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .B(_1377_),
    .C(_1383_),
    .Y(_1406_)
);

AND2X2 _19613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_30_bF$buf3),
    .Y(_9535_)
);

FILL SFILL13640x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5516_),
    .B(_5521_),
    .C(_5520_),
    .Y(_5522_)
);

AOI21X1 _15533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5050_),
    .B(_5049_),
    .C(_5045_),
    .Y(_5061_)
);

NAND2X1 _15113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4600_),
    .B(_4601_),
    .Y(_4602_)
);

FILL SFILL74200x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6364_),
    .B(_6369_),
    .C(_6217_),
    .Y(_6382_)
);

OAI21X1 _16318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_5921__bF$buf1),
    .C(_5918_),
    .Y(_5922_)
);

AOI21X1 _21971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_204_),
    .C(_11829_),
    .Y(_211_)
);

OR2X2 _21551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11651_),
    .B(_11652_),
    .Y(_11658_)
);

AOI21X1 _21131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10852_),
    .B(_10875_),
    .C(_10878_),
    .Y(_11199_)
);

FILL SFILL64280x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8972_),
    .B(_9005_),
    .C(_10551_),
    .Y(_10562_)
);

INVX1 _12238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5947_),
    .Y(_5958_)
);

INVX1 _22756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .Y(_1070_)
);

NAND2X1 _22336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf4),
    .B(areg_24_bF$buf0),
    .Y(_610_)
);

FILL SFILL33800x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6054_),
    .B(_6109_),
    .C(_6102_),
    .Y(_6111_)
);

AOI21X1 _16071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5641_),
    .B(_5634_),
    .C(_5306_),
    .Y(_5652_)
);

OAI21X1 _14804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4256_),
    .B(_4255_),
    .C(_4242_),
    .Y(_4263_)
);

OAI21X1 _17696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7423_),
    .B(_7424_),
    .C(_7421_),
    .Y(_7432_)
);

NOR2X1 _17276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6963_),
    .B(_6964_),
    .Y(_6972_)
);

NAND3X1 _20822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10854_),
    .B(_10859_),
    .C(_10857_),
    .Y(_10860_)
);

NOR2X1 _20402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10396_),
    .B(_10398_),
    .Y(_10399_)
);

FILL SFILL58920x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2499_),
    .B(_2498_),
    .C(_2423_),
    .Y(_2503_)
);

OAI21X1 _23294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1655_),
    .C(_1654_),
    .Y(_1656_)
);

XNOR2X1 _19842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9763_),
    .B(_9785_),
    .Y(_9786_)
);

NAND2X1 _19422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_24_bF$buf3),
    .Y(_9325_)
);

AOI21X1 _19002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8864_),
    .B(_8858_),
    .C(_8475_),
    .Y(_8865_)
);

FILL SFILL23720x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf3),
    .B(areg_3_bF$buf4),
    .Y(_2573_)
);

NAND2X1 _21607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_23_bF$buf0),
    .Y(_11719_)
);

AND2X2 _15762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_25_bF$buf0),
    .Y(_5312_)
);

XNOR2X1 _15342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4852_),
    .B(_4848_),
    .Y(_4853_)
);

OAI21X1 _16967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6627_),
    .B(_6628_),
    .C(_6610_),
    .Y(_6633_)
);

NAND3X1 _16547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6167_),
    .B(_6171_),
    .C(_6170_),
    .Y(_6172_)
);

NAND3X1 _16127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5673_),
    .B(_5707_),
    .C(_5711_),
    .Y(_5712_)
);

OAI21X1 _21780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11907_),
    .B(_11906_),
    .C(_11896_),
    .Y(_11908_)
);

NOR2X1 _21360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11155_),
    .B(_11448_),
    .Y(_11449_)
);

FILL SFILL8600x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11450_),
    .B(_11461_),
    .C(_11472_),
    .Y(_1162_)
);

NAND3X1 _12467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6012_),
    .B(_8424_),
    .C(_8457_),
    .Y(_8467_)
);

NAND3X1 _22985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1298_),
    .B(_1318_),
    .C(_1316_),
    .Y(_1319_)
);

NOR3X1 _12047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3723_),
    .B(_3756_),
    .C(_3788_),
    .Y(_3865_)
);

NAND2X1 _22565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .B(_859_),
    .Y(_861_)
);

AOI21X1 _22145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .B(_152_),
    .C(_400_),
    .Y(_401_)
);

INVX1 _14613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4052_),
    .Y(_4053_)
);

NAND3X1 _17085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6761_),
    .B(_6762_),
    .C(_6760_),
    .Y(_6763_)
);

FILL SFILL74200x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_21_bF$buf2),
    .Y(_5373_)
);

NAND3X1 _20631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10344_),
    .B(_10644_),
    .C(_10647_),
    .Y(_10651_)
);

NAND3X1 _20211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10187_),
    .B(_10186_),
    .C(_10188_),
    .Y(_10190_)
);

AOI21X1 _19651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9571_),
    .B(_9575_),
    .C(_9481_),
    .Y(_9577_)
);

FILL SFILL64280x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _19231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_7217__bF$buf4),
    .D(_6300__bF$buf0),
    .Y(_9116_)
);

FILL SFILL3880x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_58_),
    .B(_59_),
    .C(_61_),
    .Y(_62_)
);

AOI21X1 _21416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11509_),
    .B(_11510_),
    .C(_11508_),
    .Y(_11511_)
);

FILL SFILL33800x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf1),
    .B(areg_26_bF$buf2),
    .Y(_5564_)
);

OAI21X1 _15571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4902_),
    .B(_4904_),
    .C(_4892_),
    .Y(_5103_)
);

NAND2X1 _15151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3513_),
    .B(_4641_),
    .Y(_4643_)
);

OAI21X1 _16776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6422_),
    .B(_6388_),
    .C(_6378_),
    .Y(_6423_)
);

NAND2X1 _16356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5962_),
    .B(_5963_),
    .Y(_5964_)
);

FILL SFILL18840x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10880_),
    .B(_10858_),
    .C(_10825_),
    .Y(_10979_)
);

INVX2 _12276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6363_),
    .Y(_6374_)
);

NOR2X1 _22794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf3),
    .B(_6815__bF$buf4),
    .Y(_1111_)
);

AOI21X1 _22374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_415_),
    .C(_419_),
    .Y(_652_)
);

XNOR2X1 _18922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8776_),
    .B(_8771_),
    .Y(_8777_)
);

AOI21X1 _18502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7930_),
    .B(_7948_),
    .C(_8316_),
    .Y(_8317_)
);

DFFPOSX1 _23999_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[53]),
    .CLK(clk_bF$buf6),
    .D(_0_[53])
);

OAI21X1 _23579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1962_),
    .B(_1965_),
    .C(_4646_),
    .Y(_1966_)
);

OAI21X1 _23159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1508_),
    .B(_1504_),
    .C(_1364_),
    .Y(_1509_)
);

OAI21X1 _19707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9307_),
    .B(_9280_),
    .C(_9315_),
    .Y(_9637_)
);

NAND2X1 _14842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4302_),
    .B(_4304_),
    .Y(_4305_)
);

AOI21X1 _14422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3844_),
    .B(_3842_),
    .C(_3834_),
    .Y(_3845_)
);

AND2X2 _14002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3384_),
    .B(_3379_),
    .Y(_3385_)
);

FILL SFILL48920x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4831_),
    .B(_4849_),
    .Y(_5164_)
);

XOR2X1 _15207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4682_),
    .B(_4678_),
    .Y(_4704_)
);

AOI21X1 _20860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10556_),
    .B(_10589_),
    .C(_10900_),
    .Y(_10901_)
);

AOI21X1 _20440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10428_),
    .B(_10424_),
    .C(_10393_),
    .Y(_10440_)
);

NAND3X1 _20020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9978_),
    .B(_9979_),
    .C(_9977_),
    .Y(_9980_)
);

AOI21X1 _18099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7869_),
    .B(_7868_),
    .C(_7870_),
    .Y(_7874_)
);

FILL SFILL44120x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9825_),
    .B(_9826_),
    .C(_9793_),
    .Y(_9827_)
);

AOI21X1 _19460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9365_),
    .B(_9364_),
    .C(_9355_),
    .Y(_9366_)
);

NAND3X1 _19040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8900_),
    .B(_8904_),
    .C(_8903_),
    .Y(_8905_)
);

NAND2X1 _11967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2968_),
    .Y(_2989_)
);

NAND2X1 _21645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_11761_)
);

NOR3X1 _21225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10982_),
    .B(_10978_),
    .C(_10984_),
    .Y(_11302_)
);

AOI21X1 _15380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4526_),
    .B(_4569_),
    .C(_4893_),
    .Y(_4894_)
);

FILL SFILL38920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6207_),
    .B(_6208_),
    .C(_6210_),
    .Y(_6214_)
);

NAND2X1 _16165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_20_bF$buf3),
    .Y(_5754_)
);

NAND2X1 _12085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf4),
    .B(breg_3_bF$buf0),
    .Y(_4281_)
);

OAI21X1 _22183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_442_),
    .C(_178_),
    .Y(_443_)
);

NAND3X1 _18731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8528_),
    .B(_8565_),
    .C(_8560_),
    .Y(_8567_)
);

OAI21X1 _18311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8105_),
    .B(_8099_),
    .C(_8085_),
    .Y(_8107_)
);

NAND3X1 _20916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10962_),
    .B(_10955_),
    .C(_10960_),
    .Y(_10963_)
);

AOI21X1 _23388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1755_),
    .B(_1756_),
    .C(_1754_),
    .Y(_1759_)
);

NAND3X1 _19936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9887_),
    .B(_9888_),
    .C(_9886_),
    .Y(_9889_)
);

NAND2X1 _19516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf1),
    .B(areg_19_bF$buf4),
    .Y(_9428_)
);

NAND3X1 _14651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4086_),
    .C(_4074_),
    .Y(_4095_)
);

NOR3X1 _14231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3619_),
    .B(_3626_),
    .C(_3625_),
    .Y(_3636_)
);

NAND3X1 _15856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5410_),
    .B(_5414_),
    .C(_5413_),
    .Y(_5415_)
);

OAI21X1 _15436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4955_),
    .B(_4954_),
    .C(_4951_),
    .Y(_4956_)
);

NAND2X1 _15016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4494_),
    .B(_4490_),
    .Y(_4495_)
);

NAND2X1 _21874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf3),
    .B(areg_24_bF$buf4),
    .Y(_104_)
);

NAND3X1 _21454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11326_),
    .B(_11436_),
    .C(_11435_),
    .Y(_11553_)
);

AOI21X1 _21034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11085_),
    .B(_11086_),
    .C(_11084_),
    .Y(_11092_)
);

FILL SFILL38920x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf3),
    .B(_6427_),
    .Y(_963_)
);

INVX1 _22239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .Y(_503_)
);

NAND3X1 _13922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3291_),
    .B(_3297_),
    .C(_3294_),
    .Y(_3298_)
);

AOI21X1 _13502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2820_),
    .B(_2824_),
    .C(_2827_),
    .Y(_2838_)
);

NAND2X1 _23600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1943_),
    .B(_1865_),
    .Y(_1989_)
);

NAND3X1 _16394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .B(_5740_),
    .C(_5741_),
    .Y(_6005_)
);

FILL SFILL48920x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf0),
    .B(_2379_),
    .Y(_4156_)
);

NAND3X1 _17599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7322_),
    .B(_7324_),
    .C(_7323_),
    .Y(_7325_)
);

OAI22X1 _17179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6134_),
    .B(_6863_),
    .C(_6540_),
    .D(_6864_),
    .Y(_6865_)
);

OAI22X1 _18960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8814_),
    .B(_8815_),
    .C(_8817_),
    .D(_8816_),
    .Y(_8818_)
);

OAI21X1 _18540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8356_),
    .B(_8357_),
    .C(_8355_),
    .Y(_8358_)
);

OAI21X1 _18120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_4541__bF$buf1),
    .C(_7452_),
    .Y(_7897_)
);

OAI21X1 _20725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf3),
    .B(_5315__bF$buf4),
    .C(_10745_),
    .Y(_10753_)
);

NAND3X1 _20305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10105_),
    .B(_9999_),
    .C(_10106_),
    .Y(_10293_)
);

XNOR2X1 _13099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2395_),
    .B(_2392_),
    .Y(_2396_)
);

INVX2 _23197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .Y(_1550_)
);

AOI21X1 _19745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9673_),
    .B(_9675_),
    .C(_9649_),
    .Y(_9679_)
);

AOI21X1 _19325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9218_),
    .B(_9212_),
    .C(_9002_),
    .Y(_9219_)
);

FILL SFILL59080x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4335_),
    .B(_4344_),
    .Y(_4345_)
);

OAI21X1 _14460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .B(_3885_),
    .C(_3874_),
    .Y(_3886_)
);

AOI21X1 _14040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3421_),
    .B(_3422_),
    .C(_3420_),
    .Y(_3426_)
);

FILL SFILL38920x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34200x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5194_),
    .B(_5205_),
    .C(_5202_),
    .Y(_5206_)
);

OAI21X1 _15245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4744_),
    .B(_4745_),
    .C(_4740_),
    .Y(_4746_)
);

OAI21X1 _21683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11801_),
    .B(_11802_),
    .C(_11537_),
    .Y(_11803_)
);

NOR2X1 _21263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11030_),
    .B(_11341_),
    .Y(_11342_)
);

FILL SFILL28920x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7552_),
    .B(_7511_),
    .C(_7557_),
    .Y(_7559_)
);

XNOR2X1 _22888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_868_),
    .Y(_1214_)
);

NOR2X1 _22468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_743_),
    .Y(_754_)
);

AOI21X1 _22048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .C(_55_),
    .Y(_294_)
);

OAI21X1 _13731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3085_),
    .B(_3086_),
    .C(_3087_),
    .Y(_3089_)
);

OR2X2 _13311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2627_),
    .Y(_2629_)
);

AOI21X1 _14936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4156_),
    .B(_4406_),
    .C(_4405_),
    .Y(_4407_)
);

OAI21X1 _14516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3676_),
    .B(_3947_),
    .C(_3697_),
    .Y(_3948_)
);

AOI21X1 _20954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10985_),
    .B(_10986_),
    .C(_10692_),
    .Y(_11004_)
);

AOI21X1 _20534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10538_),
    .B(_10537_),
    .C(_10536_),
    .Y(_10544_)
);

NAND3X1 _20114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10077_),
    .B(_10042_),
    .C(_10082_),
    .Y(_10083_)
);

AOI21X1 _19974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9923_),
    .B(_9929_),
    .C(_9854_),
    .Y(_9930_)
);

OAI21X1 _19554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9468_),
    .B(_9463_),
    .C(_9469_),
    .Y(_9470_)
);

NAND2X1 _19134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_21_bF$buf4),
    .Y(_9009_)
);

NAND3X1 _21739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11862_),
    .B(_11863_),
    .C(_11861_),
    .Y(_11864_)
);

OAI21X1 _21319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11402_),
    .B(_11401_),
    .C(_11403_),
    .Y(_11404_)
);

AND2X2 _15894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5079_),
    .B(_5072_),
    .Y(_5457_)
);

NAND3X1 _15474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4993_),
    .B(_4995_),
    .C(_4994_),
    .Y(_4996_)
);

NAND2X1 _15054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf1),
    .B(areg_21_bF$buf1),
    .Y(_4537_)
);

NAND2X1 _16679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf1),
    .B(areg_27_bF$buf4),
    .Y(_6317_)
);

OAI21X1 _16259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5856_),
    .B(_5855_),
    .C(_5847_),
    .Y(_5857_)
);

OAI21X1 _21492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11315_),
    .B(_11593_),
    .C(_11591_),
    .Y(_11594_)
);

NAND2X1 _21072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .B(breg_23_bF$buf3),
    .Y(_11134_)
);

AND2X2 _17620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7286_),
    .B(_7346_),
    .Y(_7348_)
);

NAND3X1 _17200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6848_),
    .B(_6882_),
    .C(_6887_),
    .Y(_6888_)
);

NAND3X1 _12599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9839_),
    .B(_9817_),
    .C(_9762_),
    .Y(_9915_)
);

NOR3X1 _12179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5256_),
    .B(_5113_),
    .C(_5267_),
    .Y(_5310_)
);

INVX2 _22697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_981_),
    .Y(_1005_)
);

NOR2X1 _22277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf1),
    .B(_5676_),
    .Y(_545_)
);

FILL SFILL3560x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8656_),
    .B(_8652_),
    .C(_8655_),
    .Y(_8670_)
);

NAND3X1 _18405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8203_),
    .B(_8206_),
    .C(_8204_),
    .Y(_8210_)
);

FILL SFILL59080x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3338_),
    .B(_3335_),
    .C(_3320_),
    .Y(_3339_)
);

INVX2 _13540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2878_),
    .Y(_2879_)
);

OAI21X1 _13120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2411_),
    .C(_2408_),
    .Y(_2418_)
);

FILL SFILL3640x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4183_),
    .B(_4187_),
    .C(_4188_),
    .Y(_4198_)
);

NAND2X1 _14325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3737_),
    .B(_3738_),
    .Y(_3739_)
);

DFFPOSX1 _24003_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[57]),
    .CLK(clk_bF$buf9),
    .D(_0_[57])
);

FILL SFILL49080x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10739_),
    .B(_10735_),
    .Y(_10795_)
);

NOR2X1 _20343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10334_),
    .B(_9989_),
    .Y(_10335_)
);

AOI21X1 _19783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9417_),
    .B(_9398_),
    .C(_9420_),
    .Y(_9721_)
);

OAI21X1 _19363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .B(_9248_),
    .C(_9251_),
    .Y(_9260_)
);

AOI21X1 _21968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_90_),
    .C(_88_),
    .Y(_207_)
);

AOI22X1 _21548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf2),
    .B(breg_25_bF$buf2),
    .C(areg_19_bF$buf1),
    .D(breg_24_bF$buf0),
    .Y(_11654_)
);

AOI21X1 _21128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11177_),
    .B(_11180_),
    .C(_11183_),
    .Y(_11195_)
);

NOR2X1 _12811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10518_),
    .B(_10463_),
    .Y(_330_)
);

NAND3X1 _15283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4782_),
    .B(_4775_),
    .C(_4787_),
    .Y(_4788_)
);

FILL SFILL39080x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6106_),
    .B(_6105_),
    .C(_6097_),
    .Y(_6107_)
);

OAI21X1 _16068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5638_),
    .B(_5639_),
    .C(_5307_),
    .Y(_5648_)
);

FILL SFILL39000x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL4040x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _22086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .Y(_336_)
);

NAND3X1 _18634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8072_),
    .B(_8448_),
    .C(_8452_),
    .Y(_8461_)
);

NAND2X1 _18214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8000_),
    .B(_7999_),
    .Y(_8001_)
);

FILL SFILL29080x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf3),
    .B(areg_25_bF$buf3),
    .Y(_10856_)
);

FILL SFILL8760x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9780_),
    .B(_9781_),
    .C(_9779_),
    .Y(_9782_)
);

OAI21X1 _19419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8942_),
    .B(_8937_),
    .C(_8945_),
    .Y(_9321_)
);

NAND2X1 _14974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_14_bF$buf2),
    .Y(_4449_)
);

AOI21X1 _14554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3989_),
    .B(_3983_),
    .C(_3946_),
    .Y(_3990_)
);

INVX8 _14134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf2),
    .Y(_3529_)
);

FILL SFILL53960x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4662_),
    .B(_4989_),
    .C(_4985_),
    .Y(_5308_)
);

AND2X2 _15339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_21_bF$buf1),
    .Y(_4849_)
);

NAND3X1 _20992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11019_),
    .B(_11042_),
    .C(_11045_),
    .Y(_11046_)
);

NAND3X1 _20572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10579_),
    .B(_10585_),
    .C(_10263_),
    .Y(_10586_)
);

NOR3X1 _20152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10118_),
    .B(_10120_),
    .C(_10124_),
    .Y(_10125_)
);

OAI21X1 _16700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6338_),
    .B(_6339_),
    .C(_6337_),
    .Y(_6340_)
);

XNOR2X1 _19592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9486_),
    .B(_9511_),
    .Y(_9512_)
);

OAI21X1 _19172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_3958__bF$buf3),
    .C(_9041_),
    .Y(_9051_)
);

NAND2X1 _21777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_27_bF$buf4),
    .Y(_11905_)
);

OAI21X1 _21357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11157_),
    .B(_11140_),
    .C(_11148_),
    .Y(_11446_)
);

FILL SFILL3720x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _17905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7660_),
    .Y(_7661_)
);

FILL SFILL74360x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10123_),
    .B(_10134_),
    .C(_10101_),
    .Y(_10145_)
);

OR2X2 _12200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4083_),
    .B(_5530_),
    .Y(_5541_)
);

NOR3X1 _15092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4271_),
    .B(_4269_),
    .C(_4268_),
    .Y(_4579_)
);

NAND3X1 _13825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(_3188_),
    .C(_3096_),
    .Y(_3192_)
);

NAND3X1 _13405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2553_),
    .B(_2730_),
    .C(_2731_),
    .Y(_2732_)
);

BUFX2 _23923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[41]),
    .Y(y[41])
);

NOR2X1 _23503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1882_),
    .B(_1883_),
    .Y(_1884_)
);

NAND3X1 _16297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5889_),
    .B(_5897_),
    .C(_5898_),
    .Y(_5899_)
);

OAI21X1 _18863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_6300__bF$buf0),
    .C(_8305_),
    .Y(_8712_)
);

OAI21X1 _18443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8241_),
    .B(_8242_),
    .C(_8239_),
    .Y(_8252_)
);

XNOR2X1 _18023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7790_),
    .B(_7785_),
    .Y(_7791_)
);

FILL SFILL33880x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10645_),
    .B(_10646_),
    .C(_10346_),
    .Y(_10647_)
);

NAND2X1 _20208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10182_),
    .B(_10185_),
    .Y(_10186_)
);

OR2X2 _19648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9568_),
    .B(_9528_),
    .Y(_9573_)
);

NOR3X1 _19228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9106_),
    .B(_9108_),
    .C(_9111_),
    .Y(_9112_)
);

AOI21X1 _14783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4238_),
    .C(_4239_),
    .Y(_4240_)
);

AOI21X1 _14363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3739_),
    .B(_3741_),
    .C(_3728_),
    .Y(_3779_)
);

DFFPOSX1 _24041_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[31]),
    .CLK(clk_bF$buf9),
    .D(a[31])
);

FILL SFILL39080x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _15988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_26_bF$buf2),
    .C(breg_1_bF$buf1),
    .D(areg_25_bF$buf2),
    .Y(_5560_)
);

NAND3X1 _15568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5089_),
    .B(_5088_),
    .C(_5079_),
    .Y(_5099_)
);

NAND2X1 _15148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4636_),
    .B(_4639_),
    .Y(_4640_)
);

NOR3X1 _20381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10374_),
    .B(_10370_),
    .C(_10373_),
    .Y(_10376_)
);

FILL SFILL23880x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11691_),
    .B(_11695_),
    .C(_11646_),
    .Y(_11696_)
);

NAND2X1 _21166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf4),
    .B(areg_31_bF$buf3),
    .Y(_11237_)
);

NAND2X1 _17714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_22_bF$buf4),
    .Y(_7452_)
);

FILL FILL73960x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _18919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_31_bF$buf0),
    .Y(_8773_)
);

AOI21X1 _13634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2941_),
    .B(_2945_),
    .C(_2760_),
    .Y(_2982_)
);

NAND3X1 _13214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2517_),
    .C(_2522_),
    .Y(_2523_)
);

NAND2X1 _23732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2068_),
    .B(_2080_),
    .Y(_2133_)
);

NOR2X1 _23312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1417_),
    .B(_1675_),
    .Y(_1676_)
);

FILL SFILL53960x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4295_),
    .B(_4300_),
    .C(_4152_),
    .Y(_4301_)
);

AOI21X1 _14419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3539_),
    .B(_3559_),
    .C(_3840_),
    .Y(_3841_)
);

OAI21X1 _18672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8501_),
    .B(_8499_),
    .C(_8491_),
    .Y(_8502_)
);

OAI21X1 _18252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8025_),
    .B(_8032_),
    .C(_8035_),
    .Y(_8043_)
);

AOI21X1 _20857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10892_),
    .B(_10893_),
    .C(_10890_),
    .Y(_10898_)
);

NAND3X1 _20437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10417_),
    .B(_10422_),
    .C(_10427_),
    .Y(_10437_)
);

AOI21X1 _20017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9269_),
    .B(_9621_),
    .C(_9976_),
    .Y(_9977_)
);

FILL SFILL19000x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9818_),
    .B(_9819_),
    .C(_9820_),
    .Y(_9824_)
);

AOI21X1 _19457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8935_),
    .B(_8973_),
    .C(_9362_),
    .Y(_9363_)
);

AND2X2 _19037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_27_bF$buf2),
    .Y(_8902_)
);

XNOR2X1 _14592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .B(_3534_),
    .Y(_4032_)
);

OAI21X1 _14172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3568_),
    .B(_3570_),
    .C(_3567_),
    .Y(_3571_)
);

FILL SFILL64360x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1336_),
    .B(_1347_),
    .Y(_1358_)
);

NAND3X1 _15797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4980_),
    .B(_5346_),
    .C(_5345_),
    .Y(_5350_)
);

NAND3X1 _15377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4890_),
    .B(_4888_),
    .C(_4889_),
    .Y(_4891_)
);

OAI21X1 _20190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10161_),
    .B(_10162_),
    .C(_10165_),
    .Y(_10166_)
);

AOI21X1 _21395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11227_),
    .B(_11232_),
    .C(_11487_),
    .Y(_11488_)
);

OAI21X1 _17943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7699_),
    .B(_7698_),
    .C(_7697_),
    .Y(_7703_)
);

NAND3X1 _17523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7236_),
    .B(_7241_),
    .C(_7240_),
    .Y(_7242_)
);

NAND3X1 _17103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6756_),
    .B(_6763_),
    .C(_6766_),
    .Y(_6783_)
);

FILL SFILL33880x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8207_),
    .B(_8209_),
    .C(_8202_),
    .Y(_8563_)
);

AOI21X1 _18308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8101_),
    .B(_8102_),
    .C(_8087_),
    .Y(_8103_)
);

OAI21X1 _13863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3229_),
    .B(_3233_),
    .C(_2964_),
    .Y(_3234_)
);

DFFPOSX1 _23961_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[15]),
    .CLK(clk_bF$buf10),
    .D(_0_[15])
);

AOI21X1 _13443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2581_),
    .B(_2587_),
    .C(_2585_),
    .Y(_2773_)
);

AOI21X1 _13023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_823_),
    .B(_812_),
    .C(_790_),
    .Y(_2318_)
);

NAND2X1 _23541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1924_),
    .B(_1834_),
    .Y(_1926_)
);

NOR2X1 _23121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1455_),
    .Y(_1468_)
);

FILL SFILL8920x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4087_),
    .B(_4090_),
    .C(_4071_),
    .Y(_4091_)
);

NAND3X1 _14228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3593_),
    .B(_3631_),
    .C(_3627_),
    .Y(_3632_)
);

FILL SFILL23880x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54280x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_23_bF$buf2),
    .Y(_8294_)
);

OAI21X1 _18061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_3402__bF$buf0),
    .C(_7392_),
    .Y(_7833_)
);

FILL SFILL23800x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7651_),
    .B(_10687_),
    .C(_10684_),
    .Y(_10688_)
);

NOR2X1 _20246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10218_),
    .B(_10219_),
    .Y(_10227_)
);

FILL SFILL8840x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9602_),
    .B(_9603_),
    .C(_9276_),
    .Y(_9615_)
);

OAI21X1 _19266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_9153_),
    .C(_9142_),
    .Y(_9154_)
);

FILL SFILL13880x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11154_),
    .B(_11165_),
    .C(_11143_),
    .Y(_11176_)
);

NAND3X1 _22812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1105_),
    .B(_1128_),
    .C(_1130_),
    .Y(_1131_)
);

FILL SFILL29000x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _15186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_21_bF$buf1),
    .C(areg_2_bF$buf3),
    .D(breg_22_bF$buf2),
    .Y(_4681_)
);

FILL SFILL74440x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3256_),
    .B(_3292_),
    .C(_3293_),
    .Y(_3294_)
);

OAI21X1 _17752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_6300__bF$buf1),
    .C(_7493_),
    .Y(_7494_)
);

NAND2X1 _17332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_21_bF$buf2),
    .Y(_7034_)
);

FILL SFILL23960x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8756_),
    .B(_8762_),
    .C(_8766_),
    .Y(_8815_)
);

AOI21X1 _18537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7490_),
    .B(_8338_),
    .C(_7945_),
    .Y(_8355_)
);

AOI21X1 _18117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7891_),
    .B(_7893_),
    .C(_7889_),
    .Y(_7894_)
);

INVX1 _13672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2559_),
    .Y(_3024_)
);

AND2X2 _13252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2559_),
    .B(_2563_),
    .Y(_2564_)
);

NAND2X1 _23770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_2172_),
    .Y(_2173_)
);

NOR2X1 _23350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(_1715_),
    .Y(_1717_)
);

FILL SFILL64040x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _14877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4055_),
    .B(_4342_),
    .Y(_0_[22])
);

NAND2X1 _14457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3879_),
    .B(_3877_),
    .Y(_3883_)
);

NAND3X1 _14037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3421_),
    .B(_3422_),
    .C(_3420_),
    .Y(_3423_)
);

NOR2X1 _18290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_6815__bF$buf1),
    .Y(_8083_)
);

INVX2 _20895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10258_),
    .Y(_10940_)
);

OAI21X1 _20475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf0),
    .B(_3961__bF$buf1),
    .C(_10119_),
    .Y(_10479_)
);

OAI21X1 _20055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10017_),
    .B(_10016_),
    .C(_10007_),
    .Y(_10018_)
);

NAND2X1 _16603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_19_bF$buf5),
    .Y(_6234_)
);

NAND2X1 _19495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9403_),
    .B(_9404_),
    .Y(_9405_)
);

FILL SFILL54040x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _19075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8937_),
    .Y(_8944_)
);

AOI21X1 _17808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7550_),
    .B(_7549_),
    .C(_7548_),
    .Y(_7555_)
);

FILL SFILL18600x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1718_),
    .B(_1707_),
    .C(_1696_),
    .Y(_1772_)
);

AND2X2 _12523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_11_bF$buf1),
    .Y(_9092_)
);

NAND3X1 _12103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4368_),
    .C(_4412_),
    .Y(_4478_)
);

NAND2X1 _22621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .B(_489_),
    .Y(_922_)
);

OAI21X1 _22201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .B(_449_),
    .C(_452_),
    .Y(_463_)
);

FILL SFILL59080x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3081_),
    .B(_3080_),
    .C(_3079_),
    .Y(_3085_)
);

NAND2X1 _13308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2620_),
    .B(_2624_),
    .Y(_2625_)
);

XOR2X1 _23826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2233_),
    .B(_2219_),
    .Y(_2234_)
);

OAI21X1 _23406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1749_),
    .B(_1612_),
    .C(_1746_),
    .Y(_1778_)
);

BUFX2 BUFX2_insert400 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[22]),
    .Y(areg_22_bF$buf3)
);

BUFX2 BUFX2_insert401 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[22]),
    .Y(areg_22_bF$buf2)
);

BUFX2 BUFX2_insert402 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[22]),
    .Y(areg_22_bF$buf1)
);

BUFX2 BUFX2_insert403 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[22]),
    .Y(areg_22_bF$buf0)
);

NAND3X1 _17981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7709_),
    .B(_7743_),
    .C(_7738_),
    .Y(_7745_)
);

BUFX2 BUFX2_insert404 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf5)
);

BUFX2 BUFX2_insert405 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf4)
);

OR2X2 _17561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6857_),
    .B(_7278_),
    .Y(_7284_)
);

AND2X2 _17141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_28_bF$buf5),
    .Y(_6824_)
);

BUFX2 BUFX2_insert406 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf3)
);

BUFX2 BUFX2_insert407 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf2)
);

BUFX2 BUFX2_insert408 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf1)
);

BUFX2 BUFX2_insert409 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[19]),
    .Y(areg_19_bF$buf0)
);

NAND2X1 _18766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_21_bF$buf4),
    .Y(_8605_)
);

INVX1 _18346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8124_),
    .Y(_8145_)
);

NAND2X1 _13481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf4),
    .B(breg_9_bF$buf3),
    .Y(_2815_)
);

NOR2X1 _13061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .B(_2354_),
    .Y(_2355_)
);

OAI21X1 _14686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4131_),
    .B(_4132_),
    .C(_4128_),
    .Y(_4133_)
);

AOI22X1 _14266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_17_bF$buf1),
    .C(breg_4_bF$buf4),
    .D(areg_16_bF$buf2),
    .Y(_3674_)
);

FILL SFILL28920x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28840x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74040x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10264_),
    .B(_10268_),
    .C(_10269_),
    .Y(_10270_)
);

AOI21X1 _16832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6484_),
    .B(_6482_),
    .C(_6481_),
    .Y(_6485_)
);

NAND3X1 _16412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6003_),
    .B(_6009_),
    .C(_6011_),
    .Y(_6025_)
);

XNOR2X1 _21489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11315_),
    .B(_11590_),
    .Y(_0_[42])
);

NAND2X1 _21069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11125_),
    .B(_11129_),
    .Y(_11130_)
);

FILL SFILL64120x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _17617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf2),
    .B(_5369_),
    .Y(_7345_)
);

INVX1 _12752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9762_),
    .Y(_11592_)
);

AOI21X1 _12332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6900_),
    .B(_6834_),
    .C(_6099_),
    .Y(_6988_)
);

OAI21X1 _22850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1170_),
    .B(_1171_),
    .C(_1167_),
    .Y(_1172_)
);

NOR2X1 _22430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_712_),
    .Y(_0_[46])
);

INVX1 _22010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_251_),
    .Y(_252_)
);

FILL SFILL64040x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3323_),
    .B(_3332_),
    .C(_3333_),
    .Y(_3336_)
);

AOI21X1 _13537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2664_),
    .B(_2670_),
    .C(_2667_),
    .Y(_2876_)
);

NAND3X1 _13117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .B(_2414_),
    .C(_2409_),
    .Y(_2415_)
);

NAND2X1 _23635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1909_),
    .Y(_2028_)
);

XNOR2X1 _23215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1569_),
    .B(_1560_),
    .Y(_1570_)
);

NAND3X1 _17790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7530_),
    .B(_7534_),
    .C(_7532_),
    .Y(_7535_)
);

OAI21X1 _17370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_5921__bF$buf0),
    .C(_7069_),
    .Y(_7075_)
);

AOI21X1 _18995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8855_),
    .B(_8856_),
    .C(_8479_),
    .Y(_8857_)
);

FILL SFILL54040x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8379_),
    .B(_8381_),
    .Y(_8396_)
);

NAND2X1 _18155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7934_),
    .B(_7935_),
    .Y(_7936_)
);

NAND3X1 _13290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2590_),
    .B(_2600_),
    .C(_2603_),
    .Y(_2604_)
);

OAI21X1 _21701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11806_),
    .B(_11807_),
    .C(_11805_),
    .Y(_11823_)
);

INVX1 _14495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3918_),
    .Y(_3925_)
);

OAI21X1 _14075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3463_),
    .B(_3464_),
    .C(_3462_),
    .Y(_3465_)
);

INVX1 _12808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .Y(_297_)
);

OAI21X1 _22906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1233_),
    .C(_1101_),
    .Y(_1234_)
);

AOI21X1 _20093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10054_),
    .B(_10053_),
    .C(_10052_),
    .Y(_10060_)
);

OAI21X1 _16641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf0),
    .B(_3961__bF$buf4),
    .C(_6270_),
    .Y(_6276_)
);

AOI21X1 _16221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5798_),
    .B(_5803_),
    .C(_5782_),
    .Y(_5816_)
);

INVX1 _21298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11377_),
    .Y(_11381_)
);

NAND3X1 _17846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7589_),
    .B(_7596_),
    .C(_7343_),
    .Y(_7597_)
);

AOI21X1 _17426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6693_),
    .B(_6715_),
    .C(_7136_),
    .Y(_7137_)
);

NAND3X1 _17006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6673_),
    .B(_6675_),
    .C(_6674_),
    .Y(_6676_)
);

NOR2X1 _12981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1979_),
    .B(_2174_),
    .Y(_2185_)
);

OAI21X1 _12561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9455_),
    .B(_9444_),
    .C(_8709_),
    .Y(_9499_)
);

NAND2X1 _12141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4840_),
    .B(_4884_),
    .Y(_4895_)
);

FILL SFILL69160x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3125_),
    .B(_3121_),
    .Y(_3126_)
);

NOR2X1 _23864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2273_),
    .B(_2272_),
    .Y(_2274_)
);

NOR2X1 _13346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2665_),
    .B(_2666_),
    .Y(_2667_)
);

NAND2X1 _23444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1719_),
    .B(_1819_),
    .Y(_1820_)
);

INVX2 _23024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .Y(_1362_)
);

NAND2X1 _15912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5114_),
    .B(_5476_),
    .Y(_5477_)
);

OAI21X1 _18384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7878_),
    .B(_8186_),
    .C(_8016_),
    .Y(_8187_)
);

FILL SFILL59160x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11040_),
    .B(_11034_),
    .C(_11020_),
    .Y(_11041_)
);

OAI21X1 _20569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10577_),
    .B(_10576_),
    .C(_10561_),
    .Y(_10582_)
);

AND2X2 _20149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf4),
    .B(breg_19_bF$buf3),
    .Y(_10121_)
);

NOR3X1 _21930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_11818_),
    .C(_164_),
    .Y(_165_)
);

FILL SFILL28680x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_28_bF$buf1),
    .Y(_11613_)
);

OAI21X1 _19589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9506_),
    .B(_9507_),
    .C(_9503_),
    .Y(_9508_)
);

OAI22X1 _19169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_3958__bF$buf3),
    .C(_2560__bF$buf2),
    .D(_3402__bF$buf1),
    .Y(_9047_)
);

FILL SFILL14040x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_9_bF$buf2),
    .Y(_10112_)
);

AOI21X1 _22715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1016_),
    .B(_1010_),
    .C(_979_),
    .Y(_1025_)
);

NAND3X1 _15089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4558_),
    .B(_4562_),
    .C(_4565_),
    .Y(_4575_)
);

FILL SFILL49160x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6523_),
    .B(_6521_),
    .Y(_6526_)
);

OAI21X1 _16450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_5315__bF$buf0),
    .C(_5685_),
    .Y(_6065_)
);

NAND3X1 _16030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5599_),
    .B(_5605_),
    .C(_5463_),
    .Y(_5606_)
);

FILL SFILL18680x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _17655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf1),
    .B(_2560__bF$buf1),
    .C(_2362__bF$buf3),
    .D(_2669__bF$buf3),
    .Y(_7387_)
);

NAND2X1 _17235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_21_bF$buf0),
    .Y(_6927_)
);

NAND3X1 _12790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11866_),
    .B(_1_),
    .C(_67_),
    .Y(_100_)
);

NAND2X1 _12370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7393_),
    .B(_7371_),
    .Y(_7404_)
);

AOI21X1 _13995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3129_),
    .B(_3133_),
    .C(_3136_),
    .Y(_3377_)
);

NAND3X1 _13575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2916_),
    .B(_2917_),
    .C(_2915_),
    .Y(_2918_)
);

INVX2 _13155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .Y(_2458_)
);

INVX1 _23673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .Y(_2069_)
);

NAND3X1 _23253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1611_),
    .C(_1606_),
    .Y(_1612_)
);

NAND3X1 _19801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9737_),
    .B(_9738_),
    .C(_9739_),
    .Y(_9741_)
);

DFFPOSX1 _24038_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[28]),
    .CLK(clk_bF$buf4),
    .D(a[28])
);

AOI21X1 _15721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5249_),
    .B(_5255_),
    .C(_5008_),
    .Y(_5268_)
);

AND2X2 _15301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4475_),
    .B(_4468_),
    .Y(_4808_)
);

AOI21X1 _18193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7976_),
    .B(_7977_),
    .C(_7974_),
    .Y(_7978_)
);

AOI21X1 _20798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10832_),
    .B(_10830_),
    .C(_10829_),
    .Y(_10833_)
);

OAI21X1 _20378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf1),
    .B(_5668__bF$buf0),
    .C(_10359_),
    .Y(_10372_)
);

OAI21X1 _16926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6251_),
    .B(_6258_),
    .C(_6260_),
    .Y(_6588_)
);

NOR2X1 _16506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6122_),
    .B(_6126_),
    .Y(_6127_)
);

FILL SFILL69240x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8900_),
    .B(_8904_),
    .C(_8908_),
    .Y(_9298_)
);

FILL SFILL38760x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .B(_703_),
    .C(_691_),
    .Y(_713_)
);

AOI21X1 _12426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6769_),
    .B(_6341_),
    .C(_6802_),
    .Y(_8029_)
);

NAND2X1 _22944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf4),
    .B(breg_28_bF$buf3),
    .Y(_1275_)
);

NAND3X1 _12006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg[0]),
    .C(_2738_),
    .Y(_3416_)
);

NAND3X1 _22524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_772_),
    .B(_810_),
    .C(_815_),
    .Y(_816_)
);

AOI21X1 _22104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_351_),
    .C(_349_),
    .Y(_356_)
);

FILL SFILL3800x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _23729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2090_),
    .C(_2128_),
    .Y(_2129_)
);

NOR2X1 _23309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf2),
    .B(_6815__bF$buf4),
    .Y(_1672_)
);

FILL SFILL59240x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74200x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _17884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7215_),
    .B(_7638_),
    .Y(_0_[31])
);

NOR3X1 _17464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6753_),
    .B(_6754_),
    .C(_6752_),
    .Y(_7178_)
);

OAI21X1 _17044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6713_),
    .B(_6712_),
    .C(_6694_),
    .Y(_6718_)
);

FILL SFILL28760x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_27_bF$buf2),
    .Y(_8498_)
);

NAND3X1 _18249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8036_),
    .B(_8037_),
    .C(_8035_),
    .Y(_8038_)
);

NAND3X1 _13384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2697_),
    .C(_2699_),
    .Y(_2709_)
);

NAND2X1 _23482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1776_),
    .B(_1861_),
    .Y(_1862_)
);

INVX1 _23062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .Y(_1403_)
);

INVX2 _19610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9530_),
    .Y(_9531_)
);

NAND3X1 _14589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4012_),
    .B(_4016_),
    .C(_3866_),
    .Y(_4028_)
);

AOI21X1 _14169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3260_),
    .B(_3278_),
    .C(_3282_),
    .Y(_3567_)
);

FILL SFILL18760x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_20_bF$buf1),
    .Y(_5518_)
);

OAI22X1 _15530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4451_),
    .B(_5055_),
    .C(_5056_),
    .D(_4770_),
    .Y(_5057_)
);

NAND3X1 _15110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4592_),
    .B(_4597_),
    .C(_4444_),
    .Y(_4598_)
);

NOR2X1 _20187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9811_),
    .B(_9858_),
    .Y(_10163_)
);

NOR3X1 _16735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5985_),
    .B(_5986_),
    .C(_5984_),
    .Y(_6379_)
);

NAND2X1 _16315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_24_bF$buf2),
    .Y(_5919_)
);

XOR2X1 _12655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10518_),
    .B(_10463_),
    .Y(_10529_)
);

AOI22X1 _12235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5804_),
    .B(_5848_),
    .C(_4895_),
    .D(_3953_),
    .Y(_5925_)
);

AOI21X1 _22753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .B(_1026_),
    .C(_950_),
    .Y(_1067_)
);

NAND3X1 _22333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_605_),
    .C(_606_),
    .Y(_607_)
);

DFFPOSX1 _23958_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[12]),
    .CLK(clk_bF$buf2),
    .D(_0_[12])
);

OR2X2 _23538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1916_),
    .B(_1917_),
    .Y(_1922_)
);

NAND3X1 _23118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1463_),
    .C(_1460_),
    .Y(_1464_)
);

NAND3X1 _14801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4241_),
    .B(_4257_),
    .C(_4253_),
    .Y(_4260_)
);

NAND3X1 _17693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7422_),
    .B(_7344_),
    .C(_7428_),
    .Y(_7429_)
);

NAND3X1 _17273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6962_),
    .B(_6968_),
    .C(_6965_),
    .Y(_6969_)
);

NAND3X1 _18898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8746_),
    .B(_8749_),
    .C(_8748_),
    .Y(_8750_)
);

NAND2X1 _18478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf2),
    .B(areg_22_bF$buf4),
    .Y(_8290_)
);

OAI21X1 _18058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_2884__bF$buf3),
    .C(_7818_),
    .Y(_7829_)
);

OAI21X1 _13193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2499_),
    .B(_2498_),
    .C(_2496_),
    .Y(_2500_)
);

XNOR2X1 _23291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1652_),
    .Y(_0_[52])
);

NAND2X1 _11926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf3),
    .B(areg_4_bF$buf4),
    .Y(_2540_)
);

INVX1 _21604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11541_),
    .Y(_11716_)
);

OAI21X1 _14398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3542_),
    .B(_3817_),
    .C(_3815_),
    .Y(_3818_)
);

OAI21X1 _22809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1126_),
    .C(_1106_),
    .Y(_1127_)
);

NAND3X1 _16964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6622_),
    .B(_6629_),
    .C(_6609_),
    .Y(_6630_)
);

AND2X2 _16544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_15_bF$buf3),
    .Y(_6169_)
);

AOI21X1 _16124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5699_),
    .B(_5690_),
    .C(_5675_),
    .Y(_5709_)
);

AND2X2 _17749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .B(areg_25_bF$buf0),
    .Y(_7490_)
);

NAND2X1 _17329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7027_),
    .B(_7028_),
    .Y(_7029_)
);

AOI21X1 _12884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(_965_),
    .C(_11668_),
    .Y(_1129_)
);

NAND3X1 _12464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6955_),
    .B(_8260_),
    .C(_8271_),
    .Y(_8435_)
);

NAND2X1 _22982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1311_),
    .B(_1315_),
    .Y(_1316_)
);

OAI21X1 _12044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3810_),
    .B(_3821_),
    .C(_3558_),
    .Y(_3832_)
);

OAI21X1 _22562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_7100__bF$buf1),
    .C(_855_),
    .Y(_858_)
);

AOI21X1 _22142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_395_),
    .B(_397_),
    .C(_394_),
    .Y(_398_)
);

FILL SFILL33960x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3018_),
    .B(_3010_),
    .C(_3019_),
    .Y(_3020_)
);

NAND2X1 _23767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2148_),
    .B(_2147_),
    .Y(_2170_)
);

INVX8 _13249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .Y(_2560_)
);

XOR2X1 _23347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .B(_1710_),
    .Y(_1714_)
);

FILL SFILL18760x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4045_),
    .B(_4049_),
    .Y(_4050_)
);

NAND2X1 _17082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6757_),
    .B(_6759_),
    .Y(_6760_)
);

FILL SFILL74280x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5369_),
    .Y(_5370_)
);

NOR2X1 _18287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf0),
    .B(_7225__bF$buf3),
    .Y(_8080_)
);

FILL SFILL23960x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_48_),
    .C(_28_),
    .Y(_59_)
);

NOR2X1 _21413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11465_),
    .B(_11470_),
    .Y(_11508_)
);

OAI21X1 _22618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_917_),
    .C(_918_),
    .Y(_919_)
);

OAI21X1 _16773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6402_),
    .B(_6400_),
    .C(_6392_),
    .Y(_6420_)
);

NAND3X1 _16353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5954_),
    .B(_5912_),
    .C(_5960_),
    .Y(_5961_)
);

BUFX2 BUFX2_insert370 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf4)
);

BUFX2 BUFX2_insert371 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf3)
);

BUFX2 BUFX2_insert372 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf2)
);

BUFX2 BUFX2_insert373 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf1)
);

NOR3X1 _17978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7367_),
    .B(_7365_),
    .C(_7361_),
    .Y(_7741_)
);

BUFX2 BUFX2_insert374 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf0)
);

OAI21X1 _17558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7279_),
    .B(_7277_),
    .C(_7276_),
    .Y(_7280_)
);

BUFX2 BUFX2_insert375 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .Y(_2560__bF$buf4)
);

NAND2X1 _17138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg_29_bF$buf0),
    .Y(_6820_)
);

BUFX2 BUFX2_insert376 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .Y(_2560__bF$buf3)
);

BUFX2 BUFX2_insert377 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .Y(_2560__bF$buf2)
);

BUFX2 BUFX2_insert378 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .Y(_2560__bF$buf1)
);

NAND3X1 _12693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10891_),
    .B(_10803_),
    .C(_10935_),
    .Y(_10946_)
);

BUFX2 BUFX2_insert379 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560_),
    .Y(_2560__bF$buf0)
);

AND2X2 _12273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6286_),
    .B(_6330_),
    .Y(_6341_)
);

NAND3X1 _22791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(_967_),
    .C(_958_),
    .Y(_1108_)
);

XOR2X1 _22371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_647_),
    .B(_643_),
    .Y(_649_)
);

AOI21X1 _13898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3051_),
    .B(_3270_),
    .C(_3054_),
    .Y(_3271_)
);

NAND2X1 _13478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2805_),
    .B(_2810_),
    .Y(_2811_)
);

DFFPOSX1 _23996_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[50]),
    .CLK(clk_bF$buf6),
    .D(_0_[50])
);

NAND2X1 _13058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(_2349_),
    .Y(_2353_)
);

AOI21X1 _23576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3766_),
    .B(_3769_),
    .C(_4050_),
    .Y(_1963_)
);

AOI21X1 _23156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1483_),
    .B(_1488_),
    .C(_1408_),
    .Y(_1506_)
);

OAI21X1 _19704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9632_),
    .B(_9630_),
    .C(_9633_),
    .Y(_9634_)
);

FILL SFILL33720x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49320x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf3),
    .B(_3146__bF$buf0),
    .C(_5156_),
    .Y(_5161_)
);

AOI21X1 _15204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4692_),
    .B(_4691_),
    .C(_4687_),
    .Y(_4701_)
);

NAND3X1 _18096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7869_),
    .B(_7868_),
    .C(_7870_),
    .Y(_7871_)
);

NAND2X1 _16829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6073_),
    .B(_6081_),
    .Y(_6481_)
);

NAND3X1 _16409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6016_),
    .B(_5665_),
    .C(_6020_),
    .Y(_6021_)
);

OAI21X1 _11964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2924_),
    .B(_2946_),
    .C(_2901_),
    .Y(_2957_)
);

AND2X2 _21642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_27_bF$buf0),
    .Y(_11758_)
);

OAI21X1 _21222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11285_),
    .B(_11289_),
    .C(_11292_),
    .Y(_11299_)
);

AOI21X1 _12749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11417_),
    .B(_11483_),
    .C(_9959_),
    .Y(_11560_)
);

NAND3X1 _12329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6911_),
    .B(_6034_),
    .C(_6944_),
    .Y(_6955_)
);

NAND2X1 _22847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1156_),
    .B(_1154_),
    .Y(_1169_)
);

OAI21X1 _22427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11879_),
    .B(_709_),
    .C(_488_),
    .Y(_710_)
);

OAI21X1 _22007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_211_),
    .C(_194_),
    .Y(_249_)
);

NOR3X1 _16582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6210_),
    .B(_6208_),
    .C(_6207_),
    .Y(_6211_)
);

XOR2X1 _16162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5688_),
    .B(_5750_),
    .Y(_5751_)
);

NAND2X1 _17787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7111_),
    .B(_7531_),
    .Y(_7532_)
);

OAI22X1 _17367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_5921__bF$buf0),
    .C(_4116__bF$buf0),
    .D(_4541__bF$buf3),
    .Y(_7072_)
);

INVX8 _12082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf0),
    .Y(_4258_)
);

NAND3X1 _22180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .B(_438_),
    .C(_433_),
    .Y(_439_)
);

FILL SFILL8680x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10602_),
    .B(_10614_),
    .C(_10959_),
    .Y(_10960_)
);

FILL SFILL13640x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .Y(_2601_)
);

NAND3X1 _23385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1623_),
    .B(_1742_),
    .C(_1746_),
    .Y(_1756_)
);

FILL SFILL69000x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _19933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9859_),
    .B(_9885_),
    .Y(_9886_)
);

OAI21X1 _19513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9075_),
    .B(_9042_),
    .C(_9067_),
    .Y(_9425_)
);

FILL SFILL74280x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_15_bF$buf5),
    .Y(_5412_)
);

NAND3X1 _15433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4932_),
    .B(_4936_),
    .C(_4940_),
    .Y(_4953_)
);

OAI21X1 _15013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4485_),
    .B(_4486_),
    .C(_4487_),
    .Y(_4492_)
);

OAI22X1 _16638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_4551__bF$buf1),
    .C(_4116__bF$buf0),
    .D(_3961__bF$buf2),
    .Y(_6272_)
);

NAND3X1 _16218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5802_),
    .B(_5789_),
    .C(_5794_),
    .Y(_5812_)
);

NOR2X1 _21871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_99_),
    .Y(_101_)
);

NAND3X1 _21451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11547_),
    .B(_11546_),
    .C(_11548_),
    .Y(_11550_)
);

AOI21X1 _21031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10837_),
    .B(_10841_),
    .C(_10821_),
    .Y(_11089_)
);

FILL SFILL64280x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf0),
    .B(_6582__bF$buf3),
    .Y(_2153_)
);

OAI21X1 _12558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9455_),
    .B(_9444_),
    .C(_9433_),
    .Y(_9466_)
);

NAND3X1 _12138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3449_),
    .B(_4785_),
    .C(_4697_),
    .Y(_4862_)
);

OAI21X1 _22656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf3),
    .B(_5668__bF$buf1),
    .C(_742_),
    .Y(_960_)
);

OAI21X1 _22236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_365_),
    .C(_448_),
    .Y(_500_)
);

FILL SFILL64200x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5999_),
    .B(_6000_),
    .C(_5998_),
    .Y(_6002_)
);

AOI21X1 _14704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .B(_4002_),
    .C(_3915_),
    .Y(_4153_)
);

NAND2X1 _17596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7269_),
    .B(_7266_),
    .Y(_7322_)
);

OAI21X1 _17176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6861_),
    .B(_6860_),
    .C(_6851_),
    .Y(_6862_)
);

NAND2X1 _15909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf1),
    .B(areg_15_bF$buf2),
    .Y(_5473_)
);

OAI21X1 _20722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10749_),
    .B(_10747_),
    .C(_10744_),
    .Y(_10750_)
);

OAI21X1 _20302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10287_),
    .B(_10289_),
    .C(_10284_),
    .Y(_10290_)
);

NAND2X1 _13096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_10_bF$buf3),
    .Y(_2393_)
);

AOI21X1 _23194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1546_),
    .B(_942_),
    .C(_1545_),
    .Y(_1547_)
);

NAND3X1 _19742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9649_),
    .B(_9673_),
    .C(_9675_),
    .Y(_9676_)
);

NAND3X1 _19322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9209_),
    .B(_9210_),
    .C(_9208_),
    .Y(_9216_)
);

NAND3X1 _21927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_158_),
    .C(_127_),
    .Y(_162_)
);

OAI21X1 _21507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11343_),
    .B(_11334_),
    .C(_11338_),
    .Y(_11610_)
);

NAND2X1 _15662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_25_bF$buf2),
    .Y(_5203_)
);

OAI21X1 _15242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4727_),
    .B(_4728_),
    .C(_4725_),
    .Y(_4743_)
);

AND2X2 _16867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_19_bF$buf1),
    .Y(_6523_)
);

AND2X2 _16447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_25_bF$buf3),
    .Y(_6062_)
);

OAI21X1 _16027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5595_),
    .B(_5597_),
    .C(_5513_),
    .Y(_5603_)
);

NAND3X1 _21680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11718_),
    .B(_11794_),
    .C(_11798_),
    .Y(_11799_)
);

OAI21X1 _21260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf4),
    .B(_5668__bF$buf5),
    .C(_11030_),
    .Y(_11339_)
);

FILL SFILL8600x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_23_),
    .Y(_67_)
);

XNOR2X1 _12367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7360_),
    .B(_7327_),
    .Y(_7371_)
);

NAND2X1 _22885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1210_),
    .Y(_1211_)
);

INVX1 _22465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .Y(_751_)
);

NAND3X1 _22045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_282_),
    .C(_279_),
    .Y(_291_)
);

FILL SFILL74280x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4403_),
    .B(_4402_),
    .C(_4392_),
    .Y(_4404_)
);

OAI21X1 _14513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3943_),
    .B(_3944_),
    .C(_3941_),
    .Y(_3945_)
);

FILL SFILL74200x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5263_),
    .B(_5007_),
    .C(_5257_),
    .Y(_5264_)
);

NAND2X1 _20951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10995_),
    .B(_10996_),
    .Y(_11001_)
);

AOI21X1 _20531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10238_),
    .B(_10243_),
    .C(_10246_),
    .Y(_10541_)
);

NOR3X1 _20111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10073_),
    .B(_10074_),
    .C(_10075_),
    .Y(_10080_)
);

AOI21X1 _19971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9562_),
    .B(_9924_),
    .C(_9925_),
    .Y(_9927_)
);

OAI21X1 _19551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9450_),
    .B(_9454_),
    .C(_9457_),
    .Y(_9467_)
);

NAND2X1 _19131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8677_),
    .B(_8682_),
    .Y(_9006_)
);

AOI21X1 _21736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11319_),
    .B(_11581_),
    .C(_11860_),
    .Y(_11861_)
);

AOI21X1 _21316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11396_),
    .B(_11397_),
    .C(_11394_),
    .Y(_11401_)
);

FILL SFILL28840x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5104_),
    .B(_5144_),
    .C(_5141_),
    .Y(_5454_)
);

AND2X2 _15471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4665_),
    .B(_4657_),
    .Y(_4993_)
);

AOI21X1 _15051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4530_),
    .B(_4531_),
    .C(_4532_),
    .Y(_4534_)
);

AOI22X1 _16676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_28_bF$buf4),
    .C(breg_1_bF$buf1),
    .D(areg_27_bF$buf4),
    .Y(_6314_)
);

NAND2X1 _16256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_18_bF$buf0),
    .Y(_5854_)
);

FILL SFILL54200x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9828_),
    .B(_9872_),
    .Y(_9883_)
);

OAI21X1 _12176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5267_),
    .B(_5256_),
    .C(_5113_),
    .Y(_5278_)
);

AOI21X1 _22694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1000_),
    .B(_861_),
    .C(_1001_),
    .Y(_1002_)
);

OAI21X1 _22274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_541_),
    .C(_327_),
    .Y(_542_)
);

OAI21X1 _18822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8661_),
    .B(_8666_),
    .C(_8636_),
    .Y(_8667_)
);

AOI21X1 _18402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8206_),
    .B(_8204_),
    .C(_8203_),
    .Y(_8207_)
);

BUFX2 _23899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[17]),
    .Y(y[17])
);

AOI21X1 _23479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(_1845_),
    .C(_1778_),
    .Y(_1858_)
);

OAI21X1 _23059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1387_),
    .B(_1390_),
    .C(_1393_),
    .Y(_1399_)
);

NAND2X1 _19607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9523_),
    .B(_9527_),
    .Y(_9528_)
);

OAI21X1 _14742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4194_),
    .B(_4189_),
    .C(_4155_),
    .Y(_4195_)
);

NOR3X1 _14322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3728_),
    .B(_3590_),
    .C(_3735_),
    .Y(_3736_)
);

DFFPOSX1 _24000_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[54]),
    .CLK(clk_bF$buf6),
    .D(_0_[54])
);

OAI21X1 _15947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5151_),
    .B(_5514_),
    .C(_5160_),
    .Y(_5515_)
);

NAND3X1 _15527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5044_),
    .B(_5052_),
    .C(_5053_),
    .Y(_5054_)
);

AOI21X1 _15107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4590_),
    .B(_4589_),
    .C(_4587_),
    .Y(_4595_)
);

AOI21X1 _20760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10779_),
    .B(_10774_),
    .C(_10742_),
    .Y(_10791_)
);

OAI21X1 _20340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10326_),
    .B(_10327_),
    .C(_10325_),
    .Y(_10331_)
);

FILL SFILL13720x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9711_),
    .B(_9715_),
    .C(_9716_),
    .Y(_9717_)
);

AOI22X1 _19360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8869_),
    .B(_8875_),
    .C(_9249_),
    .D(_9254_),
    .Y(_9256_)
);

OAI21X1 _21965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .B(_182_),
    .C(_180_),
    .Y(_204_)
);

NAND2X1 _21545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf2),
    .B(breg_25_bF$buf2),
    .Y(_11651_)
);

NAND3X1 _21125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11169_),
    .B(_11184_),
    .C(_11191_),
    .Y(_11192_)
);

NOR2X1 _15280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4463_),
    .B(_4783_),
    .Y(_4784_)
);

FILL SFILL3960x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5673_),
    .B(_5711_),
    .C(_6103_),
    .Y(_6104_)
);

OAI21X1 _16065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5643_),
    .B(_5644_),
    .C(_5305_),
    .Y(_5645_)
);

FILL SFILL3480x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_124_),
    .C(_332_),
    .Y(_333_)
);

OAI21X1 _18631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8453_),
    .B(_8456_),
    .C(_8070_),
    .Y(_8458_)
);

AOI21X1 _18211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7991_),
    .B(_7996_),
    .C(_7926_),
    .Y(_7998_)
);

NAND2X1 _20816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf3),
    .B(areg_23_bF$buf1),
    .Y(_10853_)
);

FILL SFILL28840x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1648_),
    .B(_1649_),
    .C(_1550_),
    .Y(_1650_)
);

FILL SFILL33800x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9402_),
    .B(_9406_),
    .C(_9409_),
    .Y(_9779_)
);

AOI21X1 _19416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8959_),
    .B(_8964_),
    .C(_8966_),
    .Y(_9318_)
);

AOI21X1 _14971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_4273_),
    .C(_4202_),
    .Y(_4446_)
);

NAND3X1 _14551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3981_),
    .B(_3980_),
    .C(_3979_),
    .Y(_3987_)
);

INVX4 _14131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf3),
    .Y(_3526_)
);

AOI21X1 _15756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4669_),
    .B(_5001_),
    .C(_5304_),
    .Y(_5305_)
);

AOI21X1 _15336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4543_),
    .B(_4548_),
    .C(_4536_),
    .Y(_4846_)
);

FILL SFILL54200x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_28_bF$buf1),
    .Y(_11902_)
);

OAI21X1 _21354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf3),
    .B(_3781__bF$buf3),
    .C(_11135_),
    .Y(_11443_)
);

AOI21X1 _17902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7604_),
    .B(_7610_),
    .C(_7223_),
    .Y(_7658_)
);

FILL SFILL38920x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1202_),
    .B(_1211_),
    .Y(_1312_)
);

OAI21X1 _22559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253__bF$buf0),
    .B(_7520__bF$buf1),
    .C(_853_),
    .Y(_854_)
);

XNOR2X1 _22139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_393_),
    .Y(_394_)
);

NAND3X1 _13822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(_3188_),
    .C(_3183_),
    .Y(_3189_)
);

BUFX2 _23920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[38]),
    .Y(y[38])
);

NAND3X1 _13402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2722_),
    .C(_2728_),
    .Y(_2729_)
);

NAND2X1 _23500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_27_bF$buf1),
    .B(breg_27_bF$buf0),
    .Y(_1880_)
);

NAND3X1 _16294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5890_),
    .B(_5895_),
    .C(_5894_),
    .Y(_5896_)
);

FILL SFILL48920x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4036_),
    .B(_4040_),
    .C(_3763_),
    .Y(_4047_)
);

OAI21X1 _17499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6808_),
    .B(_7214_),
    .C(_7209_),
    .Y(_7215_)
);

NAND3X1 _17079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6750_),
    .B(_6755_),
    .C(_6600_),
    .Y(_6756_)
);

AOI21X1 _18860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8705_),
    .B(_8707_),
    .C(_8703_),
    .Y(_8708_)
);

INVX1 _18440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7823_),
    .Y(_8248_)
);

NOR2X1 _18020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7721_),
    .B(_7786_),
    .Y(_7787_)
);

NAND3X1 _20625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10345_),
    .B(_10637_),
    .C(_10638_),
    .Y(_10644_)
);

NOR3X1 _20205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10131_),
    .B(_10129_),
    .C(_10125_),
    .Y(_10183_)
);

OAI21X1 _23097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1144_),
    .B(_1301_),
    .C(_1307_),
    .Y(_1441_)
);

AND2X2 _19645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9568_),
    .B(_9528_),
    .Y(_9570_)
);

AND2X2 _19225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_25_bF$buf4),
    .Y(_9109_)
);

NAND2X1 _14780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg_17_bF$buf1),
    .Y(_4236_)
);

OAI21X1 _14360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3759_),
    .B(_3521_),
    .C(_3750_),
    .Y(_3775_)
);

INVX2 _15985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5556_),
    .Y(_5557_)
);

OAI21X1 _15565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5095_),
    .B(_5090_),
    .C(_5009_),
    .Y(_5096_)
);

OAI21X1 _15145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4633_),
    .B(_4634_),
    .C(_4348_),
    .Y(_4637_)
);

AOI21X1 _21583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11688_),
    .B(_11687_),
    .C(_11686_),
    .Y(_11693_)
);

XNOR2X1 _21163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11233_),
    .B(_11227_),
    .Y(_11234_)
);

FILL SFILL28920x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7446_),
    .B(_7447_),
    .Y(_7449_)
);

NAND2X1 _22788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1010_),
    .B(_1017_),
    .Y(_1104_)
);

OR2X2 _22368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_405_),
    .B(_644_),
    .Y(_645_)
);

AOI21X1 _18916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8377_),
    .B(_8376_),
    .C(_8375_),
    .Y(_8770_)
);

OR2X2 _13631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2974_),
    .B(_2750_),
    .Y(_2979_)
);

AOI21X1 _13211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .B(_2515_),
    .C(_2373_),
    .Y(_2520_)
);

FILL SFILL18920x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4291_),
    .B(_4293_),
    .C(_4290_),
    .Y(_4298_)
);

NAND3X1 _14416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3833_),
    .B(_3808_),
    .C(_3837_),
    .Y(_3838_)
);

FILL SFILL18680x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10579_),
    .B(_10585_),
    .C(_10263_),
    .Y(_10895_)
);

OAI21X1 _20434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10432_),
    .B(_10433_),
    .C(_10431_),
    .Y(_10434_)
);

AOI21X1 _20014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9972_),
    .B(_9973_),
    .C(_9637_),
    .Y(_9974_)
);

AOI21X1 _19874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9819_),
    .B(_9820_),
    .C(_9818_),
    .Y(_9821_)
);

NAND3X1 _19454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9319_),
    .B(_9354_),
    .C(_9359_),
    .Y(_9360_)
);

NAND2X1 _19034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg_29_bF$buf3),
    .Y(_8899_)
);

NAND2X1 _21639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_27_bF$buf0),
    .Y(_11754_)
);

NAND3X1 _21219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11293_),
    .B(_11294_),
    .C(_11292_),
    .Y(_11295_)
);

AOI21X1 _12902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11538_),
    .B(_11571_),
    .C(_9762_),
    .Y(_1325_)
);

AOI21X1 _15794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5346_),
    .B(_5345_),
    .C(_4980_),
    .Y(_5347_)
);

NAND2X1 _15374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4886_),
    .B(_4887_),
    .Y(_4888_)
);

FILL SFILL69080x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6657_),
    .B(_6656_),
    .C(_6653_),
    .Y(_6668_)
);

AOI21X1 _16579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6202_),
    .B(_6203_),
    .C(_6201_),
    .Y(_6207_)
);

NAND2X1 _16159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_23_bF$buf0),
    .Y(_5747_)
);

OAI21X1 _21392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_7100__bF$buf0),
    .C(_11474_),
    .Y(_11485_)
);

NOR3X1 _17940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7684_),
    .B(_7670_),
    .C(_7691_),
    .Y(_7699_)
);

AND2X2 _17520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_27_bF$buf0),
    .Y(_7238_)
);

NOR3X1 _17100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6381_),
    .B(_6382_),
    .C(_6380_),
    .Y(_6779_)
);

INVX1 _12499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8775_),
    .Y(_8819_)
);

INVX2 _12079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4204_),
    .Y(_4215_)
);

NAND2X1 _22597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_886_),
    .Y(_896_)
);

OAI21X1 _22177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_430_),
    .C(_399_),
    .Y(_436_)
);

NAND3X1 _18725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8552_),
    .B(_8557_),
    .C(_8559_),
    .Y(_8560_)
);

AOI21X1 _18305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7673_),
    .B(_7677_),
    .C(_7681_),
    .Y(_8100_)
);

NAND3X1 _13860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3226_),
    .B(_2983_),
    .C(_3227_),
    .Y(_3230_)
);

OAI21X1 _13440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf1),
    .B(_2362__bF$buf0),
    .C(_2558_),
    .Y(_2769_)
);

NAND3X1 _13020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2299_),
    .B(_2142_),
    .C(_2304_),
    .Y(_2315_)
);

FILL SFILL3640x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4085_),
    .B(_4084_),
    .C(_4082_),
    .Y(_4088_)
);

NAND3X1 _14225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3618_),
    .B(_3611_),
    .C(_3598_),
    .Y(_3629_)
);

NAND2X1 _20663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10673_),
    .B(_9987_),
    .Y(_10685_)
);

NAND3X1 _20243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10217_),
    .B(_10223_),
    .C(_10220_),
    .Y(_10224_)
);

FILL SFILL28920x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8887_),
    .B(_9235_),
    .C(_9611_),
    .Y(_9612_)
);

NAND3X1 _19263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9145_),
    .B(_9150_),
    .C(_9147_),
    .Y(_9151_)
);

FILL SFILL49000x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf2),
    .B(areg_23_bF$buf0),
    .Y(_97_)
);

INVX2 _21448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11258_),
    .Y(_11546_)
);

NAND3X1 _21028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11081_),
    .B(_11067_),
    .C(_11071_),
    .Y(_11085_)
);

AND2X2 _12711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10639_),
    .B(_10682_),
    .Y(_11143_)
);

NAND2X1 _15183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_23_bF$buf3),
    .Y(_4678_)
);

FILL SFILL39080x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3257_),
    .B(_3286_),
    .C(_3290_),
    .Y(_3291_)
);

AOI21X1 _16388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5612_),
    .B(_5461_),
    .C(_5997_),
    .Y(_5998_)
);

FILL SFILL39000x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8770_),
    .B(_7968_),
    .C(_8777_),
    .Y(_8812_)
);

INVX1 _18534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8347_),
    .Y(_8352_)
);

OAI21X1 _18114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf4),
    .B(_4551__bF$buf1),
    .C(_7890_),
    .Y(_7891_)
);

NAND2X1 _20719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf0),
    .B(breg_24_bF$buf1),
    .Y(_10746_)
);

FILL SFILL8760x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9671_),
    .B(_9665_),
    .C(_9650_),
    .Y(_9672_)
);

OAI21X1 _19319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9205_),
    .B(_9211_),
    .C(_9004_),
    .Y(_9212_)
);

AOI21X1 _14874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4327_),
    .B(_4330_),
    .C(_4056_),
    .Y(_4340_)
);

OAI21X1 _14454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_10869__bF$buf3),
    .C(_3879_),
    .Y(_3880_)
);

XNOR2X1 _14034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3393_),
    .B(_3387_),
    .Y(_3420_)
);

AOI22X1 _15659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_25_bF$buf3),
    .C(breg_1_bF$buf4),
    .D(areg_24_bF$buf4),
    .Y(_5199_)
);

NAND3X1 _15239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4734_),
    .B(_4738_),
    .C(_4710_),
    .Y(_4739_)
);

NAND3X1 _20892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10928_),
    .B(_10922_),
    .C(_10926_),
    .Y(_10937_)
);

AOI21X1 _20472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10472_),
    .B(_10475_),
    .C(_10470_),
    .Y(_10476_)
);

NAND2X1 _20052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_27_bF$buf2),
    .Y(_10015_)
);

FILL SFILL74360x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5850_),
    .B(_6229_),
    .Y(_6230_)
);

INVX2 _19492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9401_),
    .Y(_9402_)
);

NOR2X1 _19072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8938_),
    .B(_8940_),
    .Y(_8941_)
);

XNOR2X1 _11999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3329_),
    .B(_3044_),
    .Y(_0_[5])
);

OAI21X1 _21677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11791_),
    .B(_11792_),
    .C(_11753_),
    .Y(_11796_)
);

AND2X2 _21257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_28_bF$buf1),
    .Y(_11336_)
);

FILL SFILL3720x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7513_),
    .B(_7551_),
    .C(_7546_),
    .Y(_7552_)
);

NOR2X1 _12940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_232_),
    .B(_210_),
    .Y(_1740_)
);

NAND2X1 _12520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf3),
    .B(areg_9_bF$buf1),
    .Y(_9049_)
);

OAI21X1 _12100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_4434__bF$buf2),
    .C(_3635_),
    .Y(_4445_)
);

FILL SFILL3640x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3080_),
    .B(_3081_),
    .C(_3079_),
    .Y(_3082_)
);

NOR3X1 _13305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2613_),
    .B(_2614_),
    .C(_2618_),
    .Y(_2622_)
);

AND2X2 _23823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2230_),
    .Y(_2231_)
);

AOI21X1 _23403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1753_),
    .C(_1760_),
    .Y(_1775_)
);

OAI21X1 _16197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf0),
    .B(_2362__bF$buf1),
    .C(_5781_),
    .Y(_5788_)
);

FILL SFILL49080x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8264_),
    .B(_8269_),
    .Y(_8602_)
);

NOR3X1 _18343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8125_),
    .B(_8129_),
    .C(_8130_),
    .Y(_8142_)
);

NAND2X1 _20948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10997_),
    .B(_10993_),
    .Y(_10998_)
);

OAI21X1 _20528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10532_),
    .B(_10533_),
    .C(_10497_),
    .Y(_10537_)
);

OAI21X1 _20108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10073_),
    .B(_10074_),
    .C(_10075_),
    .Y(_10076_)
);

OAI21X1 _19968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9917_),
    .B(_9922_),
    .C(_9855_),
    .Y(_9923_)
);

AOI21X1 _19548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9456_),
    .B(_9462_),
    .C(_9424_),
    .Y(_9463_)
);

NAND2X1 _19128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8997_),
    .B(_9001_),
    .Y(_9002_)
);

OAI21X1 _14683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4118_),
    .B(_4119_),
    .C(_4112_),
    .Y(_4130_)
);

AND2X2 _14263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_16_bF$buf2),
    .Y(_3671_)
);

AOI21X1 _15888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .B(_5444_),
    .C(_5449_),
    .Y(_5450_)
);

OR2X2 _15468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4984_),
    .B(_4982_),
    .Y(_4989_)
);

AND2X2 _15048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_19_bF$buf0),
    .Y(_4530_)
);

OAI21X1 _20281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10250_),
    .B(_10254_),
    .C(_10265_),
    .Y(_10267_)
);

FILL SFILL23880x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54280x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11320_),
    .B(_11570_),
    .C(_11578_),
    .Y(_11588_)
);

NAND3X1 _21066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11115_),
    .B(_11111_),
    .C(_11123_),
    .Y(_11127_)
);

AOI21X1 _17614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7156_),
    .B(_7162_),
    .C(_7015_),
    .Y(_7342_)
);

FILL SFILL8760x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8646_),
    .B(_8649_),
    .C(_8659_),
    .Y(_8663_)
);

NOR2X1 _13954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3325_),
    .B(_3326_),
    .Y(_3333_)
);

NAND2X1 _13534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_14_bF$buf4),
    .Y(_2873_)
);

AND2X2 _13114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1968_),
    .B(_1990_),
    .Y(_2412_)
);

AND2X2 _23632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .B(_2021_),
    .Y(_2025_)
);

OAI21X1 _23212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1563_),
    .B(_1564_),
    .C(_1566_),
    .Y(_1567_)
);

FILL SFILL29000x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4181_),
    .B(_4175_),
    .C(_4162_),
    .Y(_4191_)
);

AOI21X1 _14319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3718_),
    .B(_3717_),
    .C(_3639_),
    .Y(_3732_)
);

AOI21X1 _18992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8853_),
    .B(_8846_),
    .C(_8480_),
    .Y(_8854_)
);

NOR3X1 _18572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7978_),
    .C(_7981_),
    .Y(_8393_)
);

INVX1 _18152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7932_),
    .Y(_7933_)
);

NAND3X1 _20757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10766_),
    .B(_10771_),
    .C(_10778_),
    .Y(_10788_)
);

NOR3X1 _20337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10327_),
    .B(_10325_),
    .C(_10326_),
    .Y(_10328_)
);

FILL SFILL43960x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9706_),
    .B(_9705_),
    .C(_9703_),
    .Y(_9714_)
);

NAND3X1 _19357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9252_),
    .B(_9253_),
    .C(_9251_),
    .Y(_9254_)
);

NAND2X1 _14492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3919_),
    .B(_3921_),
    .Y(_3922_)
);

NAND2X1 _14072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3459_),
    .B(_3461_),
    .Y(_3462_)
);

FILL SFILL43800x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _12805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10452_),
    .B(_253_),
    .Y(_264_)
);

NAND3X1 _22903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1227_),
    .C(_1068_),
    .Y(_1231_)
);

NAND3X1 _15697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5223_),
    .B(_5227_),
    .C(_5230_),
    .Y(_5240_)
);

OAI22X1 _15277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_2465__bF$buf0),
    .C(_7217__bF$buf2),
    .D(_2287__bF$buf0),
    .Y(_4781_)
);

NAND2X1 _20090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf1),
    .B(breg_22_bF$buf1),
    .Y(_10056_)
);

OAI21X1 _21295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11376_),
    .B(_11377_),
    .C(_11372_),
    .Y(_11378_)
);

OAI21X1 _17843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7586_),
    .B(_7587_),
    .C(_7436_),
    .Y(_7594_)
);

NAND3X1 _17423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7130_),
    .B(_7133_),
    .C(_7132_),
    .Y(_7134_)
);

AND2X2 _17003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .B(_6271_),
    .Y(_6673_)
);

FILL SFILL33880x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8450_),
    .B(_8451_),
    .C(_8074_),
    .Y(_8454_)
);

NAND3X1 _18208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7988_),
    .B(_7989_),
    .C(_7987_),
    .Y(_7994_)
);

NOR3X1 _13763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3116_),
    .B(_3119_),
    .C(_3115_),
    .Y(_3123_)
);

INVX2 _13343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2663_),
    .Y(_2664_)
);

NAND2X1 _23861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .B(_2268_),
    .Y(_2271_)
);

XOR2X1 _23441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_1809_),
    .Y(_1817_)
);

INVX1 _23021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1357_),
    .Y(_1359_)
);

OAI21X1 _14968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4436_),
    .B(_4435_),
    .C(_4432_),
    .Y(_4442_)
);

OAI21X1 _14548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_3982_),
    .C(_3948_),
    .Y(_3983_)
);

OAI21X1 _14128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3464_),
    .B(_3462_),
    .C(_3451_),
    .Y(_3522_)
);

FILL SFILL23880x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53960x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8181_),
    .B(_8180_),
    .C(_8182_),
    .Y(_8184_)
);

AOI21X1 _20986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11036_),
    .B(_11037_),
    .C(_11023_),
    .Y(_11038_)
);

NAND3X1 _20566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10574_),
    .B(_10578_),
    .C(_10560_),
    .Y(_10579_)
);

NAND2X1 _20146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf3),
    .B(breg_20_bF$buf1),
    .Y(_10118_)
);

FILL SFILL8840x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_7100__bF$buf2),
    .C(_9492_),
    .Y(_9505_)
);

INVX1 _19166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9043_),
    .Y(_9044_)
);

FILL SFILL13880x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10068_),
    .Y(_10079_)
);

NAND3X1 _22712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1018_),
    .B(_1019_),
    .C(_1021_),
    .Y(_1022_)
);

FILL SFILL29000x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4523_),
    .B(_4524_),
    .C(_4501_),
    .Y(_4572_)
);

FILL SFILL13800x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3164_),
    .B(_3169_),
    .C(_3171_),
    .Y(_3185_)
);

BUFX2 _23917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[35]),
    .Y(y[35])
);

AND2X2 _17652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf2),
    .B(breg_16_bF$buf3),
    .Y(_7384_)
);

INVX2 _17232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6923_),
    .Y(_6924_)
);

FILL SFILL23960x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf4),
    .B(_5921__bF$buf2),
    .C(_8704_),
    .Y(_8705_)
);

OAI22X1 _18437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7440_),
    .B(_8243_),
    .C(_8244_),
    .D(_7882_),
    .Y(_8245_)
);

NOR2X1 _18017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf1),
    .B(_5369_),
    .Y(_7784_)
);

NAND3X1 _13992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3368_),
    .B(_3371_),
    .C(_3373_),
    .Y(_3374_)
);

NOR2X1 _13572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2912_),
    .B(_2914_),
    .Y(_2915_)
);

NOR2X1 _13152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_2454_),
    .Y(_2455_)
);

INVX1 _23670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2010_),
    .Y(_2065_)
);

AOI21X1 _23250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1608_)
);

FILL SFILL64040x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4232_),
    .B(_4229_),
    .Y(_4233_)
);

INVX1 _14357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3770_),
    .Y(_3772_)
);

DFFPOSX1 _24035_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[25]),
    .CLK(clk_bF$buf4),
    .D(a[25])
);

XNOR2X1 _18190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7963_),
    .B(_7958_),
    .Y(_7974_)
);

NAND2X1 _20795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10826_),
    .B(_10823_),
    .Y(_10830_)
);

AOI21X1 _20375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10363_),
    .B(_10368_),
    .C(_10356_),
    .Y(_10369_)
);

OAI21X1 _16923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6579_),
    .B(_6580_),
    .C(_6546_),
    .Y(_6585_)
);

NAND3X1 _16503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6111_),
    .B(_6119_),
    .C(_6114_),
    .Y(_6124_)
);

NOR2X1 _19395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9287_),
    .B(_9288_),
    .Y(_9295_)
);

INVX2 _17708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7444_),
    .Y(_7445_)
);

FILL SFILL18600x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_407_),
    .Y(_691_)
);

AOI21X1 _12423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7821_),
    .B(_7865_),
    .C(_7558_),
    .Y(_7986_)
);

NAND2X1 _22941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1269_),
    .B(_1270_),
    .Y(_1272_)
);

OAI21X1 _12003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3022_),
    .B(_2420_),
    .C(_2978_),
    .Y(_3383_)
);

NAND3X1 _22521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_798_),
    .C(_808_),
    .Y(_813_)
);

NAND3X1 _22101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_350_),
    .C(_351_),
    .Y(_353_)
);

NOR2X1 _13628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2972_),
    .B(_2970_),
    .Y(_2975_)
);

NAND3X1 _13208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2514_),
    .C(_2515_),
    .Y(_2516_)
);

NAND2X1 _23726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2061_),
    .B(_2096_),
    .Y(_2126_)
);

NAND3X1 _23306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1667_),
    .B(_1668_),
    .C(_1561_),
    .Y(_1669_)
);

NAND3X1 _17881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7219_),
    .B(_7631_),
    .C(_7630_),
    .Y(_7636_)
);

NAND3X1 _17461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7156_),
    .B(_7162_),
    .C(_7166_),
    .Y(_7175_)
);

OAI21X1 _17041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6713_),
    .B(_6712_),
    .C(_6709_),
    .Y(_6715_)
);

NAND2X1 _18666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8493_),
    .B(_8494_),
    .Y(_8495_)
);

AOI21X1 _18246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7341_),
    .B(_7603_),
    .C(_8034_),
    .Y(_8035_)
);

OAI21X1 _13381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2622_),
    .B(_2623_),
    .C(_2580_),
    .Y(_2706_)
);

NOR3X1 _14586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4017_),
    .B(_4024_),
    .C(_3779_),
    .Y(_4025_)
);

OAI21X1 _14166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3556_),
    .B(_3557_),
    .C(_3552_),
    .Y(_3564_)
);

FILL SFILL74120x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28840x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10152_),
    .B(_10155_),
    .C(_10159_),
    .Y(_10160_)
);

NAND3X1 _16732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .B(_6362_),
    .C(_6366_),
    .Y(_6376_)
);

NAND2X1 _16312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_22_bF$buf0),
    .Y(_5916_)
);

OAI21X1 _21389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_7100__bF$buf1),
    .C(_11480_),
    .Y(_11481_)
);

AOI21X1 _17937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7695_),
    .B(_7692_),
    .C(_7668_),
    .Y(_7696_)
);

NAND2X1 _17517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_29_bF$buf0),
    .Y(_7235_)
);

OAI21X1 _12652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf2),
    .B(_5420__bF$buf2),
    .C(_10485_),
    .Y(_10496_)
);

NAND3X1 _12232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3953_),
    .B(_5881_),
    .C(_5870_),
    .Y(_5892_)
);

INVX1 _22750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1062_),
    .Y(_1063_)
);

NAND2X1 _22330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_348_),
    .Y(_603_)
);

NAND3X1 _13857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2985_),
    .B(_3212_),
    .C(_3217_),
    .Y(_3227_)
);

XOR2X1 _13437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2765_),
    .Y(_2766_)
);

DFFPOSX1 _23955_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[9]),
    .CLK(clk_bF$buf2),
    .D(_0_[9])
);

OAI21X1 _13017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2305_),
    .C(_2131_),
    .Y(_2312_)
);

OAI21X1 _23535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1918_),
    .B(_1915_),
    .C(_1875_),
    .Y(_1919_)
);

XNOR2X1 _23115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(_1441_),
    .Y(_1461_)
);

NOR3X1 _17690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7053_),
    .B(_7055_),
    .C(_7052_),
    .Y(_7425_)
);

NAND2X1 _17270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6963_),
    .B(_6964_),
    .Y(_6965_)
);

FILL SFILL18680x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38680x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_28_bF$buf5),
    .Y(_8747_)
);

XOR2X1 _18475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8243_),
    .B(_8286_),
    .Y(_8287_)
);

OAI21X1 _18055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_2884__bF$buf3),
    .C(_7825_),
    .Y(_7826_)
);

AOI21X1 _13190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2314_),
    .B(_2313_),
    .C(_2311_),
    .Y(_2496_)
);

INVX4 _11923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf2),
    .Y(_2508_)
);

OAI21X1 _21601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11705_),
    .B(_11704_),
    .C(_11702_),
    .Y(_11713_)
);

OAI21X1 _14395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf2),
    .B(_2362__bF$buf0),
    .C(_3554_),
    .Y(_3815_)
);

DFFPOSX1 _24073_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[31]),
    .CLK(clk_bF$buf3),
    .D(b[31])
);

AOI21X1 _12708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10990_),
    .B(_10946_),
    .C(_10792_),
    .Y(_11110_)
);

XOR2X1 _22806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(_1111_),
    .Y(_1124_)
);

FILL SFILL8520x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6624_),
    .B(_6625_),
    .C(_6611_),
    .Y(_6627_)
);

NAND2X1 _16541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_17_bF$buf3),
    .Y(_6166_)
);

OAI21X1 _16121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5400_),
    .B(_5402_),
    .C(_5393_),
    .Y(_5706_)
);

NAND3X1 _21198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11254_),
    .B(_11258_),
    .C(_11271_),
    .Y(_11272_)
);

AOI21X1 _17746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6655_),
    .B(_7486_),
    .C(_7080_),
    .Y(_7487_)
);

INVX2 _17326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7025_),
    .Y(_7026_)
);

NAND3X1 _12881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_1086_),
    .C(_11657_),
    .Y(_1096_)
);

NOR3X1 _12461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5947_),
    .B(_8359_),
    .C(_7164_),
    .Y(_8402_)
);

NAND3X1 _12041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3547_),
    .B(_3734_),
    .C(_3745_),
    .Y(_3799_)
);

FILL SFILL38760x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3008_),
    .B(_3007_),
    .C(_3004_),
    .Y(_3017_)
);

INVX1 _13246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .Y(_2557_)
);

NAND2X1 _23764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2130_),
    .B(_2146_),
    .Y(_2167_)
);

XNOR2X1 _23344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .B(_1710_),
    .Y(_1711_)
);

FILL SFILL64120x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5252_),
    .B(_5254_),
    .C(_5242_),
    .Y(_5367_)
);

AOI21X1 _18284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8022_),
    .B(_8023_),
    .C(_7782_),
    .Y(_8077_)
);

FILL SFILL28760x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL9000x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _20889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10911_),
    .Y(_10933_)
);

OAI21X1 _20469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253__bF$buf2),
    .B(_3958__bF$buf2),
    .C(_10471_),
    .Y(_10472_)
);

NAND2X1 _20049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10009_),
    .B(_10010_),
    .Y(_10011_)
);

OAI21X1 _21830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11726_),
    .B(_54_),
    .C(_11748_),
    .Y(_55_)
);

NAND3X1 _21410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11475_),
    .B(_11489_),
    .C(_11495_),
    .Y(_11504_)
);

XNOR2X1 _19489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9397_),
    .B(_9393_),
    .Y(_9398_)
);

NAND2X1 _19069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_26_bF$buf2),
    .Y(_8937_)
);

FILL SFILL54120x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1565_),
    .B(_1663_),
    .Y(_1707_)
);

NOR2X1 _12517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8994_),
    .B(_9005_),
    .Y(_9016_)
);

NAND3X1 _22615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_715_),
    .B(_915_),
    .C(_722_),
    .Y(_916_)
);

XOR2X1 _16770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6042_),
    .B(_6416_),
    .Y(_0_[28])
);

AOI21X1 _16350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5952_),
    .B(_5951_),
    .C(_5950_),
    .Y(_5957_)
);

FILL SFILL18680x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert340 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf1)
);

BUFX2 BUFX2_insert341 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf0)
);

BUFX2 BUFX2_insert342 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf5)
);

BUFX2 BUFX2_insert343 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf4)
);

NAND3X1 _17975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7730_),
    .B(_7735_),
    .C(_7737_),
    .Y(_7738_)
);

BUFX2 BUFX2_insert344 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf3)
);

BUFX2 BUFX2_insert345 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf2)
);

AOI22X1 _17555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_25_bF$buf3),
    .C(areg_7_bF$buf3),
    .D(breg_24_bF$buf4),
    .Y(_7277_)
);

INVX2 _17135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6816_),
    .Y(_6817_)
);

BUFX2 BUFX2_insert346 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf1)
);

BUFX2 BUFX2_insert347 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(breg_3_bF$buf0)
);

BUFX2 BUFX2_insert348 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104_),
    .Y(_9104__bF$buf3)
);

NOR2X1 _12690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9137_),
    .B(_10902_),
    .Y(_10913_)
);

BUFX2 BUFX2_insert349 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104_),
    .Y(_9104__bF$buf2)
);

NAND2X1 _12270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6264_),
    .B(_6176_),
    .Y(_6308_)
);

OAI21X1 _13895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2993_),
    .B(_3266_),
    .C(_3267_),
    .Y(_3268_)
);

OAI21X1 _13475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf1),
    .B(_6044__bF$buf2),
    .C(_2596_),
    .Y(_2808_)
);

DFFPOSX1 _23993_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[47]),
    .CLK(clk_bF$buf8),
    .D(_0_[47])
);

NAND2X1 _23573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2969_),
    .B(_1959_),
    .Y(_1960_)
);

AOI21X1 _13055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2342_),
    .B(_2343_),
    .C(_1096_),
    .Y(_2350_)
);

XOR2X1 _23153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1502_),
    .Y(_1503_)
);

XNOR2X1 _19701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9265_),
    .B(_9630_),
    .Y(_0_[36])
);

NAND2X1 _15621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5155_),
    .B(_5156_),
    .Y(_5158_)
);

NAND3X1 _15201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4693_),
    .B(_4696_),
    .C(_4685_),
    .Y(_4698_)
);

NAND3X1 _18093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7863_),
    .B(_7862_),
    .C(_7861_),
    .Y(_7868_)
);

AOI21X1 _20698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10711_),
    .B(_10710_),
    .C(_10707_),
    .Y(_10723_)
);

INVX2 _20278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10262_),
    .Y(_10263_)
);

OAI21X1 _16826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6136_),
    .B(_6477_),
    .C(_6158_),
    .Y(_6478_)
);

NOR3X1 _16406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6013_),
    .B(_6014_),
    .C(_6011_),
    .Y(_6018_)
);

NOR2X1 _11961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2781_),
    .B(_2913_),
    .Y(_2924_)
);

FILL SFILL69240x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9139_),
    .B(_9138_),
    .C(_9097_),
    .Y(_9189_)
);

NAND3X1 _12746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9641_),
    .B(_11516_),
    .C(_11505_),
    .Y(_11527_)
);

NOR3X1 _12326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6889_),
    .B(_6878_),
    .C(_6845_),
    .Y(_6922_)
);

NAND3X1 _22844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1160_),
    .B(_1133_),
    .C(_1165_),
    .Y(_1166_)
);

NAND3X1 _22424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .B(_706_),
    .C(_704_),
    .Y(_707_)
);

OAI21X1 _22004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_11886_),
    .C(_215_),
    .Y(_246_)
);

FILL SFILL3800x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2019_),
    .B(_2020_),
    .C(_2006_),
    .Y(_2021_)
);

NAND2X1 _23209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf3),
    .B(breg_27_bF$buf0),
    .Y(_1563_)
);

NAND2X1 _17784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf4),
    .B(areg_29_bF$buf4),
    .Y(_7529_)
);

AND2X2 _17364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_23_bF$buf2),
    .Y(_7069_)
);

FILL SFILL59160x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10955_),
    .Y(_10956_)
);

NAND3X1 _18989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8843_),
    .B(_8844_),
    .C(_8842_),
    .Y(_8849_)
);

NAND2X1 _18569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8379_),
    .B(_8381_),
    .Y(_8389_)
);

INVX1 _18149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7490_),
    .Y(_7929_)
);

OAI21X1 _13284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .B(_2596_),
    .C(_2597_),
    .Y(_2598_)
);

OAI21X1 _23382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1752_),
    .B(_1747_),
    .C(_1662_),
    .Y(_1753_)
);

OAI21X1 _19930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9880_),
    .B(_9881_),
    .C(_9877_),
    .Y(_9882_)
);

AOI21X1 _19510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9407_),
    .B(_9412_),
    .C(_9399_),
    .Y(_9421_)
);

FILL SFILL33960x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf1),
    .B(_549__bF$buf3),
    .Y(_3918_)
);

NAND3X1 _14069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3457_),
    .B(_3309_),
    .C(_3451_),
    .Y(_3458_)
);

NAND2X1 _15850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_17_bF$buf4),
    .Y(_5408_)
);

NOR3X1 _15430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4622_),
    .B(_4623_),
    .C(_4620_),
    .Y(_4949_)
);

NOR3X1 _15010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4486_),
    .B(_4487_),
    .C(_4485_),
    .Y(_4488_)
);

OR2X2 _20087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10047_),
    .B(_10048_),
    .Y(_10053_)
);

AND2X2 _16635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_21_bF$buf2),
    .Y(_6269_)
);

OAI21X1 _16215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5807_),
    .B(_5808_),
    .C(_5806_),
    .Y(_5809_)
);

FILL SFILL23960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2088_),
    .B(_2109_),
    .C(_2099_),
    .Y(_2120_)
);

AOI21X1 _12555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7920_),
    .B(_7547_),
    .C(_7975_),
    .Y(_9433_)
);

OAI21X1 _12135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4807_),
    .B(_4818_),
    .C(_3449_),
    .Y(_4829_)
);

NOR2X1 _22653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf2),
    .B(_6815__bF$buf4),
    .Y(_957_)
);

OAI21X1 _22233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_248_),
    .C(_461_),
    .Y(_497_)
);

NOR2X1 _23858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .B(_2248_),
    .Y(_2267_)
);

OAI21X1 _23438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5318_),
    .B(_9153_),
    .C(_1812_),
    .Y(_1813_)
);

NOR2X1 _23018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(_1353_),
    .Y(_1355_)
);

OAI21X1 _14701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4143_),
    .B(_4142_),
    .C(_4140_),
    .Y(_4150_)
);

AOI21X1 _17593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7308_),
    .B(_7302_),
    .C(_7274_),
    .Y(_7319_)
);

NAND3X1 _17173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6852_),
    .B(_6858_),
    .C(_6855_),
    .Y(_6859_)
);

OAI21X1 _15906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5106_),
    .B(_5468_),
    .C(_5469_),
    .Y(_5470_)
);

INVX1 _18798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8639_),
    .Y(_8640_)
);

AND2X2 _18378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7760_),
    .B(_7750_),
    .Y(_8180_)
);

AOI21X1 _13093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1586_),
    .B(_1609_),
    .C(_2389_),
    .Y(_2390_)
);

AOI21X1 _23191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .B(_1531_),
    .C(_1542_),
    .Y(_1544_)
);

FILL SFILL59240x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_157_),
    .B(_158_),
    .C(_156_),
    .Y(_159_)
);

OAI21X1 _21504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11345_),
    .B(_11332_),
    .C(_11355_),
    .Y(_11607_)
);

OAI21X1 _14298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3663_),
    .B(_3664_),
    .C(_3641_),
    .Y(_3709_)
);

FILL SFILL3800x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3800x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_978_),
    .B(_974_),
    .Y(_1018_)
);

FILL FILL74200x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _16864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6519_),
    .Y(_6520_)
);

OAI21X1 _16444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5686_),
    .B(_5691_),
    .C(_5680_),
    .Y(_6059_)
);

NAND3X1 _16024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5465_),
    .B(_5509_),
    .C(_5507_),
    .Y(_5600_)
);

OAI21X1 _17649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6972_),
    .B(_6961_),
    .C(_6965_),
    .Y(_7380_)
);

AOI21X1 _17229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6742_),
    .B(_6749_),
    .C(_6602_),
    .Y(_6920_)
);

NAND3X1 _12784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_23_),
    .B(_11866_),
    .C(_1_),
    .Y(_34_)
);

NAND2X1 _12364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_7_bF$buf1),
    .Y(_7338_)
);

NAND3X1 _22882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1203_),
    .B(_1207_),
    .C(_1205_),
    .Y(_1208_)
);

XOR2X1 _22462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .B(_747_),
    .Y(_748_)
);

NOR3X1 _22042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_284_),
    .B(_285_),
    .C(_287_),
    .Y(_288_)
);

OAI21X1 _13989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf1),
    .B(_549__bF$buf4),
    .C(_3364_),
    .Y(_3370_)
);

OAI21X1 _13569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2860_),
    .B(_2859_),
    .C(_2855_),
    .Y(_2911_)
);

NAND2X1 _13149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_12_bF$buf1),
    .Y(_2451_)
);

NAND2X1 _23667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2042_),
    .B(_2026_),
    .Y(_2062_)
);

NAND3X1 _23247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_1601_),
    .C(_1604_),
    .Y(_1605_)
);

FILL SFILL18760x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_15_bF$buf5),
    .Y(_4400_)
);

INVX2 _14510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .Y(_3941_)
);

FILL SFILL34040x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5259_),
    .B(_5260_),
    .C(_5252_),
    .Y(_5261_)
);

AND2X2 _18187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7966_),
    .B(_7970_),
    .Y(_7971_)
);

FILL SFILL23960x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11856_),
    .B(_11857_),
    .C(_11597_),
    .Y(_11858_)
);

NAND3X1 _21313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11396_),
    .B(_11394_),
    .C(_11397_),
    .Y(_11398_)
);

FILL SFILL69320x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1174_),
    .Y(_1268_)
);

OAI21X1 _22518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_805_),
    .B(_806_),
    .C(_808_),
    .Y(_809_)
);

AND2X2 _16673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf1),
    .B(areg_27_bF$buf4),
    .Y(_6311_)
);

NAND2X1 _16253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .B(_5850_),
    .Y(_5851_)
);

NAND3X1 _17878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6843_),
    .B(_7631_),
    .C(_7630_),
    .Y(_7632_)
);

NAND3X1 _17458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6924_),
    .B(_7010_),
    .C(_7011_),
    .Y(_7172_)
);

NAND2X1 _17038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6705_),
    .B(_6697_),
    .Y(_6711_)
);

NAND3X1 _12593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9784_),
    .B(_9707_),
    .C(_9751_),
    .Y(_9850_)
);

FILL SFILL59320x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5135_),
    .Y(_5245_)
);

XNOR2X1 _22691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_982_),
    .Y(_999_)
);

NAND3X1 _22271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_537_),
    .C(_536_),
    .Y(_539_)
);

OAI21X1 _13798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3161_),
    .B(_3160_),
    .C(_3141_),
    .Y(_3162_)
);

OAI21X1 _13378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_2700_),
    .C(_2699_),
    .Y(_2702_)
);

BUFX2 _23896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[14]),
    .Y(y[14])
);

NAND3X1 _23476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .B(_1850_),
    .C(_1854_),
    .Y(_1855_)
);

NAND2X1 _23056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1396_),
    .B(_1392_),
    .Y(_1397_)
);

NAND3X1 _19604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9520_),
    .B(_9509_),
    .C(_9515_),
    .Y(_9525_)
);

FILL FILL74200x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5216_),
    .B(_5211_),
    .C(_5181_),
    .Y(_5512_)
);

NAND3X1 _15524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5045_),
    .B(_5050_),
    .C(_5049_),
    .Y(_5051_)
);

NAND3X1 _15104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4584_),
    .B(_4591_),
    .C(_4447_),
    .Y(_4592_)
);

OAI21X1 _16729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6211_),
    .B(_6206_),
    .C(_6213_),
    .Y(_6372_)
);

NAND2X1 _16309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5907_),
    .B(_5911_),
    .Y(_5912_)
);

AOI21X1 _21962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_86_),
    .C(_88_),
    .Y(_201_)
);

NAND2X1 _21542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11387_),
    .B(_11393_),
    .Y(_11648_)
);

OAI21X1 _21122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf2),
    .B(_7520__bF$buf3),
    .C(_10865_),
    .Y(_11189_)
);

FILL SFILL13880x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_6_bF$buf3),
    .Y(_10463_)
);

NAND3X1 _12229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4970_),
    .B(_5804_),
    .C(_5848_),
    .Y(_5859_)
);

INVX2 _22747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1059_),
    .Y(_1060_)
);

AOI21X1 _22327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_591_),
    .C(_540_),
    .Y(_600_)
);

OAI21X1 _16482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6098_),
    .B(_6100_),
    .C(_6097_),
    .Y(_6101_)
);

NAND3X1 _16062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5306_),
    .B(_5641_),
    .C(_5634_),
    .Y(_5642_)
);

NAND3X1 _17687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7414_),
    .B(_7421_),
    .C(_7419_),
    .Y(_7422_)
);

INVX1 _17267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6961_),
    .Y(_6962_)
);

FILL SFILL23640x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_318_),
    .C(_298_),
    .Y(_329_)
);

OAI21X1 _20813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10525_),
    .B(_10523_),
    .C(_10514_),
    .Y(_10850_)
);

FILL SFILL13640x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2448_),
    .B(_2474_),
    .C(_2479_),
    .Y(_2493_)
);

NAND3X1 _23285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1643_),
    .C(_1641_),
    .Y(_1647_)
);

NOR2X1 _19833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9768_),
    .B(_9769_),
    .Y(_9776_)
);

NAND3X1 _19413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9281_),
    .B(_9306_),
    .C(_9303_),
    .Y(_9315_)
);

AOI21X1 _15753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5301_),
    .B(_4648_),
    .C(_5300_),
    .Y(_5302_)
);

AOI21X1 _15333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4824_),
    .B(_4828_),
    .C(_4833_),
    .Y(_4843_)
);

FILL SFILL74200x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6228_),
    .B(_6232_),
    .C(_6235_),
    .Y(_6623_)
);

OAI21X1 _16538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5808_),
    .B(_5806_),
    .C(_5798_),
    .Y(_6162_)
);

NAND3X1 _16118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5684_),
    .B(_5698_),
    .C(_5687_),
    .Y(_5702_)
);

AND2X2 _21771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_28_bF$buf1),
    .Y(_11899_)
);

AND2X2 _21351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11205_),
    .B(_11197_),
    .Y(_11440_)
);

FILL SFILL64280x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1009_),
    .B(_1020_),
    .C(_11679_),
    .Y(_1064_)
);

OAI21X1 _12458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7164_),
    .B(_5947_),
    .C(_7109_),
    .Y(_8370_)
);

OAI21X1 _22976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1038_),
    .B(_1192_),
    .C(_1198_),
    .Y(_1309_)
);

OAI21X1 _12038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3723_),
    .B(_3756_),
    .C(_3493_),
    .Y(_3776_)
);

NAND2X1 _22556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf4),
    .B(areg_27_bF$buf5),
    .Y(_851_)
);

AOI21X1 _22136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_391_)
);

AND2X2 _16291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .B(areg_21_bF$buf2),
    .Y(_5893_)
);

AOI21X1 _14604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4042_),
    .B(_4043_),
    .C(_3763_),
    .Y(_4044_)
);

AND2X2 _17496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7209_),
    .B(_7212_),
    .Y(_7213_)
);

AOI21X1 _17076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6748_),
    .B(_6746_),
    .C(_6745_),
    .Y(_6753_)
);

NOR2X1 _15809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5355_),
    .B(_5353_),
    .Y(_5363_)
);

OAI21X1 _20622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10636_),
    .B(_10640_),
    .C(_10344_),
    .Y(_10641_)
);

OAI21X1 _20202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10177_),
    .B(_10179_),
    .C(_10174_),
    .Y(_10180_)
);

NAND3X1 _23094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1303_),
    .B(_1307_),
    .C(_1309_),
    .Y(_1438_)
);

NAND3X1 _19642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9564_),
    .B(_9566_),
    .C(_9563_),
    .Y(_9567_)
);

NAND2X1 _19222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf2),
    .B(areg_24_bF$buf1),
    .Y(_9106_)
);

OAI21X1 _21827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_44_),
    .C(_41_),
    .Y(_52_)
);

OAI21X1 _21407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11496_),
    .B(_11500_),
    .C(_11473_),
    .Y(_11501_)
);

AND2X2 _15982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5549_),
    .B(_5553_),
    .Y(_5554_)
);

AOI21X1 _15562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5072_),
    .B(_5078_),
    .C(_5040_),
    .Y(_5093_)
);

AOI21X1 _15142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4618_),
    .B(_4624_),
    .C(_4350_),
    .Y(_4634_)
);

FILL SFILL8680x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6405_),
    .B(_6399_),
    .C(_6403_),
    .Y(_6414_)
);

NAND3X1 _16347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5915_),
    .B(_5953_),
    .C(_5949_),
    .Y(_5954_)
);

NAND3X1 _21580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11687_),
    .B(_11688_),
    .C(_11686_),
    .Y(_11689_)
);

NAND2X1 _21160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_29_bF$buf2),
    .Y(_11230_)
);

FILL SFILL8600x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53800x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_10869__bF$buf3),
    .C(_9137_),
    .Y(_10880_)
);

OAI21X1 _12267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6253_),
    .B(_6242_),
    .C(_6264_),
    .Y(_6275_)
);

OAI21X1 _22785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1077_),
    .B(_1076_),
    .C(_1073_),
    .Y(_1101_)
);

OR2X2 _22365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_406_),
    .Y(_642_)
);

NOR3X1 _18913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8758_),
    .B(_8761_),
    .C(_8757_),
    .Y(_8767_)
);

FILL SFILL74280x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4287_),
    .B(_4294_),
    .C(_4154_),
    .Y(_4295_)
);

NOR3X1 _14413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3830_),
    .B(_3823_),
    .C(_3829_),
    .Y(_3835_)
);

FILL SFILL74200x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5153_),
    .Y(_5154_)
);

FILL SFILL3480x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10887_),
    .B(_10886_),
    .C(_10850_),
    .Y(_10892_)
);

INVX2 _20431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10393_),
    .Y(_10431_)
);

AOI21X1 _20011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9965_),
    .B(_9969_),
    .C(_9638_),
    .Y(_9971_)
);

OAI21X1 _19871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9432_),
    .B(_9816_),
    .C(_9435_),
    .Y(_9818_)
);

NOR3X1 _19451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9351_),
    .B(_9350_),
    .C(_9352_),
    .Y(_9357_)
);

NOR2X1 _19031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf4),
    .B(_6815__bF$buf1),
    .Y(_8896_)
);

INVX1 _11958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2749_),
    .Y(_2901_)
);

NOR2X1 _21636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11746_),
    .B(_11750_),
    .Y(_11751_)
);

AOI21X1 _21216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10981_),
    .B(_10694_),
    .C(_11291_),
    .Y(_11292_)
);

FILL SFILL28840x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5342_),
    .B(_5338_),
    .C(_4979_),
    .Y(_5344_)
);

NAND3X1 _15371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4878_),
    .B(_4883_),
    .C(_4845_),
    .Y(_4885_)
);

OAI21X1 _16996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6304_),
    .B(_6294_),
    .C(_6299_),
    .Y(_6665_)
);

NAND3X1 _16576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6202_),
    .B(_6203_),
    .C(_6201_),
    .Y(_6204_)
);

AOI21X1 _16156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5599_),
    .B(_5605_),
    .C(_5463_),
    .Y(_5744_)
);

OAI21X1 _12496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8764_),
    .B(_8775_),
    .C(_8742_),
    .Y(_8786_)
);

OAI21X1 _12076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .B(_4160_),
    .C(_4171_),
    .Y(_4182_)
);

INVX1 _22594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .Y(_893_)
);

NAND3X1 _22174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_432_),
    .C(_366_),
    .Y(_433_)
);

NAND3X1 _18722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8553_),
    .B(_8554_),
    .C(_8556_),
    .Y(_8557_)
);

NOR2X1 _18302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8089_),
    .B(_8090_),
    .Y(_8097_)
);

FILL SFILL23720x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10906_),
    .B(_10907_),
    .C(_10905_),
    .Y(_10953_)
);

NAND2X1 _23799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2159_),
    .B(_2119_),
    .Y(_2205_)
);

AOI22X1 _23379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1748_),
    .B(_1621_),
    .C(_1744_),
    .D(_1745_),
    .Y(_1749_)
);

OAI21X1 _19927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_7520__bF$buf2),
    .C(_9865_),
    .Y(_9879_)
);

NAND3X1 _19507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9413_),
    .B(_9417_),
    .C(_9398_),
    .Y(_9418_)
);

OAI21X1 _14642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_3529__bF$buf0),
    .C(_4078_),
    .Y(_4085_)
);

AOI21X1 _14222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3378_),
    .B(_3360_),
    .C(_3381_),
    .Y(_3626_)
);

FILL SFILL48920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5070_),
    .B(_5067_),
    .C(_5059_),
    .Y(_5405_)
);

AOI21X1 _15427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4932_),
    .B(_4936_),
    .C(_4656_),
    .Y(_4946_)
);

AOI21X1 _15007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4480_),
    .B(_4481_),
    .C(_4479_),
    .Y(_4485_)
);

NOR2X1 _20660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10680_),
    .B(_10679_),
    .Y(_10681_)
);

NAND2X1 _20240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10218_),
    .B(_10219_),
    .Y(_10220_)
);

AOI21X1 _19680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9606_),
    .B(_9607_),
    .C(_9273_),
    .Y(_9608_)
);

NAND2X1 _19260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9142_),
    .B(_9146_),
    .Y(_9147_)
);

AND2X2 _21865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11794_),
    .B(_11785_),
    .Y(_94_)
);

INVX1 _21445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11522_),
    .Y(_11543_)
);

OAI21X1 _21025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11078_),
    .B(_11076_),
    .C(_11081_),
    .Y(_11082_)
);

AOI21X1 _15180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4584_),
    .B(_4591_),
    .C(_4447_),
    .Y(_4674_)
);

NOR3X1 _13913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3281_),
    .B(_3283_),
    .C(_3282_),
    .Y(_3288_)
);

FILL SFILL38840x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5993_),
    .B(_5992_),
    .C(_5994_),
    .Y(_5995_)
);

FILL SFILL69240x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8806_),
    .B(_8807_),
    .C(_8766_),
    .Y(_8809_)
);

NAND3X1 _18531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8347_),
    .B(_8342_),
    .C(_8345_),
    .Y(_8349_)
);

OAI21X1 _18111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7454_),
    .B(_7444_),
    .C(_7449_),
    .Y(_7888_)
);

FILL SFILL3880x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10400_),
    .B(_10395_),
    .C(_10403_),
    .Y(_10743_)
);

FILL SFILL28840x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24120x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _23188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1531_),
    .B(_1536_),
    .C(_1397_),
    .Y(_1540_)
);

AOI21X1 _19736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9667_),
    .B(_9668_),
    .C(_9653_),
    .Y(_9669_)
);

NAND3X1 _19316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9202_),
    .B(_9096_),
    .C(_9199_),
    .Y(_9209_)
);

NOR3X1 _14871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3749_),
    .B(_3752_),
    .C(_3755_),
    .Y(_4337_)
);

AND2X2 _14451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_12_bF$buf0),
    .Y(_3877_)
);

AOI21X1 _14031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3404_),
    .B(_3401_),
    .C(_3398_),
    .Y(_3417_)
);

INVX2 _15656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5195_),
    .Y(_5196_)
);

NOR3X1 _15236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4728_),
    .B(_4732_),
    .C(_4727_),
    .Y(_4736_)
);

FILL SFILL54200x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _11996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3209_),
    .B(_3187_),
    .Y(_3307_)
);

OAI21X1 _21674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11791_),
    .B(_11792_),
    .C(_11787_),
    .Y(_11793_)
);

OAI21X1 _21254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11032_),
    .B(_11023_),
    .C(_11027_),
    .Y(_11333_)
);

OAI21X1 _17802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7544_),
    .B(_7543_),
    .C(_7528_),
    .Y(_7549_)
);

FILL SFILL38840x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_31_bF$buf2),
    .Y(_1204_)
);

OAI21X1 _22459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf2),
    .B(_6427_),
    .C(_743_),
    .Y(_744_)
);

AOI21X1 _22039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11893_),
    .B(_10_),
    .C(_8_),
    .Y(_284_)
);

INVX1 _13722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3058_),
    .Y(_3079_)
);

OAI21X1 _13302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2613_),
    .B(_2614_),
    .C(_2618_),
    .Y(_2619_)
);

INVX1 _23820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .Y(_2227_)
);

NOR2X1 _23400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(_1655_),
    .Y(_1771_)
);

AND2X2 _16194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_16_bF$buf4),
    .Y(_5785_)
);

NAND2X1 _14927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_16_bF$buf2),
    .Y(_4397_)
);

AOI22X1 _14507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3671_),
    .B(_3673_),
    .C(_3937_),
    .D(_3670_),
    .Y(_3938_)
);

OAI21X1 _17399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6695_),
    .B(_6700_),
    .C(_6699_),
    .Y(_7107_)
);

NAND2X1 _18760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8593_),
    .B(_8597_),
    .Y(_8598_)
);

INVX1 _18340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8137_),
    .Y(_8138_)
);

NAND3X1 _20945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10690_),
    .B(_10989_),
    .C(_10991_),
    .Y(_10995_)
);

OAI21X1 _20525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10532_),
    .B(_10533_),
    .C(_10528_),
    .Y(_10534_)
);

AOI21X1 _20105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10067_),
    .B(_10069_),
    .C(_10066_),
    .Y(_10073_)
);

NAND2X1 _19965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9912_),
    .B(_9555_),
    .Y(_9920_)
);

AOI21X1 _19545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9435_),
    .B(_9438_),
    .C(_9448_),
    .Y(_9460_)
);

NAND3X1 _19125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8989_),
    .B(_8995_),
    .C(_8985_),
    .Y(_8999_)
);

NAND3X1 _14680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4098_),
    .B(_4121_),
    .C(_4125_),
    .Y(_4126_)
);

AOI21X1 _14260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3406_),
    .B(_3410_),
    .C(_3396_),
    .Y(_3667_)
);

NAND3X1 _15885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5437_),
    .B(_5430_),
    .C(_5435_),
    .Y(_5447_)
);

NOR2X1 _15465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4982_),
    .B(_4984_),
    .Y(_4986_)
);

AOI21X1 _15045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4252_),
    .B(_4249_),
    .C(_4242_),
    .Y(_4527_)
);

FILL SFILL48680x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3560x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11285_),
    .B(_11289_),
    .C(_11292_),
    .Y(_11585_)
);

OAI21X1 _21063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11120_),
    .B(_11119_),
    .C(_11123_),
    .Y(_11124_)
);

FILL SFILL28920x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7331_),
    .B(_7330_),
    .C(_7328_),
    .Y(_7339_)
);

XOR2X1 _22688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_994_),
    .B(_982_),
    .Y(_995_)
);

OAI21X1 _22268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_534_),
    .B(_530_),
    .C(_503_),
    .Y(_535_)
);

OAI21X1 _18816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8655_),
    .B(_8656_),
    .C(_8659_),
    .Y(_8660_)
);

NAND3X1 _13951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3324_),
    .B(_3328_),
    .C(_3327_),
    .Y(_3330_)
);

OAI21X1 _13531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2682_),
    .B(_2680_),
    .C(_2675_),
    .Y(_2870_)
);

NAND3X1 _13111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2402_),
    .B(_2406_),
    .C(_2408_),
    .Y(_2409_)
);

FILL SFILL18920x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3941_),
    .B(_3944_),
    .C(_3934_),
    .Y(_4188_)
);

OAI21X1 _14316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3448_),
    .B(_3446_),
    .C(_3435_),
    .Y(_3729_)
);

FILL SFILL18680x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10783_),
    .B(_10784_),
    .C(_10782_),
    .Y(_10785_)
);

OAI21X1 _20334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10324_),
    .B(_9638_),
    .C(_9972_),
    .Y(_10325_)
);

NAND3X1 _19774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9690_),
    .B(_9710_),
    .C(_9704_),
    .Y(_9711_)
);

AOI21X1 _19354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8474_),
    .B(_8867_),
    .C(_9250_),
    .Y(_9251_)
);

OAI21X1 _21959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_196_),
    .C(_11888_),
    .Y(_197_)
);

NAND3X1 _21539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11605_),
    .B(_11644_),
    .C(_11643_),
    .Y(_11645_)
);

AOI21X1 _21119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11178_),
    .B(_11179_),
    .C(_11170_),
    .Y(_11185_)
);

OAI22X1 _12802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8983_),
    .B(_221_),
    .C(_10726_),
    .D(_10770_),
    .Y(_232_)
);

OAI21X1 _22900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .B(_1222_),
    .C(_1219_),
    .Y(_1227_)
);

OAI21X1 _15694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5141_),
    .B(_5137_),
    .C(_5143_),
    .Y(_5237_)
);

AND2X2 _15274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_14_bF$buf0),
    .Y(_4778_)
);

FILL SFILL69080x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf0),
    .B(_2362__bF$buf3),
    .C(_6552_),
    .Y(_6558_)
);

AND2X2 _16479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5690_),
    .Y(_6097_)
);

AOI21X1 _16059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5637_),
    .B(_5636_),
    .C(_5630_),
    .Y(_5638_)
);

NAND2X1 _21292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf2),
    .B(breg_24_bF$buf0),
    .Y(_11375_)
);

FILL SFILL38600x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7430_),
    .B(_7422_),
    .C(_7428_),
    .Y(_7590_)
);

NAND2X1 _17420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7105_),
    .B(_7102_),
    .Y(_7130_)
);

AOI21X1 _17000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6295_),
    .B(_6301_),
    .C(_6303_),
    .Y(_6669_)
);

OAI21X1 _12399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf0),
    .B(_7711__bF$buf1),
    .C(_6571_),
    .Y(_7722_)
);

AND2X2 _22497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_610_),
    .B(_611_),
    .Y(_786_)
);

OAI21X1 _22077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_325_),
    .C(_123_),
    .Y(_326_)
);

NAND3X1 _18625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8076_),
    .B(_8437_),
    .C(_8442_),
    .Y(_8451_)
);

OAI21X1 _18205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7985_),
    .B(_7990_),
    .C(_7928_),
    .Y(_7991_)
);

FILL SFILL59080x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3115_),
    .B(_3116_),
    .C(_3119_),
    .Y(_3120_)
);

AOI21X1 _13340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2460_),
    .B(_2466_),
    .C(_2462_),
    .Y(_2660_)
);

FILL SFILL59000x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .B(_4433_),
    .C(_4438_),
    .Y(_4439_)
);

NAND3X1 _14545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3956_),
    .B(_3971_),
    .C(_3976_),
    .Y(_3980_)
);

OAI21X1 _14125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3518_),
    .B(_3476_),
    .C(_3466_),
    .Y(_3519_)
);

FILL SFILL3560x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10707_),
    .B(_10711_),
    .C(_10714_),
    .Y(_11035_)
);

NOR3X1 _20563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10563_),
    .B(_10567_),
    .C(_10571_),
    .Y(_10576_)
);

XOR2X1 _20143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10056_),
    .B(_10114_),
    .Y(_10115_)
);

FILL SFILL28920x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9496_),
    .B(_9489_),
    .C(_9501_),
    .Y(_9502_)
);

AND2X2 _19163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_19_bF$buf4),
    .Y(_9041_)
);

FILL SFILL49000x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11622_),
    .B(_11611_),
    .C(_11616_),
    .Y(_11895_)
);

OAI21X1 _21348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11429_),
    .B(_11427_),
    .C(_11425_),
    .Y(_11436_)
);

NAND2X1 _12611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_9_bF$buf2),
    .Y(_10046_)
);

OAI21X1 _15083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4567_),
    .B(_4568_),
    .C(_4565_),
    .Y(_4569_)
);

FILL SFILL39080x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3178_),
    .B(_3181_),
    .C(_3096_),
    .Y(_3182_)
);

BUFX2 _23914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[32]),
    .Y(y[32])
);

NAND2X1 _16288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_19_bF$buf3),
    .Y(_5889_)
);

FILL SFILL63960x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL4040x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8307_),
    .B(_8290_),
    .C(_8298_),
    .Y(_8702_)
);

AOI21X1 _18434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8231_),
    .B(_8230_),
    .C(_8228_),
    .Y(_8242_)
);

AOI21X1 _18014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7582_),
    .B(_7573_),
    .C(_7436_),
    .Y(_7781_)
);

NAND3X1 _20619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10633_),
    .B(_10634_),
    .C(_10348_),
    .Y(_10637_)
);

NOR3X1 _19639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9166_),
    .B(_9175_),
    .C(_9172_),
    .Y(_9563_)
);

XOR2X1 _19219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9059_),
    .B(_9100_),
    .Y(_9101_)
);

NOR3X1 _14774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4224_),
    .B(_4227_),
    .C(_4223_),
    .Y(_4230_)
);

NAND2X1 _14354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3766_),
    .B(_3769_),
    .Y(_3770_)
);

DFFPOSX1 _24032_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[22]),
    .CLK(clk_bF$buf8),
    .D(a[22])
);

NOR2X1 _15979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .B(_5546_),
    .Y(_5550_)
);

OAI21X1 _15559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4801_),
    .B(_4808_),
    .C(_4810_),
    .Y(_5089_)
);

NOR3X1 _15139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4630_)
);

OAI21X1 _20792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf3),
    .B(_4551__bF$buf0),
    .C(_10826_),
    .Y(_10827_)
);

NOR2X1 _20372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10015_),
    .B(_10365_),
    .Y(_10366_)
);

FILL SFILL74360x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6579_),
    .B(_6580_),
    .C(_6578_),
    .Y(_6581_)
);

OAI21X1 _16500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6117_),
    .B(_6118_),
    .C(_6119_),
    .Y(_6120_)
);

NAND3X1 _19392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9286_),
    .B(_9291_),
    .C(_9289_),
    .Y(_9292_)
);

INVX1 _21997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .Y(_238_)
);

INVX2 _21577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11648_),
    .Y(_11686_)
);

INVX2 _21157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11226_),
    .Y(_11227_)
);

XNOR2X1 _17705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7441_),
    .B(_7439_),
    .Y(_7442_)
);

AOI21X1 _12840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_538_),
    .C(_505_),
    .Y(_648_)
);

NAND3X1 _12420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7316_),
    .B(_7514_),
    .C(_7525_),
    .Y(_7953_)
);

NOR2X1 _12000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3044_),
    .B(_3318_),
    .Y(_3350_)
);

FILL SFILL3640x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2970_),
    .B(_2972_),
    .C(_2740_),
    .Y(_2973_)
);

NAND3X1 _13205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2374_),
    .B(_2506_),
    .C(_2512_),
    .Y(_2513_)
);

INVX1 _23723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2081_),
    .Y(_2123_)
);

INVX1 _23303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .Y(_1666_)
);

AND2X2 _16097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_24_bF$buf5),
    .Y(_5679_)
);

FILL SFILL49080x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8491_),
    .Y(_8492_)
);

AOI21X1 _18243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8030_),
    .B(_8031_),
    .C(_8028_),
    .Y(_8032_)
);

FILL SFILL18600x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10887_),
    .B(_10886_),
    .C(_10883_),
    .Y(_10888_)
);

AOI21X1 _20428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10139_),
    .B(_10137_),
    .C(_10183_),
    .Y(_10427_)
);

NAND3X1 _20008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9640_),
    .B(_9962_),
    .C(_9963_),
    .Y(_9967_)
);

OAI21X1 _19868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9809_),
    .B(_9810_),
    .C(_9813_),
    .Y(_9814_)
);

OAI21X1 _19448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9351_),
    .B(_9350_),
    .C(_9352_),
    .Y(_9353_)
);

NOR2X1 _19028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf3),
    .B(_7225__bF$buf3),
    .Y(_8892_)
);

NAND3X1 _14583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4014_),
    .B(_4015_),
    .C(_3867_),
    .Y(_4022_)
);

NOR2X1 _14163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .B(_3262_),
    .Y(_3561_)
);

FILL SFILL39080x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_5330_),
    .C(_4974_),
    .Y(_5340_)
);

AOI21X1 _15368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4876_),
    .B(_4875_),
    .C(_4874_),
    .Y(_4881_)
);

NAND2X1 _20181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_25_bF$buf4),
    .Y(_10157_)
);

FILL SFILL23880x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_11478_)
);

OAI21X1 _17934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7688_),
    .B(_7690_),
    .C(_7685_),
    .Y(_7693_)
);

NOR2X1 _17514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_6815__bF$buf1),
    .Y(_7232_)
);

FILL SFILL8760x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _18719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8529_),
    .Y(_8553_)
);

NOR3X1 _13854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2950_),
    .B(_2951_),
    .C(_2949_),
    .Y(_3224_)
);

DFFPOSX1 _23952_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[6]),
    .CLK(clk_bF$buf7),
    .D(_0_[6])
);

INVX4 _13434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf3),
    .Y(_2763_)
);

AOI21X1 _13014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2308_),
    .B(_2307_),
    .C(_2300_),
    .Y(_2309_)
);

NAND2X1 _23532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .B(_1893_),
    .Y(_1916_)
);

NAND2X1 _23112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1356_),
    .Y(_1458_)
);

FILL SFILL53960x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4080_),
    .B(_4077_),
    .C(_4075_),
    .Y(_4081_)
);

NAND3X1 _14219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3614_),
    .B(_3617_),
    .C(_3600_),
    .Y(_3622_)
);

AOI21X1 _18892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7935_),
    .B(_8743_),
    .C(_8350_),
    .Y(_8744_)
);

NAND2X1 _18472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_19_bF$buf4),
    .Y(_8284_)
);

AND2X2 _18052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf2),
    .B(areg_17_bF$buf3),
    .Y(_7823_)
);

OAI22X1 _20657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10323_),
    .B(_10328_),
    .C(_10677_),
    .D(_10676_),
    .Y(_10678_)
);

INVX2 _20237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10216_),
    .Y(_10217_)
);

FILL SFILL43960x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _11920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_2453_),
    .Y(_2475_)
);

AOI21X1 _19677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9604_),
    .B(_9599_),
    .C(_9274_),
    .Y(_9605_)
);

NAND2X1 _19257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_27_bF$buf2),
    .Y(_9144_)
);

AND2X2 _14392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_16_bF$buf1),
    .Y(_3812_)
);

DFFPOSX1 _24070_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[28]),
    .CLK(clk_bF$buf5),
    .D(b[28])
);

OAI21X1 _12705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10968_),
    .B(_10979_),
    .C(_10803_),
    .Y(_11077_)
);

NAND3X1 _22803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1117_),
    .B(_1114_),
    .C(_1120_),
    .Y(_1121_)
);

XNOR2X1 _15597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5130_),
    .Y(_5131_)
);

NAND2X1 _15177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4667_),
    .B(_4670_),
    .Y(_4671_)
);

NAND2X1 _21195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11268_),
    .B(_11267_),
    .Y(_11269_)
);

AOI21X1 _17743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7134_),
    .B(_7129_),
    .C(_7093_),
    .Y(_7484_)
);

XNOR2X1 _17323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7022_),
    .B(_7017_),
    .Y(_7023_)
);

NAND3X1 _18948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8799_),
    .B(_8800_),
    .C(_8798_),
    .Y(_8805_)
);

NAND3X1 _18528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8335_),
    .B(_8343_),
    .C(_8344_),
    .Y(_8345_)
);

NAND2X1 _18108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_7884_)
);

NOR2X1 _13663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3013_),
    .B(_2771_),
    .Y(_3014_)
);

INVX2 _13243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2553_),
    .Y(_2554_)
);

NOR2X1 _23761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2152_),
    .Y(_2164_)
);

XNOR2X1 _23341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1706_),
    .B(_1702_),
    .Y(_1708_)
);

FILL SFILL8920x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4058_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4333_)
);

XNOR2X1 _14448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3872_),
    .B(_3869_),
    .Y(_3873_)
);

OAI21X1 _14028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_3146__bF$buf3),
    .C(_3400_),
    .Y(_3413_)
);

FILL SFILL23880x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8050_),
    .B(_7661_),
    .C(_8042_),
    .Y(_8074_)
);

AOI21X1 _20886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10921_),
    .B(_10920_),
    .C(_10918_),
    .Y(_10930_)
);

FILL SFILL23800x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10124_),
    .B(_10118_),
    .C(_10127_),
    .Y(_10469_)
);

INVX2 _20046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10007_),
    .Y(_10008_)
);

FILL SFILL8840x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9333_),
    .B(_9394_),
    .Y(_9395_)
);

OAI21X1 _19066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8568_),
    .B(_8570_),
    .C(_8560_),
    .Y(_8934_)
);

FILL SFILL8760x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1663_),
    .Y(_1674_)
);

NAND2X1 _12514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_8_bF$buf1),
    .Y(_8983_)
);

NAND3X1 _22612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(_903_),
    .C(_898_),
    .Y(_913_)
);

FILL SFILL29000x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3069_),
    .Y(_3075_)
);

NAND3X1 _23817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_29_bF$buf2),
    .B(areg_31_bF$buf1),
    .C(_2072_),
    .Y(_2224_)
);

BUFX2 BUFX2_insert310 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf0)
);

BUFX2 BUFX2_insert311 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf5)
);

BUFX2 BUFX2_insert312 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf4)
);

BUFX2 BUFX2_insert313 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf3)
);

BUFX2 BUFX2_insert314 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf2)
);

NAND3X1 _17972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7731_),
    .B(_7732_),
    .C(_7734_),
    .Y(_7735_)
);

NAND2X1 _17552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6866_),
    .B(_6874_),
    .Y(_7274_)
);

BUFX2 BUFX2_insert315 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf1)
);

BUFX2 BUFX2_insert316 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044_),
    .Y(_6044__bF$buf0)
);

AND2X2 _17132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6499_),
    .B(_6493_),
    .Y(_6814_)
);

BUFX2 BUFX2_insert317 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5315__bF$buf4)
);

BUFX2 BUFX2_insert318 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5315__bF$buf3)
);

BUFX2 BUFX2_insert319 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315_),
    .Y(_5315__bF$buf2)
);

FILL SFILL23960x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8591_),
    .B(_8585_),
    .C(_8581_),
    .Y(_8595_)
);

NAND3X1 _18337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8132_),
    .B(_8134_),
    .C(_8133_),
    .Y(_8135_)
);

NAND2X1 _13892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .B(_3264_),
    .Y(_3265_)
);

FILL FILL74120x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2804_),
    .Y(_2805_)
);

DFFPOSX1 _23990_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[44]),
    .CLK(clk_bF$buf8),
    .D(_0_[44])
);

AOI21X1 _13052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_1140_),
    .C(_1162_),
    .Y(_2347_)
);

AOI21X1 _23570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6038_),
    .B(_1951_),
    .C(_1955_),
    .Y(_1956_)
);

NOR2X1 _23150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1497_),
    .Y(_1499_)
);

NOR3X1 _14677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4119_),
    .B(_4111_),
    .C(_4118_),
    .Y(_4123_)
);

AOI21X1 _14257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3648_),
    .B(_3652_),
    .C(_3653_),
    .Y(_3664_)
);

AOI21X1 _18090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7863_),
    .B(_7862_),
    .C(_7861_),
    .Y(_7864_)
);

OAI21X1 _20695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_10709_),
    .Y(_10720_)
);

NOR2X1 _20275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10259_),
    .B(_10258_),
    .Y(_10260_)
);

AOI21X1 _16823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6468_),
    .B(_6469_),
    .C(_6467_),
    .Y(_6475_)
);

OAI21X1 _16403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6013_),
    .B(_6014_),
    .C(_6011_),
    .Y(_6015_)
);

NOR2X1 _19295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8816_),
    .B(_8783_),
    .Y(_9186_)
);

NAND3X1 _17608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7224_),
    .B(_7329_),
    .C(_7334_),
    .Y(_7335_)
);

FILL SFILL59160x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11417_),
    .B(_11483_),
    .C(_9959_),
    .Y(_11494_)
);

AOI21X1 _12323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6703_),
    .B(_6769_),
    .C(_6341_),
    .Y(_6889_)
);

NOR2X1 _22841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1156_),
    .Y(_1163_)
);

AOI21X1 _22421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_475_),
    .C(_702_),
    .Y(_704_)
);

OAI21X1 _22001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(_11891_),
    .C(_21_),
    .Y(_243_)
);

FILL SFILL8920x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf3),
    .B(areg_10_bF$buf0),
    .Y(_3326_)
);

AOI21X1 _13528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2852_),
    .B(_2848_),
    .C(_2855_),
    .Y(_2866_)
);

NAND3X1 _13108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2403_),
    .B(_2404_),
    .C(_2405_),
    .Y(_2406_)
);

XNOR2X1 _23626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_2010_),
    .Y(_2018_)
);

NOR2X1 _23206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf2),
    .B(_6815__bF$buf4),
    .Y(_1560_)
);

OAI21X1 _17781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7524_),
    .B(_7523_),
    .C(_7515_),
    .Y(_7526_)
);

AND2X2 _17361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6660_),
    .B(_6656_),
    .Y(_7066_)
);

OAI21X1 _18986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8839_),
    .B(_8845_),
    .C(_8482_),
    .Y(_8846_)
);

OAI21X1 _18566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8356_),
    .B(_8357_),
    .C(_8334_),
    .Y(_8386_)
);

NAND2X1 _18146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7921_),
    .B(_7925_),
    .Y(_7926_)
);

NOR2X1 _13281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf3),
    .B(_8555_),
    .Y(_2595_)
);

OAI21X1 _14486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3666_),
    .B(_3914_),
    .C(_3711_),
    .Y(_3915_)
);

AOI21X1 _14066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3454_),
    .B(_3453_),
    .C(_3446_),
    .Y(_3455_)
);

FILL SFILL8680x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10047_),
    .B(_10048_),
    .Y(_10050_)
);

INVX1 _16632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5893_),
    .Y(_6266_)
);

AOI21X1 _16212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5048_),
    .B(_5785_),
    .C(_5424_),
    .Y(_5806_)
);

OAI21X1 _21289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11065_),
    .B(_11061_),
    .C(_11069_),
    .Y(_11371_)
);

AOI21X1 _17837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7566_),
    .B(_7572_),
    .C(_7483_),
    .Y(_7587_)
);

AOI21X1 _17417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7114_),
    .B(_7112_),
    .C(_7110_),
    .Y(_7127_)
);

NOR2X1 _12972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1913_),
    .B(_286_),
    .Y(_2088_)
);

NAND3X1 _12552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9236_),
    .B(_8950_),
    .C(_9279_),
    .Y(_9400_)
);

NAND3X1 _12132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3460_),
    .B(_4785_),
    .C(_4697_),
    .Y(_4796_)
);

INVX1 _22650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .Y(_953_)
);

OAI21X1 _22230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_283_),
    .B(_252_),
    .C(_291_),
    .Y(_493_)
);

FILL SFILL54120x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2872_),
    .B(_2873_),
    .Y(_3117_)
);

AND2X2 _13337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .B(_2655_),
    .Y(_2657_)
);

NAND2X1 _23855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2244_),
    .B(_2253_),
    .Y(_2264_)
);

NAND2X1 _23435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_26_bF$buf1),
    .B(areg_28_bF$buf4),
    .Y(_1810_)
);

NAND2X1 _23015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf4),
    .B(areg_31_bF$buf2),
    .Y(_1352_)
);

NOR3X1 _17590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6886_),
    .B(_6883_),
    .C(_6884_),
    .Y(_7315_)
);

NAND2X1 _17170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6853_),
    .B(_6854_),
    .Y(_6855_)
);

INVX2 _15903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5466_),
    .Y(_5467_)
);

AND2X2 _18795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf3),
    .B(areg_18_bF$buf5),
    .Y(_8637_)
);

FILL SFILL54040x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7783_),
    .B(_7867_),
    .C(_7875_),
    .Y(_8177_)
);

AND2X2 _13090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2383_),
    .Y(_2386_)
);

AOI21X1 _21921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11755_),
    .B(_11779_),
    .C(_11782_),
    .Y(_156_)
);

NAND2X1 _21501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11411_),
    .B(_11419_),
    .Y(_11604_)
);

NAND3X1 _14295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3704_),
    .B(_3705_),
    .C(_3703_),
    .Y(_3706_)
);

AOI21X1 _12608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9367_),
    .B(_9411_),
    .C(_8709_),
    .Y(_10013_)
);

AOI21X1 _22706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1003_),
    .B(_997_),
    .C(_981_),
    .Y(_1015_)
);

FILL SFILL8520x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _16861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6515_),
    .B(_6513_),
    .Y(_6517_)
);

AOI21X1 _16441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5704_),
    .C(_5706_),
    .Y(_6056_)
);

AOI21X1 _16021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5578_),
    .B(_5583_),
    .C(_5539_),
    .Y(_5597_)
);

XNOR2X1 _21098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11137_),
    .B(_11161_),
    .Y(_11162_)
);

AOI21X1 _17646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7376_),
    .B(_7375_),
    .C(_7374_),
    .Y(_7377_)
);

OAI21X1 _17226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6909_),
    .B(_6910_),
    .C(_6907_),
    .Y(_6917_)
);

NAND3X1 _12781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11876_),
    .B(_11898_),
    .C(_11887_),
    .Y(_1_)
);

NOR2X1 _12361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .B(_6220_),
    .Y(_7305_)
);

OAI21X1 _13986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf1),
    .B(_549__bF$buf4),
    .C(_3359_),
    .Y(_3367_)
);

NOR3X1 _13566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2907_),
    .B(_2906_),
    .C(_2903_),
    .Y(_2908_)
);

OAI21X1 _13146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2303_),
    .C(_2293_),
    .Y(_2448_)
);

INVX1 _23664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .Y(_2059_)
);

NAND2X1 _23244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_1601_),
    .Y(_1602_)
);

FILL SFILL24040x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24029_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[19]),
    .CLK(clk_bF$buf5),
    .D(a[19])
);

AOI21X1 _15712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4914_),
    .B(_4766_),
    .C(_4920_),
    .Y(_5258_)
);

NOR2X1 _18184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7116_),
    .B(_7967_),
    .Y(_7968_)
);

FILL SFILL59160x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf5),
    .B(areg_22_bF$buf3),
    .Y(_10823_)
);

OAI22X1 _20369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf3),
    .B(_6050__bF$buf2),
    .C(_10869__bF$buf1),
    .D(_5668__bF$buf0),
    .Y(_10362_)
);

AOI21X1 _16917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6164_),
    .B(_6185_),
    .C(_6189_),
    .Y(_6578_)
);

AOI21X1 _21730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11853_),
    .B(_11849_),
    .C(_11598_),
    .Y(_11854_)
);

INVX1 _21310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11371_),
    .Y(_11394_)
);

AND2X2 _19389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_27_bF$buf2),
    .Y(_9288_)
);

FILL SFILL54120x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_571_),
    .B(_604_),
    .C(_494_),
    .Y(_615_)
);

OAI21X1 _12417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7898_),
    .B(_7909_),
    .C(_7887_),
    .Y(_7920_)
);

OAI21X1 _22935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1229_),
    .B(_1103_),
    .C(_1231_),
    .Y(_1265_)
);

AOI21X1 _22515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_794_),
    .C(_774_),
    .Y(_806_)
);

OAI21X1 _16670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5930_),
    .B(_5934_),
    .C(_5933_),
    .Y(_6307_)
);

NAND2X1 _16250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_16_bF$buf1),
    .Y(_5847_)
);

FILL SFILL58840x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7219_),
    .B(_7622_),
    .C(_7628_),
    .Y(_7629_)
);

OAI21X1 _17455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7167_),
    .B(_7168_),
    .C(_7166_),
    .Y(_7169_)
);

NAND3X1 _17035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6694_),
    .B(_6707_),
    .C(_6702_),
    .Y(_6708_)
);

NAND3X1 _12590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9784_),
    .B(_9795_),
    .C(_9806_),
    .Y(_9817_)
);

OAI21X1 _12170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4390_),
    .B(_5179_),
    .C(_5201_),
    .Y(_5212_)
);

NAND2X1 _13795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_3159_)
);

AOI21X1 _13375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2492_),
    .B(_2491_),
    .C(_2487_),
    .Y(_2699_)
);

BUFX2 _23893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[11]),
    .Y(y[11])
);

AOI21X1 _23473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1847_),
    .B(_1846_),
    .C(_1738_),
    .Y(_1852_)
);

NAND3X1 _23053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .B(_1388_),
    .C(_1389_),
    .Y(_1394_)
);

OAI21X1 _19601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9518_),
    .B(_9519_),
    .C(_9520_),
    .Y(_9522_)
);

NAND3X1 _15941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5498_),
    .B(_5491_),
    .C(_5495_),
    .Y(_5509_)
);

AND2X2 _15521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_15_bF$buf5),
    .Y(_5048_)
);

OAI21X1 _15101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4581_),
    .B(_4582_),
    .C(_4497_),
    .Y(_4589_)
);

FILL SFILL34040x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10613_),
    .B(_10612_),
    .Y(_10614_)
);

OAI21X1 _20178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf2),
    .B(_4551__bF$buf0),
    .C(_10149_),
    .Y(_10153_)
);

OAI21X1 _16726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6367_),
    .B(_6368_),
    .C(_6366_),
    .Y(_6369_)
);

OAI21X1 _16306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5902_),
    .B(_5904_),
    .C(_5905_),
    .Y(_5909_)
);

FILL SFILL69240x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9037_),
    .B(_9033_),
    .Y(_9079_)
);

OAI21X1 _12646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8939_),
    .B(_9290_),
    .C(_9400_),
    .Y(_10430_)
);

FILL SFILL59240x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5792_),
    .B(_5771_),
    .C(_4215_),
    .Y(_5826_)
);

AND2X2 _22744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .B(_1054_),
    .Y(_1057_)
);

NAND3X1 _22324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_594_),
    .B(_595_),
    .C(_596_),
    .Y(_597_)
);

FILL SFILL3800x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23949_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[3]),
    .CLK(clk_bF$buf2),
    .D(_0_[3])
);

XNOR2X1 _23529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .B(_1910_),
    .Y(_1911_)
);

XNOR2X1 _23109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .B(_1451_),
    .Y(_1454_)
);

NAND3X1 _17684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7417_),
    .B(_7418_),
    .C(_7416_),
    .Y(_7419_)
);

OAI21X1 _17264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6958_),
    .B(_6573_),
    .C(_6564_),
    .Y(_6959_)
);

FILL SFILL59160x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL9000x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10828_),
    .B(_10833_),
    .C(_10835_),
    .Y(_10846_)
);

NAND2X1 _18889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8735_),
    .B(_8739_),
    .Y(_8740_)
);

AOI21X1 _18469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7994_),
    .B(_7995_),
    .C(_7928_),
    .Y(_8280_)
);

AOI21X1 _18049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6964_),
    .B(_7818_),
    .C(_7396_),
    .Y(_7819_)
);

AOI21X1 _13184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .B(_2434_),
    .C(_2425_),
    .Y(_2490_)
);

AOI21X1 _23282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1641_),
    .C(_1549_),
    .Y(_1644_)
);

NAND3X1 _19830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9767_),
    .B(_9771_),
    .C(_9770_),
    .Y(_9772_)
);

NOR3X1 _19410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9308_),
    .B(_9309_),
    .C(_9310_),
    .Y(_9311_)
);

NAND2X1 _11917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf3),
    .B(areg_2_bF$buf2),
    .Y(_2442_)
);

OAI21X1 _14389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3562_),
    .B(_3807_),
    .C(_3553_),
    .Y(_3808_)
);

DFFPOSX1 _24067_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[25]),
    .CLK(clk_bF$buf4),
    .D(b[25])
);

FILL SFILL18760x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5295_),
    .B(_5297_),
    .Y(_5298_)
);

OAI21X1 _15330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4835_),
    .B(_4836_),
    .C(_4838_),
    .Y(_4839_)
);

FILL SFILL64040x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6229_),
    .B(_6613_),
    .Y(_6620_)
);

OAI21X1 _16535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6145_),
    .B(_6149_),
    .C(_6151_),
    .Y(_6159_)
);

OAI21X1 _16115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5695_),
    .B(_5696_),
    .C(_5698_),
    .Y(_5699_)
);

OAI21X1 _12875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1009_),
    .B(_1020_),
    .C(_976_),
    .Y(_1031_)
);

OAI21X1 _12455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5859_),
    .B(_7087_),
    .C(_7020_),
    .Y(_8337_)
);

OR2X2 _22973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1305_),
    .Y(_1306_)
);

NAND2X1 _12035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3612_),
    .B(_3701_),
    .Y(_3734_)
);

NAND2X1 _22553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_846_),
    .Y(_848_)
);

INVX1 _22133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .Y(_388_)
);

FILL SFILL69320x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2159_),
    .B(_2119_),
    .Y(_2161_)
);

NOR2X1 _23338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1578_),
    .B(_1703_),
    .Y(_1704_)
);

AOI22X1 _14601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3519_),
    .B(_3774_),
    .C(_4040_),
    .D(_4036_),
    .Y(_4041_)
);

OAI21X1 _17493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7205_),
    .B(_7206_),
    .C(_6810_),
    .Y(_7210_)
);

NAND3X1 _17073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6742_),
    .B(_6749_),
    .C(_6602_),
    .Y(_6750_)
);

NAND3X1 _15806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4996_),
    .B(_5359_),
    .C(_5356_),
    .Y(_5360_)
);

NAND2X1 _18698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_26_bF$buf2),
    .Y(_8530_)
);

OAI21X1 _18278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8064_),
    .B(_7657_),
    .C(_8055_),
    .Y(_8070_)
);

NAND3X1 _23091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1409_),
    .B(_1433_),
    .C(_1432_),
    .Y(_1435_)
);

FILL SFILL59240x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_28_),
    .B(_42_),
    .C(_48_),
    .Y(_49_)
);

NAND3X1 _21404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11482_),
    .B(_11486_),
    .C(_11493_),
    .Y(_11498_)
);

AOI21X1 _14198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3324_),
    .B(_3328_),
    .C(_3332_),
    .Y(_3599_)
);

NOR3X1 _22609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_679_),
    .C(_686_),
    .Y(_909_)
);

FILL FILL74200x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6409_),
    .B(_6410_),
    .C(_6405_),
    .Y(_6411_)
);

OAI21X1 _16344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5946_),
    .B(_5945_),
    .C(_5929_),
    .Y(_5951_)
);

BUFX2 BUFX2_insert280 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf2)
);

BUFX2 BUFX2_insert281 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf1)
);

BUFX2 BUFX2_insert282 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf0)
);

BUFX2 BUFX2_insert283 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf5)
);

BUFX2 BUFX2_insert284 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf4)
);

INVX1 _17969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7710_),
    .Y(_7731_)
);

AND2X2 _17549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7266_),
    .B(_7269_),
    .Y(_7270_)
);

BUFX2 BUFX2_insert285 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf3)
);

BUFX2 BUFX2_insert286 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf2)
);

NAND2X1 _17129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6778_),
    .B(_6787_),
    .Y(_6810_)
);

BUFX2 BUFX2_insert287 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf1)
);

BUFX2 BUFX2_insert288 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453_),
    .Y(_5453__bF$buf0)
);

AND2X2 _12684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_12_bF$buf1),
    .Y(_10847_)
);

BUFX2 BUFX2_insert289 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(breg_9_bF$buf5)
);

NOR2X1 _12264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6132_),
    .B(_6231_),
    .Y(_6242_)
);

OAI21X1 _22782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1097_),
    .B(_1085_),
    .C(_1083_),
    .Y(_1098_)
);

OAI21X1 _22362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(_625_),
    .C(_618_),
    .Y(_639_)
);

NAND3X1 _18910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8744_),
    .B(_8756_),
    .C(_8762_),
    .Y(_8763_)
);

NOR2X1 _13889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf1),
    .B(_2763_),
    .Y(_3261_)
);

NAND2X1 _13469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_9_bF$buf2),
    .Y(_2801_)
);

DFFPOSX1 _23987_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[41]),
    .CLK(clk_bF$buf7),
    .D(_0_[41])
);

NAND3X1 _13049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_2342_),
    .C(_2343_),
    .Y(_2344_)
);

NAND3X1 _23567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7633_),
    .B(_7637_),
    .C(_7213_),
    .Y(_1953_)
);

NAND2X1 _23147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf4),
    .B(areg_30_bF$buf4),
    .Y(_1496_)
);

OAI21X1 _14830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4284_),
    .B(_4285_),
    .C(_4202_),
    .Y(_4291_)
);

OAI21X1 _14410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3829_),
    .B(_3830_),
    .C(_3823_),
    .Y(_3831_)
);

FILL SFILL33800x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_18_bF$buf4),
    .Y(_5151_)
);

NOR2X1 _18087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7859_),
    .B(_7860_),
    .Y(_7861_)
);

XNOR2X1 _11955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2847_),
    .B(_2803_),
    .Y(_2858_)
);

NAND3X1 _21633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11742_),
    .B(_11727_),
    .C(_11743_),
    .Y(_11748_)
);

AOI21X1 _21213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11287_),
    .B(_11288_),
    .C(_11010_),
    .Y(_11289_)
);

NAND2X1 _22838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1156_),
    .Y(_1159_)
);

AOI21X1 _22418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_698_),
    .C(_493_),
    .Y(_700_)
);

OAI21X1 _16993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf0),
    .B(_4551__bF$buf1),
    .C(_6655_),
    .Y(_6662_)
);

OR2X2 _16573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6160_),
    .B(_6156_),
    .Y(_6201_)
);

OAI21X1 _16153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5733_),
    .B(_5734_),
    .C(_5731_),
    .Y(_5741_)
);

NAND3X1 _17778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7516_),
    .B(_7521_),
    .C(_7519_),
    .Y(_7522_)
);

NAND2X1 _17358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7057_),
    .B(_7061_),
    .Y(_7062_)
);

FILL SFILL43880x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_6_bF$buf2),
    .Y(_8753_)
);

AND2X2 _12073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4105_),
    .B(_4138_),
    .Y(_4149_)
);

AOI21X1 _22591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_672_),
    .B(_888_),
    .C(_731_),
    .Y(_890_)
);

AOI21X1 _22171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_425_),
    .B(_424_),
    .C(_423_),
    .Y(_430_)
);

FILL SFILL8600x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10944_),
    .B(_10949_),
    .Y(_10950_)
);

INVX1 _13698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3051_),
    .Y(_3052_)
);

NOR2X1 _13278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_2591_),
    .Y(_2592_)
);

AND2X2 _23796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2200_),
    .B(_2201_),
    .Y(_2202_)
);

NAND3X1 _23376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1745_),
    .B(_1744_),
    .C(_1743_),
    .Y(_1746_)
);

NAND3X1 _19924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9870_),
    .B(_9862_),
    .C(_9875_),
    .Y(_9876_)
);

NOR3X1 _19504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9401_),
    .B(_9409_),
    .C(_9410_),
    .Y(_9415_)
);

FILL FILL74200x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5388_),
    .B(_5392_),
    .C(_5379_),
    .Y(_5402_)
);

OAI21X1 _15424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4941_),
    .B(_4942_),
    .C(_4940_),
    .Y(_4943_)
);

NAND3X1 _15004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4480_),
    .B(_4481_),
    .C(_4479_),
    .Y(_4482_)
);

NAND2X1 _16629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6261_),
    .B(_6257_),
    .Y(_6262_)
);

AOI21X1 _16209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5467_),
    .B(_5469_),
    .C(_5801_),
    .Y(_5802_)
);

OAI21X1 _21862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_83_),
    .C(_81_),
    .Y(_91_)
);

INVX1 _21442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11539_),
    .Y(_11540_)
);

NOR2X1 _21022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10755_),
    .B(_10818_),
    .Y(_11079_)
);

FILL SFILL13880x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .Y(_2055_)
);

FILL SFILL13480x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9356_),
    .B(_9290_),
    .C(_8939_),
    .Y(_9367_)
);

AOI21X1 _12129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4752_),
    .B(_4741_),
    .C(_4653_),
    .Y(_4763_)
);

NAND2X1 _22647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_822_),
    .Y(_950_)
);

OAI21X1 _22227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11878_),
    .B(_11873_),
    .C(_489_),
    .Y(_490_)
);

OAI21X1 _13910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3282_),
    .B(_3283_),
    .C(_3281_),
    .Y(_3284_)
);

NAND2X1 _16382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5989_),
    .B(_5991_),
    .Y(_5992_)
);

FILL SFILL8680x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7303_),
    .B(_7304_),
    .C(_7301_),
    .Y(_7312_)
);

INVX1 _17167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6851_),
    .Y(_6852_)
);

FILL SFILL8600x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10735_),
    .B(_10739_),
    .Y(_10740_)
);

OAI22X1 _13087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2379_),
    .C(_2382_),
    .D(_2380_),
    .Y(_2383_)
);

XNOR2X1 _23185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1402_),
    .B(_1537_),
    .Y(_0_[51])
);

AOI21X1 _19733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9286_),
    .B(_9291_),
    .C(_9294_),
    .Y(_9666_)
);

OAI21X1 _19313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9093_),
    .B(_9091_),
    .C(_9006_),
    .Y(_9206_)
);

OAI21X1 _21918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .B(_143_),
    .C(_141_),
    .Y(_152_)
);

FILL SFILL74280x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5192_),
    .B(_5187_),
    .Y(_5193_)
);

FILL SFILL13960x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4727_),
    .B(_4728_),
    .C(_4732_),
    .Y(_4733_)
);

FILL SFILL74200x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf3),
    .B(_5369_),
    .Y(_6513_)
);

OAI21X1 _16438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf2),
    .B(_6050__bF$buf2),
    .C(_6051_),
    .Y(_6052_)
);

NOR3X1 _16018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5220_),
    .B(_5221_),
    .C(_5219_),
    .Y(_5593_)
);

NAND2X1 _11993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3252_),
    .B(_3263_),
    .Y(_3274_)
);

OAI21X1 _21671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11774_),
    .B(_11775_),
    .C(_11769_),
    .Y(_11790_)
);

OAI21X1 _21251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11034_),
    .B(_11020_),
    .C(_11045_),
    .Y(_11330_)
);

FILL SFILL64280x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11745_),
    .Y(_11876_)
);

XNOR2X1 _12358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7261_),
    .B(_7250_),
    .Y(_7272_)
);

NOR2X1 _22876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(_1045_),
    .Y(_1201_)
);

OAI21X1 _22456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf0),
    .B(_5668__bF$buf1),
    .C(_510_),
    .Y(_741_)
);

NAND3X1 _22036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_257_),
    .C(_270_),
    .Y(_281_)
);

OAI21X1 _16191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5406_),
    .B(_5781_),
    .C(_5415_),
    .Y(_5782_)
);

FILL SFILL33720x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_16_bF$buf2),
    .Y(_4394_)
);

AOI21X1 _14504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3926_),
    .B(_3927_),
    .C(_3925_),
    .Y(_3935_)
);

AND2X2 _17396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7096_),
    .B(_7097_),
    .Y(_7104_)
);

AOI21X1 _15709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5235_),
    .B(_5241_),
    .C(_5103_),
    .Y(_5254_)
);

AOI21X1 _20942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10989_),
    .B(_10991_),
    .C(_10690_),
    .Y(_10992_)
);

OAI21X1 _20522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10515_),
    .B(_10516_),
    .C(_10513_),
    .Y(_10531_)
);

NAND3X1 _20102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10066_),
    .B(_10067_),
    .C(_10069_),
    .Y(_10070_)
);

AOI22X1 _19962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9913_),
    .B(_9916_),
    .C(_9896_),
    .D(_9900_),
    .Y(_9917_)
);

AOI21X1 _19542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9066_),
    .B(_9068_),
    .C(_9074_),
    .Y(_9457_)
);

OAI21X1 _19122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8993_),
    .B(_8992_),
    .C(_8995_),
    .Y(_8996_)
);

FILL SFILL23720x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11600_),
    .B(_11846_),
    .C(_11847_),
    .Y(_11851_)
);

AOI21X1 _21307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11161_),
    .B(_11136_),
    .C(_11390_),
    .Y(_11391_)
);

NAND3X1 _15882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .B(_5443_),
    .C(_5404_),
    .Y(_5444_)
);

AOI21X1 _15462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4693_),
    .B(_4696_),
    .C(_4685_),
    .Y(_4983_)
);

AOI21X1 _15042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4507_),
    .B(_4512_),
    .C(_4514_),
    .Y(_4524_)
);

FILL SFILL8680x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6296_),
    .B(_6298_),
    .Y(_6304_)
);

OAI21X1 _16247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5795_),
    .B(_5842_),
    .C(_5843_),
    .Y(_5844_)
);

OAI21X1 _21480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11566_),
    .B(_11569_),
    .C(_11573_),
    .Y(_11581_)
);

AOI21X1 _21060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11103_),
    .B(_11109_),
    .C(_11057_),
    .Y(_11120_)
);

FILL SFILL8600x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7065_),
    .B(_9718_),
    .C(_9773_),
    .Y(_9784_)
);

NAND2X1 _12167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_8_bF$buf1),
    .Y(_5179_)
);

NAND2X1 _22685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_991_),
    .B(_986_),
    .Y(_992_)
);

AOI21X1 _22265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_526_),
    .C(_506_),
    .Y(_532_)
);

NAND2X1 _18813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_21_bF$buf3),
    .Y(_8657_)
);

FILL SFILL74280x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4179_),
    .B(_4180_),
    .C(_4163_),
    .Y(_4185_)
);

OAI21X1 _14313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3714_),
    .B(_3707_),
    .C(_3716_),
    .Y(_3726_)
);

FILL SFILL74200x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5504_),
    .B(_5499_),
    .C(_5465_),
    .Y(_5505_)
);

NAND2X1 _15518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf3),
    .B(breg_17_bF$buf4),
    .Y(_5044_)
);

INVX2 _20751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10742_),
    .Y(_10782_)
);

NAND3X1 _20331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10318_),
    .B(_10319_),
    .C(_10320_),
    .Y(_10322_)
);

OAI21X1 _19771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf3),
    .B(_3781__bF$buf1),
    .C(_9333_),
    .Y(_9708_)
);

AOI21X1 _19351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9245_),
    .B(_9246_),
    .C(_8882_),
    .Y(_9248_)
);

NAND2X1 _21956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11829_),
    .B(_186_),
    .Y(_194_)
);

OAI21X1 _21536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11641_),
    .B(_11637_),
    .C(_11606_),
    .Y(_11642_)
);

AND2X2 _21116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10865_),
    .B(_10912_),
    .Y(_11182_)
);

FILL SFILL64200x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5231_),
    .B(_5232_),
    .C(_5230_),
    .Y(_5234_)
);

OAI21X1 _15271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4465_),
    .B(_4455_),
    .C(_4459_),
    .Y(_4775_)
);

OAI21X1 _16896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf0),
    .B(_2362__bF$buf3),
    .C(_6547_),
    .Y(_6555_)
);

AOI21X1 _16476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5777_),
    .B(_5775_),
    .C(_6093_),
    .Y(_6094_)
);

AOI21X1 _16056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5007_),
    .B(_5263_),
    .C(_5266_),
    .Y(_5635_)
);

FILL SFILL58920x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_10_bF$buf4),
    .Y(_7689_)
);

NAND2X1 _22494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf0),
    .B(breg_24_bF$buf2),
    .Y(_783_)
);

OAI21X1 _22074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_314_),
    .C(_312_),
    .Y(_323_)
);

OAI21X1 _18622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8443_),
    .B(_8447_),
    .C(_8074_),
    .Y(_8448_)
);

NAND3X1 _18202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7982_),
    .B(_7983_),
    .C(_7957_),
    .Y(_7988_)
);

AOI21X1 _20807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10834_),
    .B(_10842_),
    .C(_10820_),
    .Y(_10843_)
);

XNOR2X1 _23699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_2061_),
    .Y(_2097_)
);

AOI21X1 _23279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1635_),
    .B(_1639_),
    .C(_1550_),
    .Y(_1640_)
);

AND2X2 _19827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf2),
    .B(areg_19_bF$buf4),
    .Y(_9769_)
);

AOI21X1 _19407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8896_),
    .B(_8920_),
    .C(_8918_),
    .Y(_9308_)
);

AOI21X1 _14962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4419_),
    .B(_4426_),
    .C(_4388_),
    .Y(_4436_)
);

NAND3X1 _14542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3970_),
    .B(_3971_),
    .C(_3976_),
    .Y(_3977_)
);

AOI21X1 _14122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3509_),
    .B(_3515_),
    .C(_3513_),
    .Y(_3516_)
);

NAND2X1 _15747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5295_),
    .B(_5292_),
    .Y(_5296_)
);

AOI21X1 _15327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4823_),
    .B(_4822_),
    .C(_4819_),
    .Y(_4836_)
);

NOR2X1 _20980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11025_),
    .B(_11026_),
    .Y(_11032_)
);

OAI21X1 _20560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10571_),
    .B(_10567_),
    .C(_10563_),
    .Y(_10572_)
);

NAND2X1 _20140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_10111_)
);

FILL SFILL48840x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9107_),
    .B(_9497_),
    .Y(_9498_)
);

OAI21X1 _19160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9035_),
    .B(_9036_),
    .C(_9034_),
    .Y(_9037_)
);

OAI21X1 _21765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11624_),
    .B(_11609_),
    .C(_11634_),
    .Y(_11892_)
);

NAND3X1 _21345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11326_),
    .B(_11426_),
    .C(_11432_),
    .Y(_11433_)
);

FILL SFILL33720x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4241_),
    .B(_4257_),
    .C(_4564_),
    .Y(_4565_)
);

FILL SFILL3960x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3172_),
    .B(_3175_),
    .C(_3128_),
    .Y(_3179_)
);

BUFX2 _23911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[29]),
    .Y(y[29])
);

OAI21X1 _16285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5588_),
    .B(_5885_),
    .C(_5578_),
    .Y(_5886_)
);

NAND2X1 _18851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_22_bF$buf4),
    .Y(_8699_)
);

AOI21X1 _18431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7883_),
    .B(_8237_),
    .C(_8236_),
    .Y(_8239_)
);

OAI21X1 _18011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7769_),
    .B(_7770_),
    .C(_7767_),
    .Y(_7778_)
);

NAND3X1 _20616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10616_),
    .B(_10621_),
    .C(_10460_),
    .Y(_10634_)
);

FILL SFILL28840x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1430_),
    .B(_1427_),
    .C(_1410_),
    .Y(_1431_)
);

FILL SFILL64200x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9558_),
    .B(_9559_),
    .C(_9529_),
    .Y(_9560_)
);

NAND2X1 _19216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_21_bF$buf3),
    .Y(_9098_)
);

AOI22X1 _14771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .B(_3951_),
    .C(_4225_),
    .D(_3949_),
    .Y(_4227_)
);

AOI21X1 _14351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3753_),
    .B(_3761_),
    .C(_3480_),
    .Y(_3767_)
);

OR2X2 _15976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5545_),
    .B(_5546_),
    .Y(_5547_)
);

FILL SFILL18680x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5076_),
    .B(_5077_),
    .C(_5041_),
    .Y(_5086_)
);

NAND3X1 _15136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4613_),
    .B(_4617_),
    .C(_4620_),
    .Y(_4627_)
);

FILL SFILL18840x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _21994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11879_),
    .B(_235_),
    .Y(_0_[44])
);

AOI21X1 _21574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11469_),
    .B(_11467_),
    .C(_11682_),
    .Y(_11683_)
);

AOI21X1 _21154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11222_),
    .B(_11223_),
    .C(_11221_),
    .Y(_11224_)
);

NAND2X1 _17702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf3),
    .B(areg_17_bF$buf4),
    .Y(_7439_)
);

FILL SFILL38920x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _22779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_1084_),
    .C(_1088_),
    .Y(_1094_)
);

INVX2 _22359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .Y(_635_)
);

OAI21X1 _18907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_8759_),
    .C(_8346_),
    .Y(_8760_)
);

AOI21X1 _13622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2965_),
    .B(_2966_),
    .C(_2733_),
    .Y(_2970_)
);

AOI21X1 _13202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2504_),
    .B(_2503_),
    .C(_2502_),
    .Y(_2510_)
);

OAI21X1 _23720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2118_),
    .C(_2117_),
    .Y(_2119_)
);

AOI21X1 _23300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_1633_),
    .C(_1628_),
    .Y(_1662_)
);

INVX8 _16094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_26_bF$buf0),
    .Y(_5676_)
);

NAND3X1 _14827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4155_),
    .B(_4197_),
    .C(_4198_),
    .Y(_4288_)
);

OAI21X1 _14407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf3),
    .B(_2362__bF$buf0),
    .C(_3812_),
    .Y(_3828_)
);

NAND3X1 _17299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6957_),
    .B(_6990_),
    .C(_6996_),
    .Y(_6997_)
);

INVX2 _18660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8487_),
    .Y(_8488_)
);

NAND2X1 _18240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8027_),
    .B(_8026_),
    .Y(_8028_)
);

OAI21X1 _20845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10870_),
    .B(_10871_),
    .C(_10867_),
    .Y(_10885_)
);

NAND3X1 _20425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10417_),
    .B(_10422_),
    .C(_10423_),
    .Y(_10424_)
);

AOI21X1 _20005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9962_),
    .B(_9963_),
    .C(_9640_),
    .Y(_9964_)
);

NAND2X1 _19865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_24_bF$buf1),
    .Y(_9811_)
);

AOI21X1 _19445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9344_),
    .B(_9346_),
    .C(_9343_),
    .Y(_9350_)
);

AOI21X1 _19025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8836_),
    .B(_8837_),
    .C(_8601_),
    .Y(_8889_)
);

NAND3X1 _14580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3861_),
    .B(_3859_),
    .C(_3855_),
    .Y(_4018_)
);

AOI21X1 _14160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3544_),
    .B(_3543_),
    .C(_3541_),
    .Y(_3557_)
);

AOI21X1 _15785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5035_),
    .B(_5038_),
    .C(_5082_),
    .Y(_5337_)
);

NAND3X1 _15365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4871_),
    .B(_4877_),
    .C(_4847_),
    .Y(_4878_)
);

AOI21X1 _21383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10856_),
    .B(_11474_),
    .C(_11185_),
    .Y(_11475_)
);

FILL SFILL28920x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7677_),
    .B(_7676_),
    .C(_7673_),
    .Y(_7690_)
);

NOR2X1 _17511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6831_),
    .B(_6827_),
    .Y(_7229_)
);

NAND2X1 _22588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_885_),
    .B(_881_),
    .Y(_886_)
);

NAND3X1 _22168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_425_),
    .C(_423_),
    .Y(_426_)
);

AOI21X1 _18716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8190_),
    .B(_8549_),
    .C(_8548_),
    .Y(_8550_)
);

OAI21X1 _13851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3204_),
    .B(_3211_),
    .C(_3214_),
    .Y(_3221_)
);

OAI21X1 _13431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2758_),
    .B(_2576_),
    .C(_2711_),
    .Y(_2760_)
);

AOI21X1 _13011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_659_),
    .C(_692_),
    .Y(_2306_)
);

NAND2X1 _14636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_19_bF$buf2),
    .Y(_4078_)
);

AOI21X1 _14216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3618_),
    .B(_3611_),
    .C(_3598_),
    .Y(_3619_)
);

FILL SFILL18680x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18840x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10657_),
    .B(_10658_),
    .C(_10339_),
    .Y(_10675_)
);

XNOR2X1 _20234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10213_),
    .B(_10211_),
    .Y(_10214_)
);

NAND3X1 _19674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9595_),
    .B(_9596_),
    .C(_9594_),
    .Y(_9602_)
);

NAND2X1 _19254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9135_),
    .B(_9140_),
    .Y(_9141_)
);

NAND3X1 _21859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11889_),
    .B(_82_),
    .C(_86_),
    .Y(_87_)
);

NAND2X1 _21439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11535_),
    .B(_11524_),
    .Y(_11536_)
);

NAND3X1 _21019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11067_),
    .B(_11071_),
    .C(_11074_),
    .Y(_11075_)
);

OAI21X1 _12702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11022_),
    .B(_11043_),
    .C(_11011_),
    .Y(_11044_)
);

NOR2X1 _22800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf0),
    .B(_6427_),
    .Y(_1117_)
);

OAI21X1 _15594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5126_),
    .B(_5127_),
    .C(_5122_),
    .Y(_5128_)
);

INVX1 _15174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4354_),
    .Y(_4668_)
);

NOR2X1 _13907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3280_),
    .B(_3007_),
    .Y(_3281_)
);

FILL SFILL53880x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6446_),
    .B(_6447_),
    .Y(_6448_)
);

NAND3X1 _16379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5982_),
    .B(_5987_),
    .C(_5835_),
    .Y(_5988_)
);

AOI21X1 _21192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11260_),
    .B(_11265_),
    .C(_11130_),
    .Y(_11266_)
);

AOI21X1 _17740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7464_),
    .B(_7469_),
    .C(_7471_),
    .Y(_7480_)
);

NOR2X1 _17320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6606_),
    .B(_7018_),
    .Y(_7019_)
);

NOR2X1 _12299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6472_),
    .B(_6494_),
    .Y(_6626_)
);

AOI21X1 _22397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_455_),
    .C(_675_),
    .Y(_676_)
);

FILL SFILL3560x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8794_),
    .B(_8801_),
    .C(_8694_),
    .Y(_8802_)
);

NAND3X1 _18525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8336_),
    .B(_8341_),
    .C(_8340_),
    .Y(_8342_)
);

NAND2X1 _18105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7456_),
    .B(_7464_),
    .Y(_7881_)
);

FILL SFILL59080x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2991_),
    .B(_3005_),
    .C(_3009_),
    .Y(_3010_)
);

AOI21X1 _13240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .B(_2513_),
    .C(_2361_),
    .Y(_2550_)
);

FILL SFILL38920x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4057_),
    .B(_4328_),
    .C(_4329_),
    .Y(_4330_)
);

NAND2X1 _14445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf1),
    .B(breg_13_bF$buf3),
    .Y(_3870_)
);

OAI21X1 _14025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3409_),
    .B(_3408_),
    .C(_3397_),
    .Y(_3410_)
);

FILL SFILL3560x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10916_),
    .B(_10922_),
    .C(_10926_),
    .Y(_10927_)
);

NAND2X1 _20463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .B(breg_21_bF$buf1),
    .Y(_10466_)
);

INVX2 _20043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10004_),
    .Y(_10005_)
);

FILL SFILL28920x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf2),
    .B(_5369_),
    .Y(_9392_)
);

FILL SFILL49400x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8894_),
    .B(_8922_),
    .C(_8919_),
    .Y(_8931_)
);

FILL SFILL49000x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11498_),
    .Y(_11786_)
);

NAND2X1 _21248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11103_),
    .B(_11111_),
    .Y(_11326_)
);

NAND2X1 _12931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1565_),
    .B(_1631_),
    .Y(_1642_)
);

OAI21X1 _12511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7854_),
    .B(_7832_),
    .C(_7777_),
    .Y(_8950_)
);

FILL SFILL39080x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf3),
    .B(_6044__bF$buf2),
    .C(_2807_),
    .Y(_3072_)
);

NAND2X1 _23814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2177_),
    .B(_2181_),
    .Y(_2221_)
);

NOR2X1 _16188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5774_),
    .B(_5778_),
    .Y(_5779_)
);

OAI21X1 _18754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8589_),
    .B(_8590_),
    .C(_8591_),
    .Y(_8592_)
);

INVX1 _18334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8125_),
    .Y(_8132_)
);

AOI21X1 _20939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10987_),
    .B(_10983_),
    .C(_10691_),
    .Y(_10988_)
);

NAND3X1 _20519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10497_),
    .B(_10522_),
    .C(_10526_),
    .Y(_10527_)
);

NAND2X1 _19959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9912_),
    .B(_9564_),
    .Y(_9913_)
);

OAI21X1 _19539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9443_),
    .B(_9445_),
    .C(_9441_),
    .Y(_9453_)
);

AOI21X1 _19119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8988_),
    .B(_8987_),
    .C(_8986_),
    .Y(_8992_)
);

OAI21X1 _14674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4118_),
    .B(_4119_),
    .C(_4111_),
    .Y(_4120_)
);

NAND3X1 _14254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3641_),
    .B(_3660_),
    .C(_3654_),
    .Y(_3661_)
);

AOI21X1 _15879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5438_),
    .B(_5439_),
    .C(_5432_),
    .Y(_5440_)
);

NAND2X1 _15459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4977_),
    .B(_4976_),
    .Y(_4979_)
);

OAI21X1 _15039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4516_),
    .B(_4517_),
    .C(_4519_),
    .Y(_4520_)
);

OAI21X1 _20692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10716_),
    .B(_10714_),
    .C(_10706_),
    .Y(_10717_)
);

NAND2X1 _20272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_31_bF$buf3),
    .Y(_10257_)
);

FILL SFILL74360x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _16820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6149_),
    .B(_6151_),
    .C(_6145_),
    .Y(_6471_)
);

AOI21X1 _16400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5366_),
    .B(_5625_),
    .C(_5631_),
    .Y(_6011_)
);

NAND3X1 _19292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9177_),
    .B(_9182_),
    .C(_9180_),
    .Y(_9183_)
);

INVX1 _21897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_128_),
    .Y(_129_)
);

NAND3X1 _21477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11574_),
    .B(_11577_),
    .C(_11573_),
    .Y(_11578_)
);

OAI21X1 _21057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11116_),
    .B(_10905_),
    .C(_10897_),
    .Y(_11117_)
);

NOR3X1 _17605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7006_),
    .B(_7007_),
    .C(_7005_),
    .Y(_7332_)
);

FILL SFILL59080x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11395_),
    .B(_11384_),
    .C(_11373_),
    .Y(_11461_)
);

OAI21X1 _12320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6747_),
    .B(_6758_),
    .C(_6352_),
    .Y(_6856_)
);

FILL SFILL3640x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf4),
    .B(breg_11_bF$buf3),
    .Y(_3323_)
);

NOR2X1 _13525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2427_),
    .B(_2638_),
    .Y(_2863_)
);

NAND2X1 _13105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2385_),
    .Y(_2403_)
);

AND2X2 _23623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1886_),
    .B(_2013_),
    .Y(_2015_)
);

NAND3X1 _23203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1422_),
    .C(_1415_),
    .Y(_1557_)
);

FILL SFILL49080x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8836_),
    .B(_8837_),
    .C(_8601_),
    .Y(_8843_)
);

NAND2X1 _18563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8381_),
    .B(_8382_),
    .Y(_8383_)
);

AOI21X1 _18143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7916_),
    .B(_7917_),
    .C(_7918_),
    .Y(_7923_)
);

FILL SFILL33880x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18600x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10493_),
    .B(_10491_),
    .C(_10777_),
    .Y(_10778_)
);

INVX2 _20328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9993_),
    .Y(_10318_)
);

NAND3X1 _19768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9697_),
    .B(_9701_),
    .C(_9703_),
    .Y(_9704_)
);

AOI21X1 _19348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9243_),
    .B(_9238_),
    .C(_8883_),
    .Y(_9244_)
);

OAI21X1 _14483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3911_),
    .B(_3910_),
    .C(_3908_),
    .Y(_3912_)
);

AOI21X1 _14063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3191_),
    .B(_3193_),
    .C(_3200_),
    .Y(_3452_)
);

FILL SFILL39080x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4845_),
    .B(_4883_),
    .C(_5229_),
    .Y(_5230_)
);

NAND2X1 _15268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_12_bF$buf4),
    .Y(_4771_)
);

NAND2X1 _20081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf1),
    .B(breg_25_bF$buf5),
    .Y(_10047_)
);

FILL SFILL54280x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11364_),
    .B(_11367_),
    .Y(_11368_)
);

NOR3X1 _17834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7152_),
    .B(_7154_),
    .C(_7151_),
    .Y(_7584_)
);

NAND2X1 _17414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_30_bF$buf5),
    .Y(_7124_)
);

FILL SFILL8760x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8440_),
    .B(_8441_),
    .C(_8078_),
    .Y(_8444_)
);

NAND3X1 _13754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3106_),
    .B(_3109_),
    .C(_3113_),
    .Y(_3114_)
);

INVX1 _13334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2653_),
    .Y(_2654_)
);

OAI21X1 _23852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2256_),
    .B(_2239_),
    .C(_2260_),
    .Y(_2261_)
);

INVX1 _23432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1704_),
    .Y(_1807_)
);

XOR2X1 _23012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1192_),
    .B(_1348_),
    .Y(_1349_)
);

FILL SFILL53960x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29000x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4189_),
    .B(_4196_),
    .C(_4198_),
    .Y(_4432_)
);

NOR2X1 _14539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3680_),
    .B(_3972_),
    .Y(_3973_)
);

FILL SFILL3720x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(_3511_),
    .Y(_3512_)
);

OAI21X1 _15900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5238_),
    .B(_5462_),
    .C(_5228_),
    .Y(_5463_)
);

AOI21X1 _18792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8631_),
    .B(_8633_),
    .C(_8630_),
    .Y(_8634_)
);

NAND3X1 _18372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8173_),
    .B(_8171_),
    .C(_8167_),
    .Y(_8174_)
);

NAND3X1 _20977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11024_),
    .B(_11028_),
    .C(_11027_),
    .Y(_11029_)
);

NAND3X1 _20557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10564_),
    .B(_10568_),
    .C(_10566_),
    .Y(_10569_)
);

NAND2X1 _20137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10107_),
    .B(_10103_),
    .Y(_10108_)
);

NOR3X1 _19997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9577_),
    .B(_9583_),
    .C(_9586_),
    .Y(_9955_)
);

OAI21X1 _19577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_7100__bF$buf2),
    .C(_9107_),
    .Y(_9495_)
);

XNOR2X1 _19157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9012_),
    .B(_9007_),
    .Y(_9034_)
);

AOI21X1 _14292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3418_),
    .B(_3395_),
    .C(_3702_),
    .Y(_3703_)
);

FILL SFILL43880x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64360x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9970_),
    .B(_8511_),
    .C(_9532_),
    .Y(_9981_)
);

NAND2X1 _22703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_995_),
    .Y(_1012_)
);

NAND2X1 _15497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_18_bF$buf4),
    .Y(_5021_)
);

NAND3X1 _15077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4559_),
    .B(_4560_),
    .C(_4561_),
    .Y(_4562_)
);

BUFX2 _23908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[26]),
    .Y(y[26])
);

AOI21X1 _21095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11153_),
    .B(_11158_),
    .C(_11152_),
    .Y(_11159_)
);

XNOR2X1 _17643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7350_),
    .B(_7373_),
    .Y(_7374_)
);

NAND3X1 _17223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6814_),
    .B(_6908_),
    .C(_6913_),
    .Y(_6914_)
);

FILL SFILL33880x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18600x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8312_),
    .B(_8319_),
    .Y(_8695_)
);

NAND3X1 _18428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8226_),
    .B(_8233_),
    .C(_8234_),
    .Y(_8235_)
);

NAND3X1 _18008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7664_),
    .B(_7768_),
    .C(_7773_),
    .Y(_7774_)
);

AND2X2 _13983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf5),
    .B(areg_12_bF$buf0),
    .Y(_3364_)
);

NAND3X1 _13563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2876_),
    .B(_2889_),
    .C(_2886_),
    .Y(_2905_)
);

OAI21X1 _13143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2438_),
    .C(_2433_),
    .Y(_2445_)
);

AOI21X1 _23661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1997_),
    .B(_2047_),
    .C(_2054_),
    .Y(_2056_)
);

NOR2X1 _23241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .Y(_1599_)
);

AOI21X1 _14768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4214_),
    .B(_4216_),
    .C(_4207_),
    .Y(_4223_)
);

OAI21X1 _14348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3749_),
    .C(_3755_),
    .Y(_3764_)
);

DFFPOSX1 _24026_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[16]),
    .CLK(clk_bF$buf10),
    .D(a[16])
);

FILL SFILL23880x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _18181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7963_),
    .B(_7959_),
    .Y(_7965_)
);

XNOR2X1 _20786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10819_),
    .B(_10817_),
    .Y(_10820_)
);

FILL SFILL23800x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13560x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_28_bF$buf4),
    .Y(_10359_)
);

OAI21X1 _16914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6566_),
    .C(_6563_),
    .Y(_6575_)
);

NAND2X1 _19386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_29_bF$buf3),
    .Y(_9285_)
);

FILL SFILL29080x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_13_bF$buf1),
    .Y(_582_)
);

AOI21X1 _12414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6428_),
    .B(_6637_),
    .C(_6670_),
    .Y(_7887_)
);

OAI21X1 _22932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1249_),
    .B(_1100_),
    .C(_1241_),
    .Y(_1262_)
);

NAND3X1 _22512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .B(_780_),
    .C(_785_),
    .Y(_803_)
);

FILL SFILL74440x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2953_),
    .B(_2956_),
    .C(_2960_),
    .Y(_2966_)
);

NOR2X1 _23717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2056_),
    .B(_2102_),
    .Y(_2116_)
);

AOI21X1 _17872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7620_),
    .B(_7619_),
    .C(_7618_),
    .Y(_7626_)
);

AOI21X1 _17452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6648_),
    .B(_6741_),
    .C(_7165_),
    .Y(_7166_)
);

NAND2X1 _17032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_29_bF$buf4),
    .Y(_6705_)
);

FILL SFILL3880x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _18657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8484_),
    .Y(_8485_)
);

AOI21X1 _18237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8019_),
    .B(_8024_),
    .C(_7780_),
    .Y(_8025_)
);

OAI21X1 _13792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3149_),
    .B(_3155_),
    .C(_3140_),
    .Y(_3156_)
);

NAND3X1 _13372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2679_),
    .C(_2684_),
    .Y(_2696_)
);

BUFX2 _23890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[8]),
    .Y(y[8])
);

NAND3X1 _23470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1847_),
    .C(_1846_),
    .Y(_1848_)
);

AOI21X1 _23050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1388_),
    .B(_1389_),
    .C(_1263_),
    .Y(_1390_)
);

AOI21X1 _14997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4461_),
    .B(_4459_),
    .C(_4456_),
    .Y(_4473_)
);

NAND3X1 _14577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4003_),
    .B(_3998_),
    .C(_3913_),
    .Y(_4015_)
);

NAND2X1 _14157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_16_bF$buf1),
    .Y(_3554_)
);

OAI21X1 _20595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10544_),
    .B(_10545_),
    .C(_10542_),
    .Y(_10611_)
);

NAND2X1 _20175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10148_),
    .B(_10149_),
    .Y(_10150_)
);

AOI21X1 _16723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5884_),
    .B(_5974_),
    .C(_6365_),
    .Y(_6366_)
);

NOR3X1 _16303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5904_),
    .B(_5905_),
    .C(_5902_),
    .Y(_5906_)
);

OAI21X1 _19195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9074_),
    .B(_9075_),
    .C(_9042_),
    .Y(_9076_)
);

OAI21X1 _17928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf1),
    .B(_6050__bF$buf0),
    .C(_7675_),
    .Y(_7686_)
);

INVX8 _17508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[31]),
    .Y(_7225_)
);

FILL SFILL18600x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10299_),
    .B(_10310_),
    .C(_10255_),
    .Y(_10397_)
);

NAND3X1 _12223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4215_),
    .B(_5792_),
    .C(_5771_),
    .Y(_5793_)
);

OAI21X1 _22741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_866_),
    .B(_868_),
    .C(_871_),
    .Y(_1054_)
);

NAND2X1 _22321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .B(_535_),
    .Y(_594_)
);

FILL SFILL8920x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_3216_),
    .C(_3214_),
    .Y(_3217_)
);

DFFPOSX1 _23946_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[0]),
    .CLK(clk_bF$buf0),
    .D(_0_[0])
);

NAND2X1 _13428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2572_),
    .B(_2575_),
    .Y(_2756_)
);

AOI21X1 _13008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2292_),
    .B(_2289_),
    .C(_2249_),
    .Y(_2303_)
);

NOR2X1 _23526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1905_),
    .B(_1907_),
    .Y(_1908_)
);

NAND2X1 _23106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1450_),
    .B(_1446_),
    .Y(_1451_)
);

OR2X2 _17681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7372_),
    .B(_7377_),
    .Y(_7416_)
);

AOI21X1 _17261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6954_),
    .B(_6953_),
    .C(_6952_),
    .Y(_6956_)
);

AOI21X1 _18886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8730_),
    .B(_8732_),
    .C(_8733_),
    .Y(_8737_)
);

NOR3X1 _18466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8262_),
    .B(_8266_),
    .C(_8267_),
    .Y(_8277_)
);

NAND2X1 _18046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7811_),
    .B(_7815_),
    .Y(_7816_)
);

NOR3X1 _13181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2484_),
    .B(_2485_),
    .C(_2481_),
    .Y(_2487_)
);

NAND2X1 _11914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf4),
    .B(areg_1_bF$buf3),
    .Y(_2419_)
);

NAND3X1 _14386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3782_),
    .B(_3804_),
    .C(_3803_),
    .Y(_3805_)
);

DFFPOSX1 _24064_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[22]),
    .CLK(clk_bF$buf5),
    .D(b[22])
);

FILL SFILL28840x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28760x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6612_),
    .B(_6616_),
    .C(_6614_),
    .Y(_6617_)
);

AOI21X1 _16532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6155_),
    .B(_6150_),
    .C(_6136_),
    .Y(_6156_)
);

AOI21X1 _16112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5682_),
    .B(_5680_),
    .C(_5677_),
    .Y(_5696_)
);

AOI21X1 _21189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10961_),
    .B(_11261_),
    .C(_11131_),
    .Y(_11262_)
);

NAND3X1 _17737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7472_),
    .B(_7476_),
    .C(_7438_),
    .Y(_7477_)
);

AND2X2 _17317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6630_),
    .B(_6622_),
    .Y(_7016_)
);

FILL SFILL64440x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .B(_801_),
    .C(_845_),
    .Y(_998_)
);

OAI21X1 _12452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8238_),
    .B(_8282_),
    .C(_8293_),
    .Y(_8304_)
);

OAI21X1 _22970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf1),
    .B(_5676_),
    .C(_1302_),
    .Y(_1303_)
);

XNOR2X1 _12032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3668_),
    .B(_3613_),
    .Y(_3701_)
);

NOR2X1 _22550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_842_),
    .Y(_844_)
);

OR2X2 _22130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_379_),
    .B(_383_),
    .Y(_384_)
);

FILL SFILL28680x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3006_),
    .B(_2998_),
    .Y(_3007_)
);

NAND3X1 _13237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2358_),
    .B(_2528_),
    .C(_2529_),
    .Y(_2547_)
);

NAND2X1 _23755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2157_),
    .B(_2156_),
    .Y(_2158_)
);

OAI21X1 _23335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1580_),
    .B(_1700_),
    .C(_1583_),
    .Y(_1701_)
);

AOI21X1 _17490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7191_),
    .B(_7195_),
    .C(_6811_),
    .Y(_7206_)
);

OAI21X1 _17070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6739_),
    .B(_6740_),
    .C(_6650_),
    .Y(_6746_)
);

NAND2X1 _15803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .B(_5348_),
    .Y(_5357_)
);

OAI21X1 _18695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8526_),
    .B(_8157_),
    .C(_8151_),
    .Y(_8527_)
);

XOR2X1 _18275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7652_),
    .B(_8067_),
    .Y(_0_[32])
);

OAI21X1 _21821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781__bF$buf3),
    .B(_4551__bF$buf4),
    .C(_11442_),
    .Y(_46_)
);

OAI21X1 _21401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11490_),
    .B(_11491_),
    .C(_11493_),
    .Y(_11495_)
);

NAND2X1 _14195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf1),
    .B(breg_12_bF$buf4),
    .Y(_3596_)
);

OAI21X1 _12928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf3),
    .B(_6044__bF$buf2),
    .C(_11767_),
    .Y(_1609_)
);

NAND3X1 _12508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8786_),
    .B(_8830_),
    .C(_8851_),
    .Y(_8917_)
);

OAI21X1 _22606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_897_),
    .C(_899_),
    .Y(_906_)
);

FILL SFILL44040x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6391_),
    .B(_6384_),
    .C(_6394_),
    .Y(_6408_)
);

OAI21X1 _16341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5946_),
    .B(_5945_),
    .C(_5942_),
    .Y(_5948_)
);

BUFX2 BUFX2_insert250 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf3)
);

BUFX2 BUFX2_insert251 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf2)
);

BUFX2 BUFX2_insert252 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf1)
);

BUFX2 BUFX2_insert253 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf0)
);

AOI21X1 _17966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7345_),
    .B(_7727_),
    .C(_7347_),
    .Y(_7728_)
);

BUFX2 BUFX2_insert254 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4116__bF$buf4)
);

FILL SFILL74120x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7264_),
    .B(_7263_),
    .C(_7262_),
    .Y(_7267_)
);

BUFX2 BUFX2_insert255 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4116__bF$buf3)
);

BUFX2 BUFX2_insert256 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4116__bF$buf2)
);

NOR2X1 _17126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6806_),
    .B(_6042_),
    .Y(_6807_)
);

BUFX2 BUFX2_insert257 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4116__bF$buf1)
);

BUFX2 BUFX2_insert258 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116_),
    .Y(_4116__bF$buf0)
);

NAND2X1 _12681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf2),
    .B(areg_10_bF$buf4),
    .Y(_10814_)
);

BUFX2 BUFX2_insert259 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300_),
    .Y(_6300__bF$buf3)
);

NAND2X1 _12261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6198_),
    .B(_6176_),
    .Y(_6209_)
);

FILL SFILL69160x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2999_),
    .B(_2995_),
    .C(_3004_),
    .Y(_3258_)
);

DFFPOSX1 _23984_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[38]),
    .CLK(clk_bF$buf3),
    .D(_0_[38])
);

OAI21X1 _13466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf3),
    .B(_2586__bF$buf0),
    .C(_2797_),
    .Y(_2798_)
);

XNOR2X1 _23564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_1950_),
    .Y(_0_[55])
);

NAND3X1 _13046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1173_),
    .B(_2336_),
    .C(_2340_),
    .Y(_2341_)
);

OAI21X1 _23144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1487_),
    .B(_1486_),
    .C(_1361_),
    .Y(_1493_)
);

FILL SFILL24040x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5147_),
    .B(_5142_),
    .Y(_5148_)
);

NAND3X1 _18084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7792_),
    .B(_7801_),
    .C(_7805_),
    .Y(_7858_)
);

NAND2X1 _20689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf2),
    .B(breg_27_bF$buf5),
    .Y(_10713_)
);

OAI21X1 _20269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10247_),
    .B(_10248_),
    .C(_10210_),
    .Y(_10253_)
);

NAND3X1 _16817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6464_),
    .B(_6451_),
    .C(_6454_),
    .Y(_6468_)
);

INVX8 _11952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .Y(_2825_)
);

NAND3X1 _21630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11741_),
    .B(_11742_),
    .C(_11743_),
    .Y(_11744_)
);

AOI21X1 _21210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11284_),
    .B(_11276_),
    .C(_11012_),
    .Y(_11285_)
);

AOI21X1 _19289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9151_),
    .B(_9155_),
    .C(_9164_),
    .Y(_9179_)
);

FILL SFILL54120x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9477_),
    .B(_9521_),
    .Y(_11428_)
);

OAI21X1 _12317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6802_),
    .B(_6812_),
    .C(_6791_),
    .Y(_6823_)
);

XNOR2X1 _22835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1137_),
    .Y(_1156_)
);

AOI21X1 _22415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_696_),
    .C(_495_),
    .Y(_697_)
);

OAI21X1 _16990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf3),
    .B(_4541__bF$buf3),
    .C(_6651_),
    .Y(_6657_)
);

AOI21X1 _16570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6180_),
    .B(_6185_),
    .C(_6164_),
    .Y(_6197_)
);

NAND3X1 _16150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5352_),
    .B(_5732_),
    .C(_5736_),
    .Y(_5737_)
);

FILL SFILL18680x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _17775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7517_),
    .B(_7518_),
    .Y(_7519_)
);

NAND3X1 _17355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7055_),
    .B(_7044_),
    .C(_7049_),
    .Y(_7059_)
);

OAI21X1 _12490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6220_),
    .B(_7338_),
    .C(_7448_),
    .Y(_8720_)
);

INVX8 _12070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf5),
    .Y(_4116_)
);

NAND3X1 _20901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10940_),
    .B(_10932_),
    .C(_10938_),
    .Y(_10947_)
);

OAI21X1 _13695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2930_),
    .B(_3048_),
    .C(_2919_),
    .Y(_3049_)
);

NOR2X1 _13275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2585_),
    .B(_2588_),
    .Y(_2589_)
);

NOR2X1 _23793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2165_),
    .Y(_2199_)
);

INVX1 _23373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .Y(_1743_)
);

NOR2X1 _19921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9868_),
    .B(_9871_),
    .Y(_9873_)
);

OAI21X1 _19501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .B(_9409_),
    .C(_9401_),
    .Y(_9412_)
);

FILL SFILL69240x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5393_),
    .B(_5397_),
    .C(_5378_),
    .Y(_5399_)
);

AOI21X1 _15421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4359_),
    .B(_4612_),
    .C(_4938_),
    .Y(_4940_)
);

XNOR2X1 _15001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4452_),
    .B(_4476_),
    .Y(_4479_)
);

FILL SFILL34040x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10502_),
    .B(_10503_),
    .Y(_10504_)
);

NAND2X1 _20078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9704_),
    .B(_9711_),
    .Y(_10043_)
);

OAI21X1 _16626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6252_),
    .B(_6254_),
    .C(_6255_),
    .Y(_6259_)
);

AOI21X1 _16206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5790_),
    .B(_5791_),
    .C(_5783_),
    .Y(_5799_)
);

AOI21X1 _19098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8952_),
    .B(_8958_),
    .C(_8936_),
    .Y(_8969_)
);

FILL SFILL69160x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _12966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_2012_),
    .Y(_2023_)
);

AOI21X1 _12546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9312_),
    .B(_9323_),
    .C(_9247_),
    .Y(_9334_)
);

FILL SFILL59240x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4708_),
    .B(_4719_),
    .C(_3865_),
    .Y(_4730_)
);

OAI21X1 _22644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_890_),
    .B(_886_),
    .C(_901_),
    .Y(_947_)
);

OAI21X1 _22224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_476_),
    .C(_479_),
    .Y(_487_)
);

FILL SFILL24040x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2256_),
    .B(_2235_),
    .Y(_2257_)
);

INVX1 _23429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .Y(_1803_)
);

NAND2X1 _23009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_868_),
    .B(_1213_),
    .Y(_1345_)
);

NAND3X1 _17584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7274_),
    .B(_7308_),
    .C(_7302_),
    .Y(_7309_)
);

NAND2X1 _17164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_25_bF$buf3),
    .Y(_6849_)
);

FILL SFILL28760x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10733_),
    .B(_10732_),
    .C(_10731_),
    .Y(_10736_)
);

XNOR2X1 _18789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8606_),
    .B(_8603_),
    .Y(_8630_)
);

NAND3X1 _18369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8156_),
    .B(_8160_),
    .C(_8163_),
    .Y(_8170_)
);

AOI22X1 _13084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_12_bF$buf4),
    .C(areg_2_bF$buf4),
    .D(breg_13_bF$buf3),
    .Y(_2380_)
);

NAND3X1 _23182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1525_),
    .C(_1520_),
    .Y(_1535_)
);

NOR2X1 _19730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9655_),
    .B(_9656_),
    .Y(_9662_)
);

OAI21X1 _19310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9200_),
    .B(_9201_),
    .C(_9141_),
    .Y(_9202_)
);

OAI21X1 _21915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_145_),
    .B(_143_),
    .C(_148_),
    .Y(_149_)
);

FILL SFILL33960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3698_),
    .B(_3697_),
    .C(_3696_),
    .Y(_3699_)
);

FILL SFILL18760x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5183_),
    .B(_5184_),
    .Y(_5189_)
);

NOR2X1 _15230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4450_),
    .B(_4451_),
    .Y(_4729_)
);

FILL SFILL18680x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6356_),
    .B(_6362_),
    .C(_6219_),
    .Y(_6510_)
);

NAND2X1 _16435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_28_bF$buf4),
    .Y(_6049_)
);

NAND3X1 _16015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5572_),
    .B(_5577_),
    .C(_5580_),
    .Y(_5590_)
);

INVX1 _11990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3231_),
    .Y(_3241_)
);

FILL SFILL54200x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11789_),
    .B(_11833_),
    .Y(_11844_)
);

OAI21X1 _12355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf3),
    .B(_7217__bF$buf0),
    .C(_7228_),
    .Y(_7239_)
);

NAND2X1 _22873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1191_),
    .B(_1196_),
    .Y(_1198_)
);

NOR2X1 _22453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf1),
    .B(_6815__bF$buf4),
    .Y(_738_)
);

NOR3X1 _22033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_277_),
    .B(_272_),
    .C(_276_),
    .Y(_278_)
);

FILL SFILL69320x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _23658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1937_),
    .B(_1946_),
    .C(_2048_),
    .Y(_2052_)
);

NAND2X1 _23238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1594_),
    .Y(_1595_)
);

FILL SFILL69240x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4107_),
    .B(_4114_),
    .C(_4103_),
    .Y(_4391_)
);

NAND2X1 _14501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .B(_3391_),
    .Y(_3932_)
);

OAI21X1 _17393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_7100__bF$buf3),
    .C(_7096_),
    .Y(_7101_)
);

OAI21X1 _15706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5095_),
    .B(_5090_),
    .C(_5097_),
    .Y(_5251_)
);

AOI21X1 _18598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8419_),
    .B(_8420_),
    .C(_8418_),
    .Y(_8421_)
);

AND2X2 _18178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_29_bF$buf0),
    .Y(_7961_)
);

FILL SFILL19160x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11846_),
    .B(_11847_),
    .C(_11600_),
    .Y(_11848_)
);

AOI21X1 _21304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11381_),
    .B(_11380_),
    .C(_11379_),
    .Y(_11388_)
);

NAND3X1 _14098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3488_),
    .C(_3489_),
    .Y(_3490_)
);

FILL SFILL3800x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3800x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3400x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1089_),
    .B(_1253_),
    .C(_1092_),
    .Y(_1258_)
);

AOI21X1 _22509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_631_),
    .C(_619_),
    .Y(_799_)
);

FILL FILL74200x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_6300__bF$buf1),
    .C(_6296_),
    .Y(_6301_)
);

INVX2 _16244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5840_),
    .Y(_5841_)
);

FILL SFILL28760x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7618_),
    .B(_7620_),
    .C(_7619_),
    .Y(_7621_)
);

NAND3X1 _17449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7159_),
    .B(_7161_),
    .C(_7160_),
    .Y(_7162_)
);

INVX2 _17029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6700_),
    .Y(_6701_)
);

NAND3X1 _12584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9718_),
    .B(_9729_),
    .C(_9740_),
    .Y(_9751_)
);

NAND2X1 _12164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_8_bF$buf1),
    .Y(_5146_)
);

NAND2X1 _22682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf0),
    .B(breg_24_bF$buf2),
    .Y(_989_)
);

NAND3X1 _22262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_506_),
    .B(_528_),
    .C(_526_),
    .Y(_529_)
);

NAND3X1 _18810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8652_),
    .B(_8646_),
    .C(_8649_),
    .Y(_8653_)
);

FILL SFILL33960x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_17_bF$buf2),
    .Y(_3152_)
);

OAI21X1 _13369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2691_),
    .B(_2685_),
    .C(_2651_),
    .Y(_2692_)
);

BUFX2 _23887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[5]),
    .Y(y[5])
);

OAI21X1 _23467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1844_),
    .B(_1841_),
    .C(_1727_),
    .Y(_1845_)
);

AOI21X1 _23047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1386_),
    .B(_1379_),
    .C(_1264_),
    .Y(_1387_)
);

OAI21X1 _14730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4179_),
    .B(_4180_),
    .C(_4176_),
    .Y(_4181_)
);

NAND3X1 _14310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3631_),
    .B(_3633_),
    .C(_3627_),
    .Y(_3722_)
);

FILL SFILL33800x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74280x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5169_),
    .B(_5171_),
    .C(_5167_),
    .Y(_5502_)
);

OAI21X1 _15515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4737_),
    .B(_4735_),
    .C(_4726_),
    .Y(_5041_)
);

NAND3X1 _21953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_82_),
    .B(_86_),
    .C(_88_),
    .Y(_191_)
);

AOI21X1 _21533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11633_),
    .B(_11634_),
    .C(_11608_),
    .Y(_11639_)
);

OAI21X1 _21113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_6686__bF$buf2),
    .C(_11172_),
    .Y(_11179_)
);

FILL SFILL69320x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_1043_),
    .Y(_1050_)
);

AOI21X1 _22318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .B(_578_),
    .C(_543_),
    .Y(_590_)
);

AND2X2 _16893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_16_bF$buf4),
    .Y(_6552_)
);

AOI21X1 _16473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6083_),
    .B(_6084_),
    .C(_6082_),
    .Y(_6091_)
);

AOI21X1 _16053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5620_),
    .C(_5367_),
    .Y(_5632_)
);

AOI21X1 _17678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7395_),
    .B(_7400_),
    .C(_7380_),
    .Y(_7412_)
);

XNOR2X1 _17258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6930_),
    .B(_6925_),
    .Y(_6952_)
);

INVX1 _12393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7645_),
    .Y(_7656_)
);

OAI21X1 _22491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_776_),
    .C(_775_),
    .Y(_780_)
);

NAND3X1 _22071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_313_),
    .C(_318_),
    .Y(_320_)
);

NOR2X1 _20804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10826_),
    .B(_10823_),
    .Y(_10840_)
);

OAI21X1 _13598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2939_),
    .B(_2938_),
    .C(_2793_),
    .Y(_2943_)
);

NAND3X1 _13178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_2469_),
    .C(_2467_),
    .Y(_2483_)
);

NAND2X1 _23696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2092_),
    .B(_2083_),
    .Y(_2094_)
);

NAND3X1 _23276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_1633_),
    .C(_1632_),
    .Y(_1637_)
);

FILL SFILL3800x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf2),
    .B(breg_20_bF$buf1),
    .Y(_9766_)
);

NAND3X1 _19404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9292_),
    .B(_9284_),
    .C(_9296_),
    .Y(_9305_)
);

FILL FILL74200x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5288_),
    .B(_5290_),
    .C(_4965_),
    .Y(_5293_)
);

OAI21X1 _15324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4830_),
    .B(_4532_),
    .C(_4832_),
    .Y(_4833_)
);

AND2X2 _16949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_20_bF$buf2),
    .Y(_6613_)
);

NAND3X1 _16529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6146_),
    .B(_6148_),
    .C(_6147_),
    .Y(_6152_)
);

OAI21X1 _16109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf0),
    .B(_5318_),
    .C(_5679_),
    .Y(_5692_)
);

NAND2X1 _21762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11691_),
    .B(_11696_),
    .Y(_11889_)
);

NOR3X1 _21342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11212_),
    .B(_11215_),
    .C(_11214_),
    .Y(_11430_)
);

FILL SFILL13560x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11679_),
    .B(_911_),
    .C(_954_),
    .Y(_965_)
);

NAND3X1 _12449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7185_),
    .B(_8205_),
    .C(_8216_),
    .Y(_8271_)
);

OAI21X1 _22967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5315__bF$buf2),
    .B(_6686__bF$buf0),
    .C(_1139_),
    .Y(_1300_)
);

OAI21X1 _12029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3569_),
    .B(_3635_),
    .C(_3657_),
    .Y(_3668_)
);

NAND2X1 _22547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_22_bF$buf4),
    .B(areg_26_bF$buf0),
    .Y(_841_)
);

OAI21X1 _22127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_105_),
    .B(_378_),
    .C(_380_),
    .Y(_381_)
);

OAI21X1 _13810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3173_),
    .B(_3174_),
    .C(_3139_),
    .Y(_3175_)
);

NAND3X1 _16282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5879_),
    .B(_5880_),
    .C(_5882_),
    .Y(_5883_)
);

INVX1 _17487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6778_),
    .Y(_7203_)
);

NAND3X1 _17067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6603_),
    .B(_6645_),
    .C(_6646_),
    .Y(_6743_)
);

NOR3X1 _20613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10287_),
    .B(_10289_),
    .C(_10284_),
    .Y(_10631_)
);

FILL SFILL13640x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _23085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .Y(_1428_)
);

NAND3X1 _19633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9550_),
    .B(_9551_),
    .C(_9552_),
    .Y(_9557_)
);

NAND2X1 _19213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9089_),
    .B(_9094_),
    .Y(_9095_)
);

NAND3X1 _21818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_39_),
    .C(_41_),
    .Y(_42_)
);

FILL SFILL74280x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5543_),
    .Y(_5544_)
);

AOI21X1 _15553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5032_),
    .B(_5031_),
    .C(_5019_),
    .Y(_5083_)
);

FILL SFILL13960x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4622_),
    .B(_4623_),
    .C(_4620_),
    .Y(_4624_)
);

NAND3X1 _16758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6043_),
    .B(_6399_),
    .C(_6403_),
    .Y(_6404_)
);

NAND2X1 _16338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5938_),
    .B(_5558_),
    .Y(_5944_)
);

FILL SFILL43720x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11882_),
    .B(_224_),
    .C(_218_),
    .Y(_233_)
);

AOI21X1 _21571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11673_),
    .B(_11674_),
    .C(_11672_),
    .Y(_11680_)
);

NAND2X1 _21151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10882_),
    .B(_10889_),
    .Y(_11221_)
);

NOR2X1 _12678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10759_),
    .B(_10770_),
    .Y(_10781_)
);

XNOR2X1 _12258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6165_),
    .B(_6132_),
    .Y(_6176_)
);

NAND3X1 _22776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_944_),
    .B(_1090_),
    .C(_1091_),
    .Y(_1092_)
);

OAI21X1 _22356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_6686__bF$buf0),
    .C(_624_),
    .Y(_632_)
);

AOI21X1 _18904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8751_),
    .B(_8752_),
    .C(_8745_),
    .Y(_8757_)
);

NAND2X1 _16091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5325_),
    .B(_5331_),
    .Y(_5673_)
);

AOI21X1 _14824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4266_),
    .B(_4272_),
    .C(_4233_),
    .Y(_4285_)
);

NAND3X1 _14404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3816_),
    .B(_3819_),
    .C(_3824_),
    .Y(_3825_)
);

AOI21X1 _17296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6992_),
    .B(_6993_),
    .C(_6985_),
    .Y(_6994_)
);

OAI21X1 _15609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5138_),
    .B(_5139_),
    .C(_5140_),
    .Y(_5144_)
);

NAND3X1 _20842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10850_),
    .B(_10876_),
    .C(_10881_),
    .Y(_10882_)
);

OAI21X1 _20422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10412_),
    .B(_10411_),
    .C(_10409_),
    .Y(_10421_)
);

AOI21X1 _20002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9954_),
    .B(_9960_),
    .C(_9642_),
    .Y(_9961_)
);

NAND3X1 _19862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9807_),
    .B(_9800_),
    .C(_9803_),
    .Y(_9808_)
);

NAND3X1 _19442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9343_),
    .B(_9344_),
    .C(_9346_),
    .Y(_9347_)
);

OAI21X1 _19022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8885_),
    .B(_8480_),
    .C(_8855_),
    .Y(_8886_)
);

INVX8 _11949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf4),
    .Y(_2792_)
);

AOI21X1 _21627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11455_),
    .B(_11457_),
    .C(_11449_),
    .Y(_11741_)
);

AOI21X1 _21207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11254_),
    .B(_11258_),
    .C(_11271_),
    .Y(_11282_)
);

NAND3X1 _15782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5329_),
    .B(_5317_),
    .C(_5322_),
    .Y(_5334_)
);

OAI21X1 _15362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4869_),
    .B(_4868_),
    .C(_4854_),
    .Y(_4875_)
);

FILL SFILL8680x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_22_bF$buf4),
    .Y(_6654_)
);

NAND3X1 _16567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6184_),
    .B(_6172_),
    .C(_6175_),
    .Y(_6194_)
);

AOI21X1 _16147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5718_),
    .B(_5724_),
    .C(_5669_),
    .Y(_5734_)
);

OR2X2 _21380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11470_),
    .B(_11465_),
    .Y(_11471_)
);

FILL SFILL44120x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7459_),
    .B(_7470_),
    .C(_7942_),
    .Y(_8687_)
);

NAND2X1 _12067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg_7_bF$buf5),
    .Y(_4083_)
);

NAND3X1 _22585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_828_),
    .C(_832_),
    .Y(_883_)
);

NAND2X1 _22165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .B(_157_),
    .Y(_423_)
);

NOR3X1 _18713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8530_),
    .B(_8534_),
    .C(_8535_),
    .Y(_8547_)
);

FILL SFILL74280x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_7520__bF$buf3),
    .C(_9868_),
    .Y(_9869_)
);

NAND2X1 _14633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_20_bF$buf2),
    .Y(_4075_)
);

NOR2X1 _14213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(_3602_),
    .Y(_3616_)
);

FILL SFILL74200x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5380_),
    .B(_5390_),
    .C(_5391_),
    .Y(_5395_)
);

NAND3X1 _15418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4933_),
    .B(_4934_),
    .C(_4935_),
    .Y(_4936_)
);

OAI21X1 _20651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10668_),
    .B(_10663_),
    .C(_10670_),
    .Y(_10672_)
);

NAND2X1 _20231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf0),
    .B(areg_24_bF$buf2),
    .Y(_10211_)
);

OAI21X1 _19671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9591_),
    .B(_9597_),
    .C(_9276_),
    .Y(_9599_)
);

AOI21X1 _19251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9131_),
    .B(_9132_),
    .C(_9133_),
    .Y(_9138_)
);

AOI21X1 _21856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_74_),
    .C(_24_),
    .Y(_84_)
);

OR2X2 _21436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10565_),
    .B(_11237_),
    .Y(_11533_)
);

NAND2X1 _21016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf3),
    .B(breg_22_bF$buf2),
    .Y(_11072_)
);

FILL SFILL33800x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64200x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf3),
    .B(_2669__bF$buf2),
    .C(_5112_),
    .Y(_5125_)
);

NOR2X1 _15171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4663_),
    .B(_4662_),
    .Y(_4665_)
);

OAI21X1 _13904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3277_),
    .B(_3276_),
    .C(_3271_),
    .Y(_3278_)
);

INVX1 _16796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6444_),
    .Y(_6445_)
);

AOI21X1 _16376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5979_),
    .B(_5980_),
    .C(_5978_),
    .Y(_5985_)
);

FILL SFILL58920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_6582__bF$buf0),
    .C(_5179_),
    .Y(_6593_)
);

AOI21X1 _22394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_671_),
    .C(_672_),
    .Y(_673_)
);

OAI21X1 _18942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8384_),
    .B(_8396_),
    .C(_8792_),
    .Y(_8799_)
);

AND2X2 _18522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_27_bF$buf2),
    .Y(_8339_)
);

NAND2X1 _18102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7872_),
    .B(_7877_),
    .Y(_7878_)
);

NOR3X1 _20707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10718_),
    .B(_10703_),
    .C(_10724_),
    .Y(_10733_)
);

INVX1 _23599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1983_),
    .Y(_1988_)
);

OAI21X1 _23179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1530_),
    .B(_1526_),
    .C(_1404_),
    .Y(_1531_)
);

NAND3X1 _19727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9654_),
    .B(_9658_),
    .C(_9657_),
    .Y(_9659_)
);

NAND3X1 _19307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9194_),
    .B(_9195_),
    .C(_9191_),
    .Y(_9199_)
);

NAND3X1 _14862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4058_),
    .B(_4326_),
    .C(_4321_),
    .Y(_4327_)
);

OAI21X1 _14442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3638_),
    .B(_3732_),
    .C(_3725_),
    .Y(_3867_)
);

NAND2X1 _14022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_19_bF$buf2),
    .Y(_3407_)
);

OAI21X1 _15647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_4551__bF$buf4),
    .C(_5183_),
    .Y(_5186_)
);

NAND3X1 _15227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4718_),
    .B(_4722_),
    .C(_4725_),
    .Y(_4726_)
);

OAI21X1 _20880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf3),
    .B(_8759_),
    .C(_10919_),
    .Y(_10923_)
);

NAND2X1 _20460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10173_),
    .B(_10181_),
    .Y(_10462_)
);

INVX1 _20040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10000_),
    .Y(_10001_)
);

FILL SFILL48840x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9202_),
    .B(_9199_),
    .C(_9096_),
    .Y(_9388_)
);

NOR3X1 _19060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8924_),
    .B(_8925_),
    .C(_8926_),
    .Y(_8927_)
);

XNOR2X1 _11987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3198_),
    .B(_2683_),
    .Y(_3209_)
);

AOI21X1 _21665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11763_),
    .B(_11766_),
    .C(_11769_),
    .Y(_11783_)
);

NAND2X1 _21245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11118_),
    .B(_11125_),
    .Y(_11323_)
);

OAI21X1 _13713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3064_),
    .B(_3063_),
    .C(_3068_),
    .Y(_3069_)
);

NAND2X1 _23811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2183_),
    .Y(_2218_)
);

FILL SFILL38840x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5767_),
    .B(_5753_),
    .C(_5772_),
    .Y(_5776_)
);

FILL SFILL43800x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4380_),
    .B(_4384_),
    .C(_4366_),
    .Y(_4387_)
);

FILL SFILL3480x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8583_),
    .B(_8584_),
    .C(_8582_),
    .Y(_8589_)
);

NOR2X1 _18331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8126_),
    .B(_8127_),
    .Y(_8129_)
);

NAND3X1 _20936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10694_),
    .B(_10980_),
    .C(_10981_),
    .Y(_10985_)
);

NOR3X1 _20516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10516_),
    .B(_10520_),
    .C(_10515_),
    .Y(_10524_)
);

FILL SFILL33800x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_9153_),
    .C(_9909_),
    .Y(_9910_)
);

FILL SFILL64200x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9442_),
    .B(_9449_),
    .C(_9427_),
    .Y(_9450_)
);

NAND3X1 _19116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8988_),
    .B(_8986_),
    .C(_8987_),
    .Y(_8989_)
);

OAI21X1 _14671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf0),
    .B(_2362__bF$buf5),
    .C(_4101_),
    .Y(_4117_)
);

INVX1 _14251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3392_),
    .Y(_3658_)
);

AOI21X1 _15876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5043_),
    .B(_5065_),
    .C(_5068_),
    .Y(_5437_)
);

NOR2X1 _15456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4975_),
    .B(_4974_),
    .Y(_4976_)
);

AOI21X1 _15036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4506_),
    .B(_4505_),
    .C(_4502_),
    .Y(_4517_)
);

FILL SFILL18840x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _21894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_125_),
    .Y(_126_)
);

NOR3X1 _21474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11551_),
    .B(_11557_),
    .C(_11559_),
    .Y(_11575_)
);

NAND3X1 _21054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11104_),
    .B(_11097_),
    .C(_11102_),
    .Y(_11114_)
);

NAND3X1 _17602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7325_),
    .B(_7328_),
    .C(_7321_),
    .Y(_7329_)
);

FILL SFILL38840x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_984_),
    .C(_983_),
    .Y(_985_)
);

OAI21X1 _22259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_524_),
    .B(_520_),
    .C(_507_),
    .Y(_525_)
);

NOR2X1 _18807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8243_),
    .B(_8286_),
    .Y(_8650_)
);

XNOR2X1 _13942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3319_),
    .B(_3313_),
    .Y(_3320_)
);

NOR2X1 _13522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2844_),
    .B(_2846_),
    .Y(_2860_)
);

XNOR2X1 _13102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2395_),
    .B(_2399_),
    .Y(_2400_)
);

NAND2X1 _23620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_27_bF$buf1),
    .B(breg_29_bF$buf2),
    .Y(_2011_)
);

INVX2 _23200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .Y(_1553_)
);

FILL SFILL69080x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48920x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_549__bF$buf3),
    .C(_4166_),
    .Y(_4178_)
);

NAND3X1 _14307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3717_),
    .B(_3718_),
    .C(_3716_),
    .Y(_3719_)
);

OAI21X1 _17199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6884_),
    .B(_6883_),
    .C(_6886_),
    .Y(_6887_)
);

FILL SFILL13720x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8587_),
    .B(_8594_),
    .C(_8592_),
    .Y(_8840_)
);

OAI21X1 _18560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7971_),
    .C(_8379_),
    .Y(_8380_)
);

NAND3X1 _18140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7918_),
    .B(_7916_),
    .C(_7917_),
    .Y(_7919_)
);

AOI21X1 _20745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10768_),
    .B(_10769_),
    .C(_10767_),
    .Y(_10775_)
);

AOI21X1 _20325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10304_),
    .B(_10298_),
    .C(_9996_),
    .Y(_10315_)
);

NAND3X1 _19765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9698_),
    .B(_9700_),
    .C(_9699_),
    .Y(_9701_)
);

NAND3X1 _19345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8887_),
    .B(_9234_),
    .C(_9235_),
    .Y(_9241_)
);

AND2X2 _14480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3628_),
    .B(_3622_),
    .Y(_3908_)
);

AOI21X1 _14060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3430_),
    .B(_3434_),
    .C(_3358_),
    .Y(_3448_)
);

FILL SFILL38920x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5224_),
    .B(_5226_),
    .C(_5225_),
    .Y(_5227_)
);

OAI21X1 _15265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4587_),
    .B(_4767_),
    .C(_4578_),
    .Y(_4768_)
);

OAI21X1 _21283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11360_),
    .B(_11359_),
    .C(_11358_),
    .Y(_11365_)
);

FILL SFILL28920x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7559_),
    .B(_7565_),
    .C(_7568_),
    .Y(_7581_)
);

AOI21X1 _17411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6696_),
    .B(_6701_),
    .C(_6706_),
    .Y(_7121_)
);

FILL SFILL28840x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _22488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf2),
    .B(breg_25_bF$buf1),
    .C(areg_23_bF$buf0),
    .D(breg_24_bF$buf2),
    .Y(_776_)
);

OAI21X1 _22068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781__bF$buf0),
    .B(_4541__bF$buf4),
    .C(_40_),
    .Y(_316_)
);

NAND3X1 _18616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8422_),
    .B(_8428_),
    .C(_8185_),
    .Y(_8441_)
);

NAND2X1 _13751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_14_bF$buf4),
    .Y(_3111_)
);

NAND2X1 _13331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2645_),
    .B(_2649_),
    .Y(_2651_)
);

OAI21X1 _14956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4425_),
    .B(_4424_),
    .C(_4389_),
    .Y(_4429_)
);

AOI21X1 _14536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3684_),
    .B(_3687_),
    .C(_3681_),
    .Y(_3970_)
);

NAND3X1 _14116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3501_),
    .B(_3504_),
    .C(_3508_),
    .Y(_3509_)
);

FILL SFILL18680x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf2),
    .B(breg_27_bF$buf5),
    .Y(_11026_)
);

NAND2X1 _20554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10219_),
    .B(_10565_),
    .Y(_10566_)
);

NAND3X1 _20134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10100_),
    .B(_10095_),
    .C(_10091_),
    .Y(_10105_)
);

OAI21X1 _19994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9930_),
    .B(_9936_),
    .C(_9940_),
    .Y(_9952_)
);

AND2X2 _19574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf0),
    .B(areg_26_bF$buf3),
    .Y(_9492_)
);

AOI21X1 _19154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9021_),
    .B(_9020_),
    .C(_9017_),
    .Y(_9031_)
);

NAND2X1 _21759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11703_),
    .B(_11708_),
    .Y(_11885_)
);

NAND3X1 _21339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11423_),
    .B(_11425_),
    .C(_11419_),
    .Y(_11426_)
);

AOI21X1 _12602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9729_),
    .B(_9740_),
    .C(_9718_),
    .Y(_9948_)
);

OAI21X1 _22700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .B(_1006_),
    .C(_1005_),
    .Y(_1008_)
);

AOI21X1 _15494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .B(_4692_),
    .C(_4690_),
    .Y(_5018_)
);

XNOR2X1 _15074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4534_),
    .B(_4529_),
    .Y(_4559_)
);

FILL SFILL69080x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3168_),
    .B(_3167_),
    .C(_3166_),
    .Y(_3172_)
);

BUFX2 _23905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[23]),
    .Y(y[23])
);

AOI21X1 _16699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6328_),
    .C(_6306_),
    .Y(_6339_)
);

AND2X2 _16279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5491_),
    .B(_5485_),
    .Y(_5879_)
);

NOR2X1 _21092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10838_),
    .B(_11155_),
    .Y(_11156_)
);

NAND3X1 _17640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7367_),
    .B(_7368_),
    .C(_7369_),
    .Y(_7370_)
);

AOI21X1 _17220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6894_),
    .B(_6901_),
    .C(_6844_),
    .Y(_6910_)
);

NAND2X1 _12199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_6_bF$buf2),
    .Y(_5530_)
);

NAND3X1 _22297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_544_),
    .B(_559_),
    .C(_566_),
    .Y(_567_)
);

NAND2X1 _18845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8686_),
    .B(_8691_),
    .Y(_8692_)
);

NAND3X1 _18425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8228_),
    .B(_8231_),
    .C(_8230_),
    .Y(_8232_)
);

NOR3X1 _18005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7423_),
    .B(_7424_),
    .C(_7427_),
    .Y(_7771_)
);

FILL SFILL59080x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2845_),
    .B(_3359_),
    .C(_3106_),
    .Y(_3360_)
);

AOI21X1 _13560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2894_),
    .B(_2899_),
    .C(_2870_),
    .Y(_2900_)
);

NAND3X1 _13140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .B(_2425_),
    .C(_2434_),
    .Y(_2441_)
);

FILL SFILL38920x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59320x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_3673_),
    .Y(_4220_)
);

NAND3X1 _14345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3757_),
    .B(_3760_),
    .C(_3755_),
    .Y(_3761_)
);

DFFPOSX1 _24023_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[13]),
    .CLK(clk_bF$buf8),
    .D(a[13])
);

FILL SFILL3560x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _20783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10816_),
    .Y(_10817_)
);

OAI21X1 _20363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10017_),
    .B(_10007_),
    .C(_10011_),
    .Y(_10356_)
);

FILL SFILL28920x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6548_),
    .B(_6564_),
    .C(_6570_),
    .Y(_6572_)
);

NOR2X1 _19383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf0),
    .B(_6815__bF$buf2),
    .Y(_9282_)
);

OAI22X1 _21988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_225_),
    .B(_228_),
    .C(_11854_),
    .D(_11880_),
    .Y(_229_)
);

AOI21X1 _21568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11462_),
    .B(_11463_),
    .C(_11446_),
    .Y(_11676_)
);

OAI21X1 _21148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11216_),
    .B(_10945_),
    .C(_10939_),
    .Y(_11217_)
);

INVX8 _12831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf0),
    .Y(_549_)
);

AOI21X1 _12411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7766_),
    .B(_7733_),
    .C(_7656_),
    .Y(_7854_)
);

FILL SFILL18920x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2961_),
    .B(_2962_),
    .C(_2960_),
    .Y(_2963_)
);

AOI21X1 _23714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1983_),
    .B(_2111_),
    .C(_2112_),
    .Y(_2113_)
);

NOR2X1 _16088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf2),
    .B(_5668__bF$buf2),
    .Y(_5669_)
);

FILL SFILL49080x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8185_),
    .B(_8481_),
    .C(_8433_),
    .Y(_8482_)
);

NAND3X1 _18234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8016_),
    .B(_8017_),
    .C(_8015_),
    .Y(_8022_)
);

NOR3X1 _20839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10871_),
    .B(_10874_),
    .C(_10870_),
    .Y(_10878_)
);

NAND3X1 _20419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10394_),
    .B(_10410_),
    .C(_10416_),
    .Y(_10417_)
);

NOR2X1 _19859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9446_),
    .B(_9485_),
    .Y(_9804_)
);

INVX1 _19439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9321_),
    .Y(_9343_)
);

OAI21X1 _19019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8515_),
    .B(_8485_),
    .C(_8523_),
    .Y(_8882_)
);

OAI21X1 _14994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf2),
    .B(_549__bF$buf3),
    .C(_4458_),
    .Y(_4470_)
);

OAI21X1 _14574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4004_),
    .B(_4011_),
    .C(_3867_),
    .Y(_4012_)
);

AOI21X1 _14154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3312_),
    .B(_3550_),
    .C(_3316_),
    .Y(_3551_)
);

OAI21X1 _15779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5326_),
    .B(_5327_),
    .C(_5329_),
    .Y(_5330_)
);

NAND3X1 _15359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4853_),
    .B(_4870_),
    .C(_4866_),
    .Y(_4871_)
);

FILL SFILL3720x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10607_),
    .B(_10602_),
    .Y(_10608_)
);

INVX1 _20172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10146_),
    .Y(_10147_)
);

NAND3X1 _16720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6361_),
    .B(_6360_),
    .C(_6359_),
    .Y(_6362_)
);

AOI21X1 _16300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5897_),
    .B(_5898_),
    .C(_5889_),
    .Y(_5902_)
);

NAND3X1 _19192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9066_),
    .B(_9067_),
    .C(_9068_),
    .Y(_9073_)
);

OAI21X1 _21797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_18_),
    .B(_14_),
    .C(_11891_),
    .Y(_19_)
);

NAND3X1 _21377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11462_),
    .B(_11446_),
    .C(_11463_),
    .Y(_11468_)
);

OAI21X1 _17925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7682_),
    .B(_7681_),
    .C(_7672_),
    .Y(_7683_)
);

AOI21X1 _17505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7170_),
    .B(_7176_),
    .C(_6921_),
    .Y(_7222_)
);

FILL SFILL59080x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10332_),
    .B(_10353_),
    .C(_10342_),
    .Y(_10364_)
);

OAI21X1 _12220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5749_),
    .B(_5705_),
    .C(_4204_),
    .Y(_5760_)
);

FILL SFILL43880x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2790_),
    .B(_2940_),
    .C(_3213_),
    .Y(_3214_)
);

NOR3X1 _13425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2737_),
    .C(_2735_),
    .Y(_2753_)
);

BUFX2 _23943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[61]),
    .Y(y[61])
);

XNOR2X1 _13005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2153_),
    .Y(_2300_)
);

NOR2X1 _23523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1812_),
    .B(_1904_),
    .Y(_1905_)
);

NAND2X1 _23103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf5),
    .B(areg_27_bF$buf4),
    .Y(_1448_)
);

NAND3X1 _18883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8733_),
    .B(_8730_),
    .C(_8732_),
    .Y(_8734_)
);

NAND3X1 _18463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8188_),
    .B(_8273_),
    .C(_8268_),
    .Y(_8274_)
);

NOR3X1 _18043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7792_),
    .B(_7808_),
    .C(_7807_),
    .Y(_7813_)
);

FILL SFILL18600x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10665_),
    .B(_10664_),
    .C(_10667_),
    .D(_10666_),
    .Y(_10668_)
);

OAI21X1 _20228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10206_),
    .B(_10207_),
    .C(_9920_),
    .Y(_10208_)
);

INVX8 _11911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(_2376_)
);

NAND3X1 _19668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9588_),
    .B(_9589_),
    .C(_9390_),
    .Y(_9595_)
);

NAND3X1 _19248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9133_),
    .B(_9131_),
    .C(_9132_),
    .Y(_9134_)
);

OAI21X1 _14383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3801_),
    .B(_3798_),
    .C(_3783_),
    .Y(_3802_)
);

DFFPOSX1 _24061_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[19]),
    .CLK(clk_bF$buf4),
    .D(b[19])
);

FILL SFILL54280x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5117_),
    .B(_5109_),
    .C(_5120_),
    .Y(_5121_)
);

OAI21X1 _15168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4068_),
    .B(_4364_),
    .C(_4660_),
    .Y(_4661_)
);

NAND2X1 _21186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11258_),
    .B(_11254_),
    .Y(_11259_)
);

AOI21X1 _17734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7456_),
    .B(_7463_),
    .C(_7442_),
    .Y(_7474_)
);

NAND2X1 _17314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7009_),
    .B(_7012_),
    .Y(_7013_)
);

FILL SFILL29080x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8738_),
    .B(_8737_),
    .C(_8695_),
    .Y(_8795_)
);

NAND2X1 _18519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_25_bF$buf4),
    .Y(_8335_)
);

INVX2 _13654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3003_),
    .Y(_3004_)
);

OAI21X1 _13234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2539_),
    .B(_2532_),
    .C(_2543_),
    .Y(_2544_)
);

NOR2X1 _23752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2154_),
    .Y(_2155_)
);

NAND2X1 _23332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1695_),
    .B(_1697_),
    .Y(_1698_)
);

AOI21X1 _14859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4318_),
    .B(_4319_),
    .C(_4317_),
    .Y(_4323_)
);

OAI21X1 _14439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3856_),
    .B(_3857_),
    .C(_3853_),
    .Y(_3863_)
);

FILL SFILL3720x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_3403_)
);

AND2X2 _15800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5348_),
    .B(_5352_),
    .Y(_5353_)
);

NAND3X1 _18692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8484_),
    .B(_8523_),
    .C(_8521_),
    .Y(_8524_)
);

OAI21X1 _18272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8062_),
    .B(_8064_),
    .C(_7657_),
    .Y(_8065_)
);

NAND2X1 _20877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10565_),
    .B(_10919_),
    .Y(_10920_)
);

NAND3X1 _20457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10457_),
    .B(_10458_),
    .C(_10456_),
    .Y(_10459_)
);

OAI21X1 _20037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9754_),
    .B(_9997_),
    .C(_9951_),
    .Y(_9998_)
);

FILL SFILL43960x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9524_),
    .B(_9845_),
    .C(_9517_),
    .Y(_9846_)
);

OAI21X1 _19477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .B(_9379_),
    .C(_9375_),
    .Y(_9385_)
);

AOI21X1 _19057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8487_),
    .B(_8512_),
    .C(_8509_),
    .Y(_8924_)
);

NAND2X1 _14192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3335_),
    .B(_3339_),
    .Y(_3593_)
);

FILL SFILL43880x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_8555_),
    .Y(_1586_)
);

NOR2X1 _12505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8874_),
    .B(_8863_),
    .Y(_8884_)
);

NAND3X1 _22603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_902_),
    .C(_899_),
    .Y(_903_)
);

AOI21X1 _15397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4892_),
    .B(_4898_),
    .C(_4812_),
    .Y(_4913_)
);

NAND3X1 _23808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2168_),
    .B(_2194_),
    .C(_2195_),
    .Y(_2214_)
);

BUFX2 BUFX2_insert220 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[23]),
    .Y(areg_23_bF$buf2)
);

BUFX2 BUFX2_insert221 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[23]),
    .Y(areg_23_bF$buf1)
);

BUFX2 BUFX2_insert222 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[23]),
    .Y(areg_23_bF$buf0)
);

BUFX2 BUFX2_insert223 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .Y(_3146__bF$buf3)
);

AOI21X1 _17963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7719_),
    .B(_7718_),
    .C(_7717_),
    .Y(_7725_)
);

BUFX2 BUFX2_insert224 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .Y(_3146__bF$buf2)
);

NOR3X1 _17543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7247_),
    .B(_7233_),
    .C(_7254_),
    .Y(_7264_)
);

BUFX2 BUFX2_insert225 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .Y(_3146__bF$buf1)
);

BUFX2 BUFX2_insert226 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146_),
    .Y(_3146__bF$buf0)
);

OAI21X1 _17123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6803_),
    .B(_6412_),
    .C(_6798_),
    .Y(_6804_)
);

BUFX2 BUFX2_insert227 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf4)
);

BUFX2 BUFX2_insert228 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf3)
);

BUFX2 BUFX2_insert229 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(areg_3_bF$buf2)
);

NAND3X1 _18748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8582_),
    .B(_8583_),
    .C(_8584_),
    .Y(_8585_)
);

NAND2X1 _18328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_26_bF$buf2),
    .Y(_8125_)
);

OAI21X1 _13883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_3253__bF$buf2),
    .C(_3254_),
    .Y(_3255_)
);

DFFPOSX1 _23981_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[35]),
    .CLK(clk_bF$buf3),
    .D(_0_[35])
);

NOR2X1 _13463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_2379_),
    .Y(_2795_)
);

INVX1 _13043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .Y(_2338_)
);

NAND3X1 _23561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1946_),
    .B(_1944_),
    .C(_1945_),
    .Y(_1948_)
);

NAND3X1 _23141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1483_),
    .C(_1488_),
    .Y(_1490_)
);

NAND3X1 _14668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_4112_),
    .C(_4108_),
    .Y(_4113_)
);

NAND3X1 _14248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3648_),
    .B(_3652_),
    .C(_3653_),
    .Y(_3654_)
);

FILL SFILL53960x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7849_),
    .B(_7850_),
    .C(_7853_),
    .Y(_7855_)
);

NAND2X1 _20686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10708_),
    .B(_10709_),
    .Y(_10710_)
);

FILL SFILL23800x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10245_),
    .B(_10249_),
    .C(_10209_),
    .Y(_10250_)
);

OAI21X1 _16814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6459_),
    .B(_6460_),
    .C(_6464_),
    .Y(_6465_)
);

OAI21X1 _19286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9172_),
    .B(_9166_),
    .C(_9175_),
    .Y(_9176_)
);

FILL SFILL29080x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10024_),
    .B(_11242_),
    .C(_11286_),
    .Y(_11395_)
);

NAND2X1 _12314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6286_),
    .B(_6330_),
    .Y(_6791_)
);

INVX1 _22832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .Y(_1153_)
);

NOR2X1 _22412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_500_),
    .B(_677_),
    .Y(_694_)
);

FILL SFILL29000x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3314_),
    .B(_3315_),
    .Y(_3316_)
);

NAND3X1 _13519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2852_),
    .B(_2855_),
    .C(_2848_),
    .Y(_2856_)
);

NOR2X1 _23617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(_1886_),
    .Y(_2008_)
);

INVX1 _17772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7515_),
    .Y(_7516_)
);

OAI21X1 _17352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7052_),
    .B(_7053_),
    .C(_7055_),
    .Y(_7056_)
);

FILL SFILL3880x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8802_),
    .B(_8824_),
    .C(_8692_),
    .Y(_8837_)
);

OAI21X1 _18557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8372_),
    .B(_8371_),
    .C(_8363_),
    .Y(_8377_)
);

NAND3X1 _18137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7911_),
    .B(_7912_),
    .C(_7910_),
    .Y(_7916_)
);

NAND3X1 _13692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3042_),
    .B(_3043_),
    .C(_3045_),
    .Y(_3046_)
);

OR2X2 _23790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2193_),
    .B(_2169_),
    .Y(_2195_)
);

INVX8 _13272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf4),
    .Y(_2586_)
);

AOI21X1 _23370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .B(_1722_),
    .C(_1664_),
    .Y(_1739_)
);

NAND2X1 _14897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_21_bF$buf1),
    .Y(_4364_)
);

OAI21X1 _14477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3662_),
    .B(_3664_),
    .C(_3654_),
    .Y(_3905_)
);

OAI21X1 _14057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3349_),
    .B(_3345_),
    .C(_3353_),
    .Y(_3445_)
);

INVX1 _20495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10500_),
    .Y(_10501_)
);

NAND3X1 _20075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10000_),
    .B(_10039_),
    .C(_10038_),
    .Y(_10040_)
);

NOR3X1 _16623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6254_),
    .B(_6255_),
    .C(_6252_),
    .Y(_6256_)
);

AND2X2 _16203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5419_),
    .B(_5795_),
    .Y(_5796_)
);

OAI21X1 _19095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8607_),
    .B(_8965_),
    .C(_8631_),
    .Y(_8966_)
);

NAND3X1 _17828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7575_),
    .B(_7576_),
    .C(_7438_),
    .Y(_7577_)
);

NOR2X1 _17408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6705_),
    .B(_7116_),
    .Y(_7117_)
);

OAI22X1 _12963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10748_),
    .B(_1979_),
    .C(_418_),
    .D(_451_),
    .Y(_1990_)
);

AOI21X1 _12543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7810_),
    .B(_7635_),
    .C(_7843_),
    .Y(_9301_)
);

NAND3X1 _12123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4642_),
    .B(_4072_),
    .C(_4686_),
    .Y(_4697_)
);

NAND2X1 _22641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_905_),
    .B(_912_),
    .Y(_944_)
);

XOR2X1 _22221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_239_),
    .B(_483_),
    .Y(_0_[45])
);

FILL SFILL59080x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf1),
    .B(_9104__bF$buf1),
    .C(_3103_),
    .Y(_3107_)
);

NAND2X1 _13328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2643_),
    .B(_2634_),
    .Y(_2647_)
);

XOR2X1 _23846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2242_),
    .B(_2254_),
    .Y(_2255_)
);

XNOR2X1 _23426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1799_),
    .B(_1788_),
    .Y(_1800_)
);

NAND3X1 _23006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(_1334_),
    .C(_1330_),
    .Y(_1342_)
);

NOR3X1 _17581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6947_),
    .B(_6945_),
    .C(_6940_),
    .Y(_7306_)
);

AOI21X1 _17161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6466_),
    .B(_6470_),
    .C(_6478_),
    .Y(_6846_)
);

OAI21X1 _18786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8626_),
    .B(_8625_),
    .C(_8611_),
    .Y(_8627_)
);

NAND3X1 _18366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8162_),
    .B(_8166_),
    .C(_8121_),
    .Y(_8167_)
);

OAI21X1 _13081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2323_),
    .B(_2375_),
    .C(_2317_),
    .Y(_2377_)
);

INVX1 _21912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11812_),
    .Y(_146_)
);

XOR2X1 _14286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .B(_3670_),
    .Y(_3696_)
);

FILL SFILL28840x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28760x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8680x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6491_),
    .B(_6496_),
    .C(_6497_),
    .Y(_6507_)
);

AOI21X1 _16432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5988_),
    .B(_5995_),
    .C(_5745_),
    .Y(_6046_)
);

OAI21X1 _16012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5529_),
    .B(_5533_),
    .C(_5535_),
    .Y(_5587_)
);

OAI21X1 _21089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10840_),
    .B(_10822_),
    .C(_10830_),
    .Y(_11152_)
);

AOI21X1 _17637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6941_),
    .B(_6943_),
    .C(_6936_),
    .Y(_7367_)
);

OAI21X1 _17217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6589_),
    .B(_6596_),
    .C(_6598_),
    .Y(_6907_)
);

OAI21X1 _12772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10123_),
    .B(_10233_),
    .C(_11800_),
    .Y(_11811_)
);

NAND3X1 _12352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg_10_bF$buf5),
    .C(_6055_),
    .Y(_7207_)
);

AOI22X1 _22870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_28_bF$buf2),
    .C(breg_22_bF$buf4),
    .D(areg_27_bF$buf5),
    .Y(_1194_)
);

INVX1 _22450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .Y(_734_)
);

OAI21X1 _22030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3146__bF$buf0),
    .B(_5668__bF$buf2),
    .C(_260_),
    .Y(_274_)
);

NAND2X1 _13977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3356_),
    .B(_3351_),
    .Y(_3357_)
);

NOR3X1 _13557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2892_),
    .B(_2876_),
    .C(_2891_),
    .Y(_2897_)
);

NOR2X1 _13137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2426_),
    .B(_2436_),
    .Y(_2438_)
);

AND2X2 _23655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1994_),
    .B(_2049_),
    .Y(_2050_)
);

INVX1 _23235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .Y(_1592_)
);

NAND2X1 _17390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_27_bF$buf1),
    .Y(_7097_)
);

OAI21X1 _15703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5246_),
    .B(_5247_),
    .C(_5243_),
    .Y(_5248_)
);

NAND2X1 _18595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8417_),
    .B(_8416_),
    .Y(_8418_)
);

FILL SFILL54040x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_27_bF$buf2),
    .Y(_7958_)
);

OAI21X1 _16908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf1),
    .B(_2669__bF$buf3),
    .C(_5842_),
    .Y(_6568_)
);

AOI21X1 _21721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11843_),
    .B(_11839_),
    .C(_11601_),
    .Y(_11845_)
);

AND2X2 _21301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11072_),
    .B(_11383_),
    .Y(_11385_)
);

NAND3X1 _14095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3480_),
    .B(_3486_),
    .C(_3243_),
    .Y(_3487_)
);

FILL SFILL8920x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_12_bF$buf1),
    .Y(_516_)
);

NAND3X1 _12408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7635_),
    .B(_7810_),
    .C(_7777_),
    .Y(_7821_)
);

OAI21X1 _22926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1240_),
    .B(_1243_),
    .C(_1246_),
    .Y(_1255_)
);

INVX2 _22506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .Y(_796_)
);

NAND2X1 _16661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .B(areg_25_bF$buf0),
    .Y(_6298_)
);

OAI21X1 _16241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5602_),
    .B(_5836_),
    .C(_5592_),
    .Y(_5838_)
);

INVX2 _17866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7221_),
    .Y(_7618_)
);

FILL SFILL74120x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7157_),
    .B(_7158_),
    .Y(_7159_)
);

AND2X2 _17026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_29_bF$buf4),
    .Y(_6698_)
);

NAND3X1 _12581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8249_),
    .B(_8260_),
    .C(_8271_),
    .Y(_9718_)
);

AOI21X1 _12161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4379_),
    .B(_4445_),
    .C(_5102_),
    .Y(_5113_)
);

FILL SFILL69160x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3145_),
    .B(_3148_),
    .C(_3141_),
    .Y(_3149_)
);

AOI21X1 _13366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .B(_2687_),
    .C(_2680_),
    .Y(_2689_)
);

BUFX2 _23884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[2]),
    .Y(y[2])
);

NOR3X1 _23464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1733_),
    .B(_1839_),
    .C(_1837_),
    .Y(_1842_)
);

AOI21X1 _23044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1364_),
    .B(_1368_),
    .C(_1371_),
    .Y(_1384_)
);

FILL SFILL64120x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5495_),
    .B(_5491_),
    .C(_5498_),
    .Y(_5499_)
);

OAI21X1 _15512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5029_),
    .B(_5024_),
    .C(_5018_),
    .Y(_5038_)
);

OAI21X1 _20589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10599_),
    .B(_10598_),
    .C(_10600_),
    .Y(_10604_)
);

NAND2X1 _20169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf5),
    .B(areg_22_bF$buf3),
    .Y(_10143_)
);

NAND2X1 _16717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6357_),
    .B(_6358_),
    .Y(_6359_)
);

NAND2X1 _21950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11826_),
    .B(_186_),
    .Y(_187_)
);

NAND3X1 _21530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11608_),
    .B(_11633_),
    .C(_11634_),
    .Y(_11635_)
);

OAI22X1 _21110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_6686__bF$buf2),
    .C(_2560__bF$buf3),
    .D(_6300__bF$buf3),
    .Y(_11175_)
);

AOI21X1 _19189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9067_),
    .B(_9068_),
    .C(_9066_),
    .Y(_9069_)
);

FILL SFILL54120x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10288_),
    .B(_10277_),
    .C(_10266_),
    .Y(_10332_)
);

AOI21X1 _12217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5661_),
    .B(_5672_),
    .C(_5683_),
    .Y(_5727_)
);

OAI21X1 _22735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_853_),
    .B(_1045_),
    .C(_1046_),
    .Y(_1047_)
);

NOR2X1 _22315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .B(_586_),
    .Y(_587_)
);

FILL FILL74040x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6163_),
    .B(_6547_),
    .C(_6172_),
    .Y(_6548_)
);

AOI21X1 _16470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5767_),
    .B(_5772_),
    .C(_5753_),
    .Y(_6086_)
);

OAI21X1 _16050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5363_),
    .B(_5362_),
    .C(_4996_),
    .Y(_5628_)
);

NAND3X1 _17675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7399_),
    .B(_7388_),
    .C(_7391_),
    .Y(_7409_)
);

OAI21X1 _17255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6939_),
    .B(_6936_),
    .C(_6934_),
    .Y(_6949_)
);

NOR2X1 _12390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7623_),
    .B(_7602_),
    .Y(_7624_)
);

NAND3X1 _20801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10829_),
    .B(_10832_),
    .C(_10830_),
    .Y(_10837_)
);

OAI21X1 _13595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2939_),
    .B(_2938_),
    .C(_2937_),
    .Y(_2940_)
);

AOI21X1 _13175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2474_),
    .B(_2479_),
    .C(_2448_),
    .Y(_2480_)
);

XOR2X1 _23693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2090_),
    .Y(_2091_)
);

AOI21X1 _23273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1633_),
    .B(_1632_),
    .C(_1552_),
    .Y(_1634_)
);

NOR2X1 _19821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9760_),
    .B(_9761_),
    .Y(_9763_)
);

NOR3X1 _19401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9300_),
    .B(_9298_),
    .C(_9299_),
    .Y(_9302_)
);

DFFPOSX1 _24058_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[16]),
    .CLK(clk_bF$buf4),
    .D(b[16])
);

AOI21X1 _15741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5277_),
    .B(_5270_),
    .C(_4967_),
    .Y(_5290_)
);

INVX1 _15321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4529_),
    .Y(_4830_)
);

OAI21X1 _20398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10050_),
    .B(_10045_),
    .C(_10053_),
    .Y(_10394_)
);

OAI21X1 _16946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6236_),
    .B(_6227_),
    .C(_6230_),
    .Y(_6610_)
);

AOI21X1 _16526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6148_),
    .B(_6147_),
    .C(_6146_),
    .Y(_6149_)
);

OAI22X1 _16106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5012_),
    .B(_5688_),
    .C(_5371_),
    .D(_5375_),
    .Y(_5689_)
);

NOR3X1 _12866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_878_),
    .B(_867_),
    .C(_889_),
    .Y(_932_)
);

AOI21X1 _12446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8183_),
    .B(_8227_),
    .C(_6955_),
    .Y(_8238_)
);

NAND2X1 _22964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1150_),
    .Y(_1297_)
);

NAND2X1 _12026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_6_bF$buf4),
    .Y(_3635_)
);

AOI21X1 _22544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_837_),
    .C(_835_),
    .Y(_838_)
);

NAND2X1 _22124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_27_bF$buf5),
    .Y(_378_)
);

XNOR2X1 _23749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2150_),
    .B(_2127_),
    .Y(_2151_)
);

OAI21X1 _23329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1597_),
    .B(_1600_),
    .C(_1593_),
    .Y(_1694_)
);

AOI21X1 _17484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7183_),
    .B(_7190_),
    .C(_6813_),
    .Y(_7200_)
);

AOI21X1 _17064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6721_),
    .B(_6727_),
    .C(_6677_),
    .Y(_6740_)
);

FILL SFILL28760x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10609_),
    .B(_10615_),
    .C(_10618_),
    .Y(_10627_)
);

OAI21X1 _18689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8519_),
    .B(_8515_),
    .C(_8485_),
    .Y(_8520_)
);

NAND3X1 _18269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7655_),
    .B(_8056_),
    .C(_8055_),
    .Y(_8061_)
);

XNOR2X1 _23082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1424_),
    .Y(_1425_)
);

AOI21X1 _19630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9551_),
    .B(_9552_),
    .C(_9550_),
    .Y(_9553_)
);

AOI21X1 _19210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9086_),
    .B(_9085_),
    .C(_9087_),
    .Y(_9091_)
);

FILL SFILL54120x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_38_),
    .C(_37_),
    .Y(_39_)
);

NAND3X1 _14189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3586_),
    .B(_3587_),
    .C(_3588_),
    .Y(_3589_)
);

FILL SFILL18760x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5205_),
    .B(_5202_),
    .C(_5194_),
    .Y(_5540_)
);

NAND3X1 _15550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5072_),
    .B(_5078_),
    .C(_5040_),
    .Y(_5079_)
);

AOI21X1 _15130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4063_),
    .B(_4315_),
    .C(_4619_),
    .Y(_4620_)
);

FILL SFILL18680x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _16755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6395_),
    .C(_6394_),
    .Y(_6401_)
);

NAND3X1 _16335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5929_),
    .B(_5940_),
    .C(_5937_),
    .Y(_5941_)
);

FILL SFILL54200x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert190 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551_),
    .Y(_4551__bF$buf1)
);

BUFX2 BUFX2_insert191 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551_),
    .Y(_4551__bF$buf0)
);

BUFX2 BUFX2_insert192 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402_),
    .Y(_3402__bF$buf3)
);

BUFX2 BUFX2_insert193 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402_),
    .Y(_3402__bF$buf2)
);

BUFX2 BUFX2_insert194 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402_),
    .Y(_3402__bF$buf1)
);

BUFX2 BUFX2_insert195 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402_),
    .Y(_3402__bF$buf0)
);

BUFX2 BUFX2_insert196 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711_),
    .Y(_7711__bF$buf3)
);

BUFX2 BUFX2_insert197 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711_),
    .Y(_7711__bF$buf2)
);

BUFX2 BUFX2_insert198 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711_),
    .Y(_7711__bF$buf1)
);

NAND2X1 _12675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_9_bF$buf1),
    .Y(_10748_)
);

BUFX2 BUFX2_insert199 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711_),
    .Y(_7711__bF$buf0)
);

NAND2X1 _12255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_7_bF$buf5),
    .Y(_6143_)
);

OAI21X1 _22773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_1084_),
    .C(_945_),
    .Y(_1089_)
);

NOR2X1 _22353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_628_),
    .Y(_629_)
);

NAND3X1 _18901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8745_),
    .B(_8751_),
    .C(_8752_),
    .Y(_8754_)
);

FILL SFILL69320x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23978_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[32]),
    .CLK(clk_bF$buf9),
    .D(_0_[32])
);

OAI21X1 _23558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(_1856_),
    .C(_1850_),
    .Y(_1944_)
);

AOI21X1 _23138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1484_),
    .B(_1485_),
    .C(_1479_),
    .Y(_1486_)
);

NOR3X1 _14821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_3982_),
    .C(_3985_),
    .Y(_4282_)
);

OAI21X1 _14401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf0),
    .B(_2586__bF$buf3),
    .C(_3595_),
    .Y(_3822_)
);

INVX1 _17293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6959_),
    .Y(_6991_)
);

NOR3X1 _15606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5138_),
    .B(_5139_),
    .C(_5140_),
    .Y(_5141_)
);

NAND3X1 _18498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8303_),
    .B(_8289_),
    .C(_8308_),
    .Y(_8312_)
);

NOR3X1 _18078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7837_),
    .B(_7834_),
    .C(_7836_),
    .Y(_7851_)
);

FILL SFILL38760x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_4_bF$buf4),
    .Y(_2759_)
);

FILL SFILL59240x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _21624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_6300__bF$buf3),
    .C(_3253__bF$buf0),
    .D(_5921__bF$buf3),
    .Y(_11738_)
);

AOI21X1 _21204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10967_),
    .B(_10970_),
    .C(_11278_),
    .Y(_11279_)
);

FILL SFILL24200x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64360x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3800x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_1038_),
    .C(_1148_),
    .Y(_1149_)
);

NAND3X1 _22409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_607_),
    .C(_668_),
    .Y(_689_)
);

FILL FILL74200x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_22_bF$buf0),
    .Y(_6651_)
);

OAI21X1 _16564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6189_),
    .B(_6190_),
    .C(_6188_),
    .Y(_6191_)
);

OAI21X1 _16144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5457_),
    .B(_5450_),
    .C(_5459_),
    .Y(_5731_)
);

AOI21X1 _17769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7118_),
    .B(_7115_),
    .C(_7107_),
    .Y(_7512_)
);

AOI21X1 _17349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7048_),
    .B(_7047_),
    .C(_7046_),
    .Y(_7052_)
);

NOR2X1 _12484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7207_),
    .B(_8632_),
    .Y(_8654_)
);

NAND3X1 _12064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3931_),
    .B(_3887_),
    .C(_3383_),
    .Y(_4051_)
);

NAND2X1 _22582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_879_),
    .Y(_880_)
);

AOI21X1 _22162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_409_),
    .B(_411_),
    .C(_403_),
    .Y(_420_)
);

OAI22X1 _18710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7786_),
    .B(_8541_),
    .C(_8542_),
    .D(_8189_),
    .Y(_8543_)
);

FILL SFILL33960x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2988_),
    .Y(_3042_)
);

INVX1 _13269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2581_),
    .Y(_2582_)
);

OR2X2 _23787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2191_),
    .B(_2189_),
    .Y(_2192_)
);

INVX1 _23367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1735_),
    .Y(_1736_)
);

AND2X2 _19915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_28_bF$buf1),
    .Y(_9866_)
);

FILL SFILL18760x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3783_),
    .B(_4068_),
    .C(_4070_),
    .Y(_4071_)
);

OAI21X1 _14210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3606_),
    .B(_3610_),
    .C(_3600_),
    .Y(_3611_)
);

OAI21X1 _15835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5391_),
    .B(_5390_),
    .C(_5380_),
    .Y(_5392_)
);

XOR2X1 _15415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .B(_4671_),
    .Y(_4933_)
);

OAI21X1 _21853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11807_),
    .B(_11805_),
    .C(_11799_),
    .Y(_81_)
);

OAI21X1 _21433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11230_),
    .B(_11528_),
    .C(_11529_),
    .Y(_11530_)
);

OR2X2 _21013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11062_),
    .B(_11063_),
    .Y(_11069_)
);

OAI21X1 _22638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_922_),
    .C(_939_),
    .Y(_940_)
);

NAND3X1 _22218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_244_),
    .B(_465_),
    .C(_471_),
    .Y(_481_)
);

INVX1 _13901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .Y(_3275_)
);

INVX1 _16793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6063_),
    .Y(_6442_)
);

NAND3X1 _16373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5975_),
    .B(_5981_),
    .C(_5838_),
    .Y(_5982_)
);

FILL SFILL13960x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7745_),
    .B(_7749_),
    .C(_7753_),
    .Y(_7763_)
);

NAND3X1 _17578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7295_),
    .B(_7299_),
    .C(_7301_),
    .Y(_7302_)
);

INVX1 _17158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6838_),
    .Y(_6842_)
);

FILL SFILL43880x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6549_),
    .B(_6461_),
    .C(_6505_),
    .Y(_6560_)
);

NAND3X1 _22391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_598_),
    .C(_601_),
    .Y(_670_)
);

FILL SFILL8600x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10729_),
    .B(_10725_),
    .C(_10701_),
    .Y(_10730_)
);

OAI21X1 _13498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2829_),
    .B(_2830_),
    .C(_2832_),
    .Y(_2833_)
);

XNOR2X1 _13078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2372_),
    .B(_2370_),
    .Y(_2373_)
);

NOR3X1 _23596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1258_),
    .B(_1540_),
    .C(_1984_),
    .Y(_1985_)
);

AOI21X1 _23176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1524_),
    .B(_1523_),
    .C(_1521_),
    .Y(_1528_)
);

AND2X2 _19724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_27_bF$buf2),
    .Y(_9656_)
);

AOI21X1 _19304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9194_),
    .B(_9195_),
    .C(_9191_),
    .Y(_9196_)
);

NAND3X1 _21909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_135_),
    .C(_139_),
    .Y(_142_)
);

FILL FILL74200x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_21_bF$buf1),
    .Y(_5183_)
);

NAND2X1 _15224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_13_bF$buf3),
    .Y(_4723_)
);

FILL SFILL33640x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6498_),
    .B(_6502_),
    .C(_6424_),
    .Y(_6503_)
);

NOR2X1 _16429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6038_),
    .B(_6041_),
    .Y(_6042_)
);

OAI21X1 _16009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5582_),
    .C(_5580_),
    .Y(_5583_)
);

XNOR2X1 _11984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3142_),
    .B(_3165_),
    .Y(_3176_)
);

NAND3X1 _21662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11755_),
    .B(_11779_),
    .C(_11770_),
    .Y(_11780_)
);

INVX2 _21242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11319_),
    .Y(_11320_)
);

FILL SFILL13880x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf2),
    .B(_6044__bF$buf2),
    .C(_10200_),
    .Y(_11778_)
);

XOR2X1 _12349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7164_),
    .B(_5947_),
    .Y(_0_[9])
);

NOR2X1 _22867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5369_),
    .B(_6686__bF$buf0),
    .Y(_1191_)
);

NOR2X1 _22447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_667_),
    .B(_439_),
    .Y(_731_)
);

AOI21X1 _22027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_270_),
    .C(_257_),
    .Y(_271_)
);

NOR2X1 _13710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3063_),
    .B(_3064_),
    .Y(_3065_)
);

NAND3X1 _16182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5766_),
    .B(_5767_),
    .C(_5772_),
    .Y(_5773_)
);

FILL SFILL8680x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4381_),
    .B(_4383_),
    .C(_4382_),
    .Y(_4384_)
);

NAND2X1 _17387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_25_bF$buf0),
    .Y(_7094_)
);

FILL SFILL23960x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10980_),
    .B(_10981_),
    .C(_10694_),
    .Y(_10982_)
);

OAI21X1 _20513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10515_),
    .B(_10516_),
    .C(_10520_),
    .Y(_10521_)
);

AOI21X1 _19953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_31_bF$buf0),
    .C(_9901_),
    .Y(_9907_)
);

AND2X2 _19533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9059_),
    .B(_9100_),
    .Y(_9447_)
);

NAND2X1 _19113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8932_),
    .B(_8929_),
    .Y(_8986_)
);

NAND3X1 _21718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11836_),
    .B(_11837_),
    .C(_11835_),
    .Y(_11841_)
);

AOI21X1 _15873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5415_),
    .B(_5418_),
    .C(_5422_),
    .Y(_5434_)
);

NAND2X1 _15453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_25_bF$buf0),
    .Y(_4973_)
);

OAI21X1 _15033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4236_),
    .B(_4239_),
    .C(_4513_),
    .Y(_4514_)
);

FILL SFILL53960x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_23_bF$buf4),
    .Y(_6294_)
);

NAND3X1 _16238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5832_),
    .B(_5833_),
    .C(_5831_),
    .Y(_5834_)
);

FILL SFILL59320x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_118_),
    .C(_103_),
    .Y(_123_)
);

NOR3X1 _21471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11279_),
    .B(_11274_),
    .C(_11266_),
    .Y(_11572_)
);

NAND3X1 _21051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11103_),
    .B(_11109_),
    .C(_11057_),
    .Y(_11111_)
);

NAND3X1 _12998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2292_),
    .C(_2249_),
    .Y(_2293_)
);

AOI21X1 _12578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9587_),
    .B(_9532_),
    .C(_8522_),
    .Y(_9685_)
);

NOR2X1 _12158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5058_),
    .B(_5069_),
    .Y(_5080_)
);

OAI21X1 _22676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_776_),
    .C(_784_),
    .Y(_982_)
);

AOI21X1 _22256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_517_),
    .C(_515_),
    .Y(_522_)
);

OAI21X1 _18804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf0),
    .B(_3146__bF$buf1),
    .C(_8641_),
    .Y(_8647_)
);

FILL SFILL13640x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33720x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4170_),
    .B(_4163_),
    .C(_4174_),
    .Y(_4175_)
);

AOI21X1 _14304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3429_),
    .B(_3385_),
    .C(_3432_),
    .Y(_3716_)
);

AOI21X1 _17196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6873_),
    .B(_6866_),
    .C(_6850_),
    .Y(_6884_)
);

NAND3X1 _15929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5494_),
    .B(_5493_),
    .C(_5492_),
    .Y(_5495_)
);

AOI21X1 _15509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5033_),
    .B(_5030_),
    .C(_5017_),
    .Y(_5034_)
);

AOI21X1 _20742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10483_),
    .B(_10488_),
    .C(_10469_),
    .Y(_10772_)
);

NOR3X1 _20322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9946_),
    .B(_9953_),
    .C(_9956_),
    .Y(_10312_)
);

INVX1 _19762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9691_),
    .Y(_9698_)
);

OAI21X1 _19342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9233_),
    .B(_9237_),
    .C(_8886_),
    .Y(_9238_)
);

FILL SFILL23720x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_180_),
    .Y(_184_)
);

OAI21X1 _21527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11631_),
    .B(_11624_),
    .C(_11609_),
    .Y(_11632_)
);

AND2X2 _21107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf4),
    .B(areg_25_bF$buf3),
    .Y(_11172_)
);

NAND2X1 _15682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5177_),
    .B(_5173_),
    .Y(_5224_)
);

NAND3X1 _15262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4761_),
    .B(_4764_),
    .C(_4762_),
    .Y(_4765_)
);

FILL SFILL8680x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6544_),
    .B(_6539_),
    .Y(_6545_)
);

NAND3X1 _16467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6079_),
    .B(_6066_),
    .C(_6069_),
    .Y(_6083_)
);

OAI21X1 _16047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5623_),
    .B(_5624_),
    .C(_5622_),
    .Y(_5625_)
);

NOR3X1 _21280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11345_),
    .B(_11332_),
    .C(_11352_),
    .Y(_11360_)
);

FILL SFILL48840x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_7_bF$buf1),
    .Y(_7591_)
);

NAND2X1 _22485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_567_),
    .Y(_773_)
);

NAND3X1 _22065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_305_),
    .B(_310_),
    .C(_312_),
    .Y(_313_)
);

NOR3X1 _18613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8012_),
    .B(_8018_),
    .C(_8021_),
    .Y(_8438_)
);

FILL SFILL74280x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_21_bF$buf4),
    .Y(_9759_)
);

OAI21X1 _14953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4425_),
    .B(_4424_),
    .C(_4420_),
    .Y(_4426_)
);

OAI21X1 _14533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_3961__bF$buf1),
    .C(_3680_),
    .Y(_3967_)
);

INVX1 _14113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .Y(_3506_)
);

OAI21X1 _15738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5275_),
    .B(_5276_),
    .C(_4969_),
    .Y(_5286_)
);

OAI21X1 _15318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf3),
    .B(_2884__bF$buf0),
    .C(_4821_),
    .Y(_4826_)
);

NAND2X1 _20971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_29_bF$buf4),
    .Y(_11023_)
);

NAND2X1 _20551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf1),
    .B(areg_28_bF$buf1),
    .Y(_10563_)
);

OAI21X1 _20131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10099_),
    .B(_10098_),
    .C(_10100_),
    .Y(_10102_)
);

NAND3X1 _19991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9645_),
    .B(_9750_),
    .C(_9752_),
    .Y(_9949_)
);

OAI21X1 _19571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9111_),
    .B(_9106_),
    .C(_9114_),
    .Y(_9489_)
);

NAND3X1 _19151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9022_),
    .B(_9026_),
    .C(_9014_),
    .Y(_9028_)
);

FILL SFILL64280x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _21756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11881_),
    .Y(_11882_)
);

NAND3X1 _21336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11421_),
    .B(_11420_),
    .C(_11422_),
    .Y(_11423_)
);

FILL SFILL33800x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4679_),
    .B(_5012_),
    .Y(_5015_)
);

AOI21X1 _15071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4542_),
    .B(_4540_),
    .C(_4538_),
    .Y(_4556_)
);

FILL SFILL33720x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3168_),
    .B(_3167_),
    .C(_3166_),
    .Y(_3169_)
);

BUFX2 _23902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[20]),
    .Y(y[20])
);

NOR3X1 _16696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5945_),
    .B(_5942_),
    .C(_5946_),
    .Y(_6336_)
);

AOI21X1 _16276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .B(_5536_),
    .C(_5533_),
    .Y(_5876_)
);

OAI22X1 _12196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3525_),
    .B(_5036_),
    .C(_4270_),
    .D(_4303_),
    .Y(_5497_)
);

AOI21X1 _22294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_562_),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

AOI21X1 _18842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8682_),
    .B(_8683_),
    .C(_8684_),
    .Y(_8689_)
);

AND2X2 _18422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf2),
    .B(areg_18_bF$buf5),
    .Y(_8229_)
);

NAND3X1 _18002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7767_),
    .B(_7760_),
    .C(_7764_),
    .Y(_7768_)
);

FILL SFILL23720x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10349_),
    .B(_10457_),
    .C(_10458_),
    .Y(_10624_)
);

NOR2X1 _23499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300__bF$buf2),
    .B(_6815__bF$buf3),
    .Y(_1879_)
);

NAND2X1 _23079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf0),
    .B(breg_29_bF$buf1),
    .Y(_1421_)
);

OAI21X1 _19627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9167_),
    .B(_9149_),
    .C(_9151_),
    .Y(_9550_)
);

NAND3X1 _19207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9086_),
    .B(_9087_),
    .C(_9085_),
    .Y(_9088_)
);

NAND3X1 _14762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4207_),
    .B(_4214_),
    .C(_4216_),
    .Y(_4217_)
);

NOR3X1 _14342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3736_),
    .B(_3742_),
    .C(_3744_),
    .Y(_3758_)
);

DFFPOSX1 _24020_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[10]),
    .CLK(clk_bF$buf0),
    .D(a[10])
);

NAND3X1 _15967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5522_),
    .B(_5526_),
    .C(_5528_),
    .Y(_5537_)
);

AOI21X1 _15547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5074_),
    .B(_5075_),
    .C(_5067_),
    .Y(_5076_)
);

NAND3X1 _15127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4614_),
    .B(_4616_),
    .C(_4615_),
    .Y(_4617_)
);

OAI21X1 _20780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10555_),
    .B(_10812_),
    .C(_10607_),
    .Y(_10813_)
);

OAI21X1 _20360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10019_),
    .B(_10005_),
    .C(_10029_),
    .Y(_10352_)
);

FILL SFILL8600x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf4),
    .B(_7225__bF$buf3),
    .Y(_9278_)
);

NAND3X1 _21985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_223_),
    .C(_11884_),
    .Y(_226_)
);

NAND3X1 _21565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11669_),
    .B(_11655_),
    .C(_11660_),
    .Y(_11673_)
);

AOI21X1 _21145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11207_),
    .B(_11208_),
    .C(_11206_),
    .Y(_11214_)
);

AOI21X1 _13613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2728_),
    .C(_2959_),
    .Y(_2960_)
);

AOI21X1 _23711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_2107_),
    .C(_2108_),
    .Y(_2110_)
);

FILL SFILL38840x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5363_),
    .B(_4996_),
    .C(_5356_),
    .Y(_5666_)
);

FILL SFILL43800x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4260_),
    .B(_4265_),
    .C(_4268_),
    .Y(_4278_)
);

NAND2X1 _18651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8174_),
    .B(_8179_),
    .Y(_8479_)
);

FILL SFILL64280x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8012_),
    .B(_8018_),
    .C(_7782_),
    .Y(_8019_)
);

OAI21X1 _20836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10870_),
    .B(_10871_),
    .C(_10874_),
    .Y(_10875_)
);

OAI21X1 _20416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf0),
    .B(_3781__bF$buf1),
    .C(_10056_),
    .Y(_10414_)
);

FILL SFILL28840x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf2),
    .B(_3961__bF$buf0),
    .C(_9797_),
    .Y(_9801_)
);

FILL SFILL64200x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9007_),
    .B(_9339_),
    .C(_9010_),
    .Y(_9340_)
);

AOI21X1 _19016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8876_),
    .B(_8877_),
    .C(_8878_),
    .Y(_8879_)
);

OAI21X1 _14991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4465_),
    .B(_4464_),
    .C(_4455_),
    .Y(_4467_)
);

NAND3X1 _14571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4001_),
    .B(_3915_),
    .C(_4002_),
    .Y(_4009_)
);

AND2X2 _14151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3542_),
    .Y(_3548_)
);

AOI21X1 _15776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5316_),
    .B(_5314_),
    .C(_5311_),
    .Y(_5327_)
);

NOR3X1 _15356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4855_),
    .B(_4859_),
    .C(_4864_),
    .Y(_4868_)
);

FILL SFILL18840x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(_11_),
    .C(_11893_),
    .Y(_16_)
);

AOI21X1 _21374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11464_),
    .B(_11459_),
    .C(_11445_),
    .Y(_11465_)
);

NAND2X1 _17922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_27_bF$buf3),
    .Y(_7680_)
);

INVX2 _17502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6843_),
    .Y(_7219_)
);

FILL SFILL74120x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1333_),
    .B(_1331_),
    .C(_1332_),
    .Y(_1334_)
);

XNOR2X1 _22579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_875_),
    .Y(_876_)
);

AOI21X1 _22159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_412_),
    .C(_402_),
    .Y(_416_)
);

NAND3X1 _18707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8537_),
    .B(_8539_),
    .C(_8538_),
    .Y(_8540_)
);

AOI21X1 _13842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3210_),
    .B(_3208_),
    .C(_3207_),
    .Y(_3211_)
);

XOR2X1 _13422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .B(_2750_),
    .Y(_0_[16])
);

BUFX2 _23940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[58]),
    .Y(y[58])
);

AOI21X1 _13002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2286_),
    .C(_2270_),
    .Y(_2297_)
);

OAI22X1 _23520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1703_),
    .B(_1811_),
    .C(_1814_),
    .D(_1810_),
    .Y(_1901_)
);

OAI21X1 _23100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1443_),
    .C(_1442_),
    .Y(_1444_)
);

NAND2X1 _14627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_22_bF$buf2),
    .Y(_4068_)
);

NAND2X1 _14207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(_3602_),
    .Y(_3608_)
);

NAND3X1 _17099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6423_),
    .B(_6771_),
    .C(_6777_),
    .Y(_6778_)
);

FILL SFILL44120x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8725_),
    .B(_8726_),
    .C(_8724_),
    .Y(_8730_)
);

NAND3X1 _18460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8254_),
    .B(_8261_),
    .C(_8222_),
    .Y(_8270_)
);

OAI21X1 _18040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7807_),
    .B(_7808_),
    .C(_7792_),
    .Y(_7809_)
);

NOR3X1 _20645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8868_),
    .B(_8473_),
    .C(_8865_),
    .Y(_10665_)
);

NAND2X1 _20225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10204_),
    .B(_10199_),
    .Y(_10205_)
);

NAND3X1 _19665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9383_),
    .B(_9376_),
    .C(_9381_),
    .Y(_9592_)
);

NAND3X1 _19245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9125_),
    .B(_9127_),
    .C(_9124_),
    .Y(_9131_)
);

AOI21X1 _14380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .B(_3797_),
    .C(_3786_),
    .Y(_3798_)
);

FILL SFILL44120x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5112_),
    .B(_5114_),
    .Y(_5118_)
);

NAND2X1 _15165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_24_bF$buf1),
    .Y(_4658_)
);

NAND3X1 _21183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11133_),
    .B(_11213_),
    .C(_11218_),
    .Y(_11256_)
);

OAI21X1 _17731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7089_),
    .B(_7066_),
    .C(_7079_),
    .Y(_7471_)
);

NAND3X1 _17311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6997_),
    .B(_7007_),
    .C(_7002_),
    .Y(_7010_)
);

NAND2X1 _22388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_666_),
    .Y(_667_)
);

NOR2X1 _18936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8783_),
    .B(_8789_),
    .Y(_8792_)
);

OAI21X1 _18516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8331_),
    .B(_7955_),
    .C(_7988_),
    .Y(_8332_)
);

NAND2X1 _13651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_12_bF$buf3),
    .Y(_3001_)
);

NOR2X1 _13231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2533_),
    .Y(_2541_)
);

NAND3X1 _14856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4317_),
    .B(_4318_),
    .C(_4319_),
    .Y(_4320_)
);

NAND3X1 _14436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3780_),
    .B(_3859_),
    .C(_3855_),
    .Y(_3860_)
);

AND2X2 _14016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_19_bF$buf2),
    .Y(_3400_)
);

FILL SFILL18840x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf4),
    .B(areg_29_bF$buf2),
    .Y(_10917_)
);

AND2X2 _20454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10091_),
    .B(_10083_),
    .Y(_10456_)
);

OAI21X1 _20034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9994_),
    .B(_9642_),
    .C(_9962_),
    .Y(_9995_)
);

NAND3X1 _19894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9837_),
    .B(_9836_),
    .C(_9835_),
    .Y(_9843_)
);

NAND3X1 _19474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9277_),
    .B(_9376_),
    .C(_9381_),
    .Y(_9382_)
);

NAND3X1 _19054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8905_),
    .B(_8898_),
    .C(_8910_),
    .Y(_8921_)
);

NOR2X1 _21659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11230_),
    .B(_11528_),
    .Y(_11776_)
);

AOI21X1 _21239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11293_),
    .B(_11294_),
    .C(_11009_),
    .Y(_11316_)
);

NOR2X1 _12922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10112_),
    .B(_11767_),
    .Y(_1543_)
);

AOI21X1 _12502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8786_),
    .B(_8830_),
    .C(_8851_),
    .Y(_8852_)
);

AOI21X1 _22600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_682_),
    .C(_693_),
    .Y(_899_)
);

OAI21X1 _15394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4896_),
    .B(_4897_),
    .C(_4814_),
    .Y(_4910_)
);

FILL SFILL69080x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf4),
    .B(breg_9_bF$buf3),
    .Y(_3062_)
);

OAI21X1 _23805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2208_),
    .B(_2117_),
    .C(_2210_),
    .Y(_2211_)
);

AND2X2 _16599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_19_bF$buf5),
    .Y(_6229_)
);

NOR2X1 _16179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5389_),
    .B(_5768_),
    .Y(_5769_)
);

NAND2X1 _17960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_22_bF$buf0),
    .Y(_7721_)
);

OAI21X1 _17540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6827_),
    .B(_6831_),
    .C(_6819_),
    .Y(_7260_)
);

NAND3X1 _17120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6800_),
    .B(_6799_),
    .C(_6404_),
    .Y(_6801_)
);

INVX8 _12099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf1),
    .Y(_4434_)
);

OAI21X1 _22197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_454_),
    .C(_445_),
    .Y(_458_)
);

NAND2X1 _18745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8524_),
    .B(_8520_),
    .Y(_8582_)
);

OAI21X1 _18325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7746_),
    .B(_7748_),
    .C(_7738_),
    .Y(_8122_)
);

FILL SFILL59080x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg_19_bF$buf3),
    .Y(_3251_)
);

AOI21X1 _13460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2692_),
    .B(_2697_),
    .C(_2626_),
    .Y(_2791_)
);

OAI21X1 _13040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2333_),
    .B(_2334_),
    .C(_1456_),
    .Y(_2335_)
);

FILL SFILL38920x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf0),
    .B(_2586__bF$buf3),
    .C(_3870_),
    .Y(_4110_)
);

OAI21X1 _14245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf1),
    .B(_2287__bF$buf2),
    .C(_3643_),
    .Y(_3651_)
);

FILL SFILL49480x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _20683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10706_),
    .Y(_10707_)
);

AOI21X1 _20263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10241_),
    .B(_10242_),
    .C(_10240_),
    .Y(_10247_)
);

FILL SFILL28920x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6070_),
    .B(_6134_),
    .Y(_6462_)
);

NAND2X1 _19283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_31_bF$buf0),
    .Y(_9173_)
);

NAND3X1 _21888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

OAI21X1 _21468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11551_),
    .B(_11557_),
    .C(_11559_),
    .Y(_11568_)
);

AOI21X1 _21048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11106_),
    .B(_11105_),
    .C(_11098_),
    .Y(_11107_)
);

OAI21X1 _12731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11361_),
    .B(_11297_),
    .C(_10002_),
    .Y(_11362_)
);

AOI21X1 _12311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6560_),
    .B(_6637_),
    .C(_6428_),
    .Y(_6758_)
);

FILL SFILL18920x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _13936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3312_),
    .Y(_3313_)
);

OAI21X1 _13516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_549__bF$buf4),
    .C(_2635_),
    .Y(_2853_)
);

AND2X2 _23614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1890_),
    .B(_1879_),
    .Y(_2005_)
);

NOR3X1 _18974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8400_),
    .B(_8407_),
    .C(_8410_),
    .Y(_8834_)
);

NAND3X1 _18554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8361_),
    .B(_8373_),
    .C(_8367_),
    .Y(_8374_)
);

AOI21X1 _18134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7911_),
    .B(_7912_),
    .C(_7910_),
    .Y(_7913_)
);

NAND3X1 _20739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10764_),
    .B(_10750_),
    .C(_10754_),
    .Y(_10768_)
);

NAND3X1 _20319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10291_),
    .B(_10297_),
    .C(_10301_),
    .Y(_10308_)
);

NOR2X1 _19759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9692_),
    .B(_9693_),
    .Y(_9694_)
);

NAND3X1 _19339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9231_),
    .B(_8890_),
    .C(_9230_),
    .Y(_9234_)
);

OAI21X1 _14894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4305_),
    .B(_4360_),
    .C(_4295_),
    .Y(_4361_)
);

OAI21X1 _14474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3894_),
    .B(_3900_),
    .C(_3901_),
    .Y(_3902_)
);

OAI21X1 _14054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3441_),
    .B(_3440_),
    .C(_3436_),
    .Y(_3442_)
);

AOI21X1 _15679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5206_),
    .B(_5210_),
    .C(_5193_),
    .Y(_5221_)
);

AOI21X1 _15259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4389_),
    .B(_4760_),
    .C(_4435_),
    .Y(_4761_)
);

INVX1 _20492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10149_),
    .Y(_10498_)
);

OAI21X1 _20072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10036_),
    .B(_10031_),
    .C(_10001_),
    .Y(_10037_)
);

AOI21X1 _16620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6247_),
    .B(_6248_),
    .C(_6246_),
    .Y(_6252_)
);

OAI21X1 _16200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf0),
    .B(_2362__bF$buf1),
    .C(_5785_),
    .Y(_5791_)
);

OAI21X1 _19092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8954_),
    .B(_8953_),
    .C(_8951_),
    .Y(_8963_)
);

OR2X2 _21697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11810_),
    .B(_11817_),
    .Y(_11818_)
);

AOI21X1 _21277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11356_),
    .B(_11353_),
    .C(_11330_),
    .Y(_11357_)
);

NAND3X1 _17825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7478_),
    .B(_7472_),
    .C(_7476_),
    .Y(_7574_)
);

INVX2 _17405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7113_),
    .Y(_7114_)
);

OAI21X1 _12960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_253_),
    .B(_1936_),
    .C(_1947_),
    .Y(_1957_)
);

AOI21X1 _12540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9126_),
    .B(_9170_),
    .C(_9038_),
    .Y(_9268_)
);

NOR3X1 _12120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4610_),
    .B(_4621_),
    .C(_4599_),
    .Y(_4664_)
);

FILL SFILL3640x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3102_),
    .B(_3103_),
    .Y(_3104_)
);

OAI21X1 _13325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2641_),
    .B(_2642_),
    .C(_2643_),
    .Y(_2644_)
);

XNOR2X1 _23843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2251_),
    .B(_2246_),
    .Y(_2252_)
);

OAI21X1 _23423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1789_),
    .B(_1795_),
    .C(_1796_),
    .Y(_1797_)
);

OAI21X1 _23003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1338_),
    .B(_1337_),
    .C(_1218_),
    .Y(_1339_)
);

NAND2X1 _18783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_8624_)
);

AOI21X1 _18363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8158_),
    .B(_8159_),
    .C(_8157_),
    .Y(_8164_)
);

FILL SFILL49000x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf2),
    .B(_6815__bF$buf0),
    .Y(_11019_)
);

XOR2X1 _20548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10511_),
    .B(_10558_),
    .Y(_10559_)
);

AOI21X1 _20128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10093_),
    .B(_10094_),
    .C(_10092_),
    .Y(_10098_)
);

NAND3X1 _19988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9941_),
    .B(_9944_),
    .C(_9940_),
    .Y(_9945_)
);

NAND2X1 _19568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_24_bF$buf1),
    .Y(_9485_)
);

NOR2X1 _19148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8624_),
    .B(_9023_),
    .Y(_9024_)
);

OAI21X1 _14283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3681_),
    .B(_3682_),
    .C(_3678_),
    .Y(_3693_)
);

FILL SFILL54280x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _15488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5010_),
    .Y(_5011_)
);

OAI21X1 _15068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_4551__bF$buf4),
    .C(_4539_),
    .Y(_4552_)
);

FILL SFILL39000x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _21086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf3),
    .B(_4541__bF$buf4),
    .C(_3253__bF$buf0),
    .D(_4551__bF$buf4),
    .Y(_11149_)
);

OAI21X1 _17634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf2),
    .B(_3529__bF$buf4),
    .C(_7354_),
    .Y(_7364_)
);

OAI21X1 _17214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6899_),
    .B(_6898_),
    .C(_6847_),
    .Y(_6904_)
);

FILL SFILL29080x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8682_),
    .B(_8684_),
    .C(_8683_),
    .Y(_8685_)
);

AOI21X1 _18419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7385_),
    .B(_8224_),
    .C(_7836_),
    .Y(_8225_)
);

OAI21X1 _13974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3347_),
    .B(_3346_),
    .C(_3348_),
    .Y(_3354_)
);

NAND3X1 _13554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2875_),
    .B(_2893_),
    .C(_2890_),
    .Y(_2894_)
);

NAND2X1 _13134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf3),
    .B(areg_9_bF$buf4),
    .Y(_2435_)
);

XOR2X1 _23652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_1998_),
    .Y(_2047_)
);

XNOR2X1 _23232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_1588_),
    .Y(_1589_)
);

NAND3X1 _14759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4208_),
    .B(_4212_),
    .C(_4211_),
    .Y(_4213_)
);

NOR3X1 _14339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3472_),
    .C(_3468_),
    .Y(_3754_)
);

DFFPOSX1 _24017_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[7]),
    .CLK(clk_bF$buf0),
    .D(a[7])
);

FILL SFILL74360x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4898_),
    .B(_4812_),
    .C(_4903_),
    .Y(_5243_)
);

AOI21X1 _18592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8408_),
    .B(_8414_),
    .C(_8279_),
    .Y(_8415_)
);

NAND2X1 _18172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7949_),
    .B(_7954_),
    .Y(_7955_)
);

NAND3X1 _20777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10808_),
    .B(_10809_),
    .C(_10807_),
    .Y(_10810_)
);

NAND2X1 _20357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10083_),
    .B(_10091_),
    .Y(_10349_)
);

AOI21X1 _16905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6557_),
    .B(_6558_),
    .C(_6550_),
    .Y(_6565_)
);

NAND3X1 _19797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9735_),
    .B(_9728_),
    .C(_9687_),
    .Y(_9736_)
);

AOI21X1 _19377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9216_),
    .B(_9217_),
    .C(_9004_),
    .Y(_9275_)
);

AOI21X1 _14092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3477_),
    .B(_3478_),
    .C(_3476_),
    .Y(_3484_)
);

FILL SFILL43880x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10825_),
    .B(_10880_),
    .C(_10913_),
    .Y(_484_)
);

NOR3X1 _12405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7667_),
    .B(_7744_),
    .C(_7755_),
    .Y(_7788_)
);

NAND2X1 _22923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1244_),
    .B(_1252_),
    .Y(_1253_)
);

AOI21X1 _22503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_635_),
    .B(_613_),
    .C(_792_),
    .Y(_793_)
);

AOI21X1 _15297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4788_),
    .B(_4792_),
    .C(_4773_),
    .Y(_4803_)
);

AOI21X1 _23708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .B(_1535_),
    .C(_1532_),
    .Y(_2106_)
);

AOI21X1 _17863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7597_),
    .B(_7603_),
    .C(_7341_),
    .Y(_7615_)
);

NAND3X1 _17443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7149_),
    .B(_7062_),
    .C(_7155_),
    .Y(_7156_)
);

NAND2X1 _17023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf4),
    .B(areg_27_bF$buf1),
    .Y(_6695_)
);

FILL SFILL33880x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8474_),
    .Y(_8475_)
);

NAND3X1 _18228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7880_),
    .B(_8009_),
    .C(_8010_),
    .Y(_8016_)
);

INVX8 _13783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .Y(_3146_)
);

AOI21X1 _13363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2473_),
    .C(_2477_),
    .Y(_2686_)
);

XOR2X1 _23881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3307_),
    .B(_3296_),
    .Y(_0_[4])
);

AOI21X1 _23461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1828_),
    .B(_1824_),
    .C(_1781_),
    .Y(_1839_)
);

FILL SFILL54280x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _23041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1232_),
    .C(_1225_),
    .Y(_1381_)
);

FILL SFILL23480x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_14_bF$buf0),
    .Y(_4463_)
);

OAI21X1 _14568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3911_),
    .B(_3910_),
    .C(_3868_),
    .Y(_4005_)
);

OAI21X1 _14148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf1),
    .B(_2362__bF$buf0),
    .C(_3266_),
    .Y(_3544_)
);

FILL SFILL23880x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8840x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _20586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10598_),
    .B(_10600_),
    .C(_10599_),
    .Y(_10601_)
);

FILL SFILL23800x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10138_),
    .B(_10139_),
    .C(_10137_),
    .Y(_10140_)
);

NAND3X1 _16714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6349_),
    .B(_6355_),
    .C(_6262_),
    .Y(_6356_)
);

OAI21X1 _19186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8644_),
    .B(_9065_),
    .C(_8646_),
    .Y(_9066_)
);

FILL SFILL8760x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7674_),
    .B(_7675_),
    .Y(_7676_)
);

NAND3X1 _12634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10266_),
    .B(_10288_),
    .C(_10277_),
    .Y(_10299_)
);

NAND3X1 _12214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5683_),
    .B(_5661_),
    .C(_5672_),
    .Y(_5694_)
);

NAND2X1 _22732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf4),
    .B(areg_28_bF$buf2),
    .Y(_1044_)
);

NAND3X1 _22312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(_581_),
    .C(_583_),
    .Y(_584_)
);

FILL SFILL29000x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3205_),
    .B(_3206_),
    .Y(_3207_)
);

NAND3X1 _13419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2549_),
    .B(_2741_),
    .C(_2742_),
    .Y(_2747_)
);

BUFX2 _23937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[55]),
    .Y(y[55])
);

NAND2X1 _23517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1815_),
    .Y(_1898_)
);

FILL SFILL43960x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7403_),
    .B(_7405_),
    .C(_7402_),
    .Y(_7406_)
);

OAI21X1 _17252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6940_),
    .B(_6945_),
    .C(_6932_),
    .Y(_6946_)
);

FILL SFILL49240x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8725_),
    .B(_8726_),
    .C(_8724_),
    .Y(_8727_)
);

AOI21X1 _18457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7881_),
    .B(_7915_),
    .C(_7924_),
    .Y(_8267_)
);

NAND3X1 _18037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7801_),
    .B(_7805_),
    .C(_7793_),
    .Y(_7806_)
);

AOI21X1 _13592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2625_),
    .B(_2702_),
    .C(_2936_),
    .Y(_2937_)
);

FILL FILL74120x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2471_),
    .B(_2457_),
    .C(_2472_),
    .Y(_2477_)
);

OAI21X1 _23690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1906_),
    .B(_2086_),
    .C(_2035_),
    .Y(_2087_)
);

NOR3X1 _23270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1628_),
    .B(_1553_),
    .C(_1629_),
    .Y(_1630_)
);

AOI21X1 _14797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3965_),
    .B(_3967_),
    .C(_3973_),
    .Y(_4254_)
);

OR2X2 _14377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3790_),
    .Y(_3795_)
);

DFFPOSX1 _24055_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[13]),
    .CLK(clk_bF$buf1),
    .D(b[13])
);

AND2X2 _20395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10387_),
    .B(_10390_),
    .Y(_10391_)
);

OAI21X1 _16943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf1),
    .B(_2884__bF$buf1),
    .C(_6561_),
    .Y(_6607_)
);

INVX2 _16523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6138_),
    .Y(_6146_)
);

OAI21X1 _16103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5674_),
    .B(_5685_),
    .C(_5682_),
    .Y(_5686_)
);

OAI21X1 _17728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7461_),
    .B(_7462_),
    .C(_7443_),
    .Y(_7467_)
);

AOI21X1 _17308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6603_),
    .B(_6645_),
    .C(_6642_),
    .Y(_7007_)
);

OAI21X1 _12863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(_878_),
    .C(_867_),
    .Y(_900_)
);

OAI21X1 _12443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8150_),
    .B(_8161_),
    .C(_7196_),
    .Y(_8205_)
);

AND2X2 _22961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1292_),
    .Y(_1294_)
);

INVX1 _12023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3591_),
    .Y(_3612_)
);

NAND2X1 _22541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_592_),
    .Y(_835_)
);

AOI21X1 _22121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_113_),
    .C(_106_),
    .Y(_375_)
);

FILL SFILL59080x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8920x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_2362__bF$buf0),
    .C(_2768_),
    .Y(_2997_)
);

AOI22X1 _13228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2349_),
    .B(_2352_),
    .C(_2534_),
    .D(_2535_),
    .Y(_2537_)
);

OAI21X1 _23746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1811_),
    .B(_2086_),
    .C(_2089_),
    .Y(_2148_)
);

NAND3X1 _23326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1665_),
    .B(_1690_),
    .C(_1689_),
    .Y(_1691_)
);

NAND3X1 _17481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6811_),
    .B(_7191_),
    .C(_7195_),
    .Y(_7197_)
);

NOR3X1 _17061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6338_),
    .B(_6339_),
    .C(_6337_),
    .Y(_6737_)
);

AOI21X1 _18686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8512_),
    .B(_8513_),
    .C(_8487_),
    .Y(_8517_)
);

OAI21X1 _18266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8054_),
    .B(_8057_),
    .C(_7654_),
    .Y(_8058_)
);

FILL SFILL13800x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .Y(_36_)
);

FILL SFILL29000x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3257_),
    .B(_3290_),
    .C(_3585_),
    .Y(_3586_)
);

FILL SFILL28840x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_12_bF$buf3),
    .Y(_1511_)
);

FILL SFILL64120x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6395_),
    .C(_6394_),
    .Y(_6398_)
);

NAND2X1 _16332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_27_bF$buf5),
    .Y(_5938_)
);

FILL SFILL19000x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert160 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf2)
);

BUFX2 BUFX2_insert161 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf1)
);

BUFX2 BUFX2_insert162 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf0)
);

BUFX2 BUFX2_insert163 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf5)
);

BUFX2 BUFX2_insert164 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf4)
);

OR2X2 _17957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7278_),
    .B(_7713_),
    .Y(_7718_)
);

BUFX2 BUFX2_insert165 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf3)
);

NAND3X1 _17537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7242_),
    .B(_7234_),
    .C(_7246_),
    .Y(_7257_)
);

BUFX2 BUFX2_insert166 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf2)
);

NAND3X1 _17117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6793_),
    .B(_6797_),
    .C(_6419_),
    .Y(_6798_)
);

BUFX2 BUFX2_insert167 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf1)
);

BUFX2 BUFX2_insert168 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[29]),
    .Y(areg_29_bF$buf0)
);

NOR2X1 _12672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf2),
    .B(_4434__bF$buf2),
    .Y(_10715_)
);

BUFX2 BUFX2_insert169 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884_),
    .Y(_2884__bF$buf3)
);

OAI21X1 _12252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5640_),
    .B(_5343_),
    .C(_5672_),
    .Y(_6110_)
);

INVX2 _22770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .Y(_1085_)
);

NOR2X1 _22350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_621_),
    .B(_624_),
    .Y(_625_)
);

OAI21X1 _13877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3047_),
    .B(_3247_),
    .C(_3208_),
    .Y(_3248_)
);

NAND2X1 _13457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2784_),
    .B(_2762_),
    .Y(_2788_)
);

DFFPOSX1 _23975_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[29]),
    .CLK(clk_bF$buf6),
    .D(_0_[29])
);

NAND3X1 _13037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .B(_2327_),
    .C(_2331_),
    .Y(_2332_)
);

NOR3X1 _23555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1928_),
    .B(_1929_),
    .C(_1873_),
    .Y(_1941_)
);

NAND3X1 _23135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1482_),
    .C(_1477_),
    .Y(_1483_)
);

AOI21X1 _17290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6969_),
    .B(_6973_),
    .C(_6976_),
    .Y(_6987_)
);

AOI21X1 _15603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5132_),
    .B(_5133_),
    .C(_5131_),
    .Y(_5138_)
);

NAND3X1 _18495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8302_),
    .B(_8303_),
    .C(_8308_),
    .Y(_8309_)
);

OAI21X1 _18075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7842_),
    .B(_7847_),
    .C(_7817_),
    .Y(_7848_)
);

NAND3X1 _16808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6451_),
    .B(_6454_),
    .C(_6457_),
    .Y(_6458_)
);

NAND2X1 _11943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf2),
    .B(breg_3_bF$buf0),
    .Y(_2727_)
);

NOR3X1 _21621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11728_),
    .B(_11730_),
    .C(_11733_),
    .Y(_11735_)
);

OAI21X1 _21201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11266_),
    .B(_11274_),
    .C(_11014_),
    .Y(_11276_)
);

FILL SFILL44040x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8920x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11264_),
    .B(_11275_),
    .C(_11253_),
    .Y(_11329_)
);

OAI21X1 _12308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6626_),
    .B(_6615_),
    .C(_6461_),
    .Y(_6725_)
);

NAND3X1 _22826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1143_),
    .B(_1138_),
    .C(_1145_),
    .Y(_1146_)
);

AOI21X1 _22406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .B(_463_),
    .C(_685_),
    .Y(_686_)
);

NAND2X1 _16981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6647_),
    .B(_6643_),
    .Y(_6648_)
);

AOI21X1 _16561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5412_),
    .B(_6168_),
    .C(_5799_),
    .Y(_6188_)
);

OAI21X1 _16141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5722_),
    .B(_5723_),
    .C(_5671_),
    .Y(_5728_)
);

AOI21X1 _17766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7495_),
    .B(_7498_),
    .C(_7499_),
    .Y(_7509_)
);

FILL SFILL74120x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7048_),
    .B(_7047_),
    .C(_7046_),
    .Y(_7049_)
);

OAI21X1 _12481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7228_),
    .B(_8588_),
    .C(_8610_),
    .Y(_8621_)
);

INVX1 _12061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4008_),
    .Y(_4019_)
);

AOI21X1 _13686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2835_),
    .B(_2833_),
    .C(_2837_),
    .Y(_3039_)
);

OAI21X1 _13266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2578_),
    .C(_2495_),
    .Y(_2579_)
);

NAND2X1 _23784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2188_),
    .B(_2187_),
    .Y(_2189_)
);

NAND2X1 _23364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_23_bF$buf2),
    .B(areg_31_bF$buf4),
    .Y(_1733_)
);

NAND2X1 _19912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf1),
    .B(areg_26_bF$buf4),
    .Y(_9863_)
);

NAND2X1 _15832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf0),
    .B(breg_18_bF$buf0),
    .Y(_5389_)
);

AOI21X1 _15412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4914_),
    .B(_4907_),
    .C(_4766_),
    .Y(_4930_)
);

AOI21X1 _20489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10493_),
    .B(_10492_),
    .C(_10491_),
    .Y(_10494_)
);

AOI21X1 _20069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10028_),
    .B(_10029_),
    .C(_10004_),
    .Y(_10033_)
);

NAND3X1 _16617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6247_),
    .B(_6248_),
    .C(_6246_),
    .Y(_6249_)
);

OAI21X1 _21850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .B(_73_),
    .C(_26_),
    .Y(_77_)
);

INVX2 _21430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11525_),
    .Y(_11526_)
);

AND2X2 _21010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11062_),
    .B(_11063_),
    .Y(_11065_)
);

NAND3X1 _19089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8936_),
    .B(_8952_),
    .C(_8958_),
    .Y(_8959_)
);

FILL FILL74040x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf2),
    .B(_5420__bF$buf0),
    .Y(_1925_)
);

NAND3X1 _12537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9181_),
    .B(_9225_),
    .C(_9027_),
    .Y(_9236_)
);

OAI21X1 _12117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4610_),
    .B(_4621_),
    .C(_4599_),
    .Y(_4632_)
);

OAI21X1 _22635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(_697_),
    .C(_936_),
    .Y(_937_)
);

NOR3X1 _22215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_217_),
    .C(_220_),
    .Y(_478_)
);

NAND2X1 _16790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6437_),
    .B(_6436_),
    .Y(_6438_)
);

OAI21X1 _16370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5972_),
    .B(_5973_),
    .C(_5886_),
    .Y(_5979_)
);

NAND3X1 _17995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7759_),
    .B(_7750_),
    .C(_7706_),
    .Y(_7760_)
);

NAND3X1 _17575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7296_),
    .B(_7297_),
    .C(_7298_),
    .Y(_7299_)
);

OAI21X1 _17155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6837_),
    .B(_6832_),
    .C(_6817_),
    .Y(_6839_)
);

NOR2X1 _12290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5179_),
    .B(_6483_),
    .Y(_6527_)
);

OAI21X1 _20701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10722_),
    .B(_10723_),
    .C(_10719_),
    .Y(_10727_)
);

FILL SFILL44040x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2819_),
    .B(_2811_),
    .C(_2800_),
    .Y(_2830_)
);

NOR2X1 _13075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2367_),
    .B(_2369_),
    .Y(_2370_)
);

AND2X2 _23593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1763_),
    .B(_1767_),
    .Y(_1982_)
);

NAND3X1 _23173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1521_),
    .B(_1524_),
    .C(_1523_),
    .Y(_1525_)
);

NAND2X1 _19721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_29_bF$buf0),
    .Y(_9653_)
);

NAND2X1 _19301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8787_),
    .B(_8813_),
    .Y(_9193_)
);

NAND3X1 _21906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_137_),
    .C(_138_),
    .Y(_139_)
);

AOI21X1 _15641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4865_),
    .B(_4861_),
    .C(_4854_),
    .Y(_5180_)
);

OAI21X1 _15221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf0),
    .B(_2560__bF$buf4),
    .C(_4715_),
    .Y(_4720_)
);

FILL SFILL34040x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10208_),
    .B(_10273_),
    .Y(_10285_)
);

NAND3X1 _16846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6438_),
    .B(_6490_),
    .C(_6486_),
    .Y(_6500_)
);

AOI21X1 _16426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5654_),
    .B(_5657_),
    .C(_6033_),
    .Y(_6039_)
);

AOI21X1 _16006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5210_),
    .B(_5193_),
    .C(_5579_),
    .Y(_5580_)
);

NOR2X1 _11981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3110_),
    .B(_3142_),
    .Y(_3143_)
);

FILL SFILL69160x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11734_),
    .B(_11723_),
    .Y(_11745_)
);

OAI21X1 _12346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7087_),
    .B(_7065_),
    .C(_6012_),
    .Y(_7142_)
);

NAND3X1 _22864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1186_),
    .C(_1187_),
    .Y(_1188_)
);

FILL SFILL59240x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_694_),
    .B(_499_),
    .C(_681_),
    .Y(_728_)
);

NOR2X1 _22024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11905_),
    .B(_267_),
    .Y(_268_)
);

FILL SFILL24040x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _23649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .B(_2042_),
    .Y(_2043_)
);

NAND3X1 _23229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1579_),
    .C(_1583_),
    .Y(_1584_)
);

OAI21X1 _14912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4080_),
    .B(_4075_),
    .C(_4084_),
    .Y(_4381_)
);

NAND2X1 _17384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7084_),
    .B(_7090_),
    .Y(_7091_)
);

FILL SFILL59160x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10977_),
    .B(_10972_),
    .C(_10695_),
    .Y(_10978_)
);

NOR2X1 _20510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10157_),
    .B(_10212_),
    .Y(_10517_)
);

NAND3X1 _18589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8405_),
    .B(_8406_),
    .C(_8404_),
    .Y(_8411_)
);

NAND3X1 _18169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7947_),
    .B(_7938_),
    .C(_7941_),
    .Y(_7951_)
);

NOR2X1 _19950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_9153_),
    .Y(_9903_)
);

AOI21X1 _19530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9436_),
    .B(_9437_),
    .C(_9428_),
    .Y(_9443_)
);

AOI21X1 _19110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8973_),
    .B(_8967_),
    .C(_8935_),
    .Y(_8982_)
);

FILL SFILL54120x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11836_),
    .B(_11837_),
    .C(_11835_),
    .Y(_11838_)
);

NAND3X1 _14089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3475_),
    .B(_3245_),
    .C(_3479_),
    .Y(_3480_)
);

FILL SFILL49160x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5407_),
    .B(_5423_),
    .C(_5429_),
    .Y(_5430_)
);

OAI21X1 _15450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4968_),
    .B(_4933_),
    .C(_4923_),
    .Y(_4969_)
);

OAI21X1 _15030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_2884__bF$buf0),
    .C(_4503_),
    .Y(_4510_)
);

FILL SFILL39160x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6290_),
    .B(_6285_),
    .Y(_6291_)
);

AND2X2 _16235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5444_),
    .B(_5436_),
    .Y(_5831_)
);

FILL SFILL59400x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_2280_),
    .Y(_2290_)
);

NOR3X1 _12575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8150_),
    .B(_8161_),
    .C(_8139_),
    .Y(_9652_)
);

NAND2X1 _12155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_3_bF$buf0),
    .Y(_5047_)
);

AND2X2 _22673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_978_),
    .Y(_979_)
);

NAND3X1 _22253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_518_),
    .C(_517_),
    .Y(_519_)
);

NAND2X1 _18801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf3),
    .B(areg_18_bF$buf5),
    .Y(_8644_)
);

FILL SFILL69320x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf3),
    .B(_2376__bF$buf3),
    .Y(_0_[0])
);

NAND2X1 _23458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1826_),
    .Y(_1835_)
);

NAND3X1 _23038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1372_),
    .C(_1373_),
    .Y(_1377_)
);

FILL SFILL69240x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4166_),
    .B(_4167_),
    .Y(_4172_)
);

OAI21X1 _14301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3699_),
    .B(_3695_),
    .C(_3703_),
    .Y(_3713_)
);

OAI21X1 _17193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6517_),
    .B(_6880_),
    .C(_6542_),
    .Y(_6881_)
);

XNOR2X1 _15926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5470_),
    .B(_5466_),
    .Y(_5492_)
);

NAND3X1 _15506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5026_),
    .B(_5028_),
    .C(_5027_),
    .Y(_5031_)
);

AOI21X1 _18398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8199_),
    .B(_8201_),
    .C(_8197_),
    .Y(_8202_)
);

NAND3X1 _21944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_180_),
    .C(_171_),
    .Y(_181_)
);

AOI21X1 _21524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11627_),
    .B(_11628_),
    .C(_11611_),
    .Y(_11629_)
);

OAI21X1 _21104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10863_),
    .B(_10853_),
    .C(_10857_),
    .Y(_11169_)
);

FILL SFILL3800x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _22729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1039_),
    .B(_1037_),
    .Y(_1040_)
);

INVX2 _22309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .Y(_580_)
);

FILL FILL74200x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6532_),
    .B(_6518_),
    .C(_6536_),
    .Y(_6542_)
);

OAI21X1 _16464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6074_),
    .B(_6075_),
    .C(_6079_),
    .Y(_6080_)
);

AOI21X1 _16044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5248_),
    .B(_5101_),
    .C(_5253_),
    .Y(_5622_)
);

FILL SFILL28760x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _17669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7380_),
    .Y(_7402_)
);

NAND2X1 _17249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6937_),
    .B(_6938_),
    .Y(_6942_)
);

OAI21X1 _12384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6681_),
    .B(_6659_),
    .C(_6560_),
    .Y(_7558_)
);

AND2X2 _22482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_769_),
    .Y(_770_)
);

NAND3X1 _22062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_309_),
    .C(_307_),
    .Y(_310_)
);

OAI21X1 _18610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8415_),
    .B(_8421_),
    .C(_8425_),
    .Y(_8434_)
);

FILL SFILL8600x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2931_),
    .B(_2932_),
    .C(_2930_),
    .Y(_2933_)
);

OAI21X1 _13169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2472_),
    .B(_2471_),
    .C(_2457_),
    .Y(_2473_)
);

INVX1 _23687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .Y(_2084_)
);

NAND2X1 _23267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .B(_1626_),
    .Y(_1627_)
);

OAI21X1 _19815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9481_),
    .B(_9755_),
    .C(_9581_),
    .Y(_9756_)
);

FILL SFILL18760x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4410_),
    .B(_4411_),
    .C(_4408_),
    .Y(_4422_)
);

AOI21X1 _14530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3960_),
    .B(_3962_),
    .C(_3957_),
    .Y(_3963_)
);

AND2X2 _14110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1228_),
    .B(_1282_),
    .Y(_3502_)
);

FILL SFILL33720x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39160x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5281_),
    .B(_5282_),
    .C(_5280_),
    .Y(_5283_)
);

OAI22X1 _15315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_3146__bF$buf0),
    .C(_4116__bF$buf3),
    .D(_2884__bF$buf2),
    .Y(_4823_)
);

BUFX2 BUFX2_insert70 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .Y(_6815__bF$buf3)
);

BUFX2 BUFX2_insert71 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .Y(_6815__bF$buf2)
);

BUFX2 BUFX2_insert72 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .Y(_6815__bF$buf1)
);

BUFX2 BUFX2_insert73 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .Y(_6815__bF$buf0)
);

BUFX2 BUFX2_insert74 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(areg_12_bF$buf4)
);

BUFX2 BUFX2_insert75 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(areg_12_bF$buf3)
);

BUFX2 BUFX2_insert76 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(areg_12_bF$buf2)
);

BUFX2 BUFX2_insert77 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(areg_12_bF$buf1)
);

BUFX2 BUFX2_insert78 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[12]),
    .Y(areg_12_bF$buf0)
);

BUFX2 BUFX2_insert79 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[22]),
    .Y(breg_22_bF$buf4)
);

FILL SFILL23960x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11873_),
    .B(_11878_),
    .Y(_11879_)
);

NAND2X1 _21333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11367_),
    .B(_11364_),
    .Y(_11420_)
);

FILL SFILL69320x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf3),
    .B(_7225__bF$buf0),
    .C(_1289_),
    .Y(_1290_)
);

AOI21X1 _22538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_816_),
    .B(_821_),
    .C(_770_),
    .Y(_831_)
);

AND2X2 _22118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_368_),
    .Y(_370_)
);

AND2X2 _13801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3138_),
    .B(_3134_),
    .Y(_3166_)
);

NAND3X1 _16693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6321_),
    .B(_6323_),
    .C(_6316_),
    .Y(_6333_)
);

AOI21X1 _16273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5871_),
    .B(_5866_),
    .C(_5872_),
    .Y(_5873_)
);

AOI21X1 _17898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7617_),
    .B(_7621_),
    .C(_7220_),
    .Y(_7653_)
);

AOI21X1 _17478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7189_),
    .B(_7188_),
    .C(_7187_),
    .Y(_7193_)
);

NAND3X1 _17058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6716_),
    .B(_6720_),
    .C(_6723_),
    .Y(_6733_)
);

OAI21X1 _12193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf2),
    .B(_5453__bF$buf1),
    .C(_4083_),
    .Y(_5464_)
);

INVX1 _22291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_545_),
    .Y(_561_)
);

FILL SFILL8600x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10619_),
    .B(_10620_),
    .C(_10618_),
    .Y(_10621_)
);

AOI21X1 _13398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2374_),
    .B(_2512_),
    .C(_2723_),
    .Y(_2724_)
);

NOR2X1 _23496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .B(_1792_),
    .Y(_1876_)
);

OAI21X1 _23076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921__bF$buf1),
    .B(_5668__bF$buf1),
    .C(_1275_),
    .Y(_1418_)
);

AOI21X1 _19624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9538_),
    .B(_9536_),
    .C(_9534_),
    .Y(_9547_)
);

NAND3X1 _19204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9080_),
    .B(_9081_),
    .C(_9079_),
    .Y(_9085_)
);

NOR2X1 _21809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_31_),
    .Y(_32_)
);

FILL FILL74200x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5529_),
    .B(_5533_),
    .C(_5515_),
    .Y(_5534_)
);

AOI21X1 _15544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4711_),
    .B(_4733_),
    .C(_4736_),
    .Y(_5073_)
);

XNOR2X1 _15124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4358_),
    .B(_4356_),
    .Y(_4614_)
);

AOI21X1 _16749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5743_),
    .B(_6002_),
    .C(_6393_),
    .Y(_6394_)
);

AOI22X1 _16329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf5),
    .B(areg_27_bF$buf3),
    .C(breg_1_bF$buf1),
    .D(areg_26_bF$buf2),
    .Y(_5934_)
);

NAND3X1 _21982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11886_),
    .B(_197_),
    .C(_213_),
    .Y(_223_)
);

OAI21X1 _21562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11665_),
    .B(_11666_),
    .C(_11669_),
    .Y(_11670_)
);

NOR3X1 _21142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10942_),
    .B(_10940_),
    .C(_10941_),
    .Y(_11211_)
);

FILL SFILL38600x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10650_),
    .B(_10661_),
    .C(_10671_),
    .Y(_10682_)
);

OAI21X1 _12249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6076_),
    .B(_4105_),
    .C(_5508_),
    .Y(_6087_)
);

NAND3X1 _22767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_1073_),
    .C(_1069_),
    .Y(_1082_)
);

NAND2X1 _22347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_28_bF$buf2),
    .Y(_622_)
);

NAND3X1 _13610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2756_),
    .B(_2954_),
    .C(_2955_),
    .Y(_2956_)
);

OAI21X1 _16082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5302_),
    .B(_5662_),
    .C(_5660_),
    .Y(_5663_)
);

OAI21X1 _14815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4230_),
    .B(_4231_),
    .C(_4206_),
    .Y(_4275_)
);

NAND3X1 _17287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6960_),
    .B(_6983_),
    .C(_6978_),
    .Y(_6984_)
);

FILL SFILL23960x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10511_),
    .B(_10558_),
    .Y(_10872_)
);

AOI21X1 _20413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10404_),
    .B(_10403_),
    .C(_10402_),
    .Y(_10411_)
);

NAND2X1 _19853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9792_),
    .B(_9797_),
    .Y(_9798_)
);

AOI21X1 _19433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9331_),
    .B(_9330_),
    .C(_9329_),
    .Y(_9337_)
);

XNOR2X1 _19013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8471_),
    .B(_8876_),
    .Y(_0_[34])
);

AND2X2 _21618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_24_bF$buf4),
    .Y(_11731_)
);

OAI21X1 _15773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5015_),
    .B(_5010_),
    .C(_5323_),
    .Y(_5324_)
);

OAI21X1 _15353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4864_),
    .B(_4859_),
    .C(_4855_),
    .Y(_4865_)
);

FILL SFILL13560x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6639_),
    .B(_6640_),
    .C(_6641_),
    .Y(_6645_)
);

AOI21X1 _16558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5841_),
    .B(_5843_),
    .C(_6183_),
    .Y(_6184_)
);

OAI21X1 _16138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5722_),
    .B(_5723_),
    .C(_5721_),
    .Y(_5724_)
);

FILL SFILL59320x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11893_),
    .B(_10_),
    .C(_11_),
    .Y(_13_)
);

NAND3X1 _21371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11455_),
    .B(_11457_),
    .C(_11456_),
    .Y(_11462_)
);

AOI21X1 _12898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11603_),
    .B(_11614_),
    .C(_9762_),
    .Y(_1282_)
);

NAND2X1 _12478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_10_bF$buf5),
    .Y(_8588_)
);

NAND2X1 _22996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1292_),
    .B(_1290_),
    .Y(_1331_)
);

INVX1 _12058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3975_),
    .Y(_3986_)
);

NOR2X1 _22576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_870_),
    .B(_865_),
    .Y(_873_)
);

OR2X2 _22156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_11528_),
    .Y(_413_)
);

INVX1 _18704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8530_),
    .Y(_8537_)
);

XOR2X1 _19909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9811_),
    .B(_9858_),
    .Y(_9859_)
);

OAI21X1 _14624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3866_),
    .B(_4064_),
    .C(_4022_),
    .Y(_4065_)
);

OAI21X1 _14204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_9104__bF$buf2),
    .C(_3604_),
    .Y(_3605_)
);

NOR3X1 _17096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6767_),
    .B(_6768_),
    .C(_6766_),
    .Y(_6775_)
);

NAND2X1 _15829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf4),
    .B(breg_19_bF$buf2),
    .Y(_5385_)
);

OAI21X1 _15409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4912_),
    .B(_4913_),
    .C(_4768_),
    .Y(_4926_)
);

NOR3X1 _20642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8453_),
    .B(_8456_),
    .C(_8459_),
    .Y(_10662_)
);

OAI21X1 _20222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10195_),
    .B(_10194_),
    .C(_10197_),
    .Y(_10202_)
);

NAND3X1 _19662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9571_),
    .B(_9575_),
    .C(_9481_),
    .Y(_9589_)
);

AOI21X1 _19242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9125_),
    .B(_9127_),
    .C(_9124_),
    .Y(_9128_)
);

OAI21X1 _21847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_72_),
    .B(_73_),
    .C(_71_),
    .Y(_74_)
);

INVX1 _21427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11241_),
    .Y(_11523_)
);

NAND2X1 _21007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf4),
    .B(breg_25_bF$buf0),
    .Y(_11062_)
);

NAND2X1 _15582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5112_),
    .B(_5114_),
    .Y(_5115_)
);

AOI21X1 _15162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4598_),
    .B(_4605_),
    .C(_4361_),
    .Y(_4655_)
);

NOR2X1 _16787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6426_),
    .B(_6434_),
    .Y(_6435_)
);

NAND3X1 _16367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5839_),
    .B(_5880_),
    .C(_5882_),
    .Y(_5976_)
);

NAND2X1 _21180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11251_),
    .B(_11248_),
    .Y(_11252_)
);

FILL SFILL8600x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _12287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5179_),
    .B(_6483_),
    .Y(_6494_)
);

NOR3X1 _22385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_657_),
    .B(_656_),
    .C(_660_),
    .Y(_664_)
);

AOI22X1 _18933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8787_),
    .B(_8788_),
    .C(_8785_),
    .D(_8784_),
    .Y(_8789_)
);

OAI21X1 _18513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8328_),
    .B(_8327_),
    .C(_8325_),
    .Y(_8329_)
);

FILL SFILL74280x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf1),
    .B(_6815__bF$buf2),
    .Y(_9649_)
);

XNOR2X1 _14853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4062_),
    .B(_4060_),
    .Y(_4317_)
);

AOI22X1 _14433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3802_),
    .B(_3805_),
    .C(_3847_),
    .D(_3838_),
    .Y(_3857_)
);

NAND2X1 _14013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf1),
    .B(areg_17_bF$buf1),
    .Y(_3397_)
);

OAI21X1 _15638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5167_),
    .B(_5169_),
    .C(_5165_),
    .Y(_5176_)
);

NAND2X1 _15218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4714_),
    .B(_4715_),
    .Y(_4716_)
);

XOR2X1 _20871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10865_),
    .B(_10912_),
    .Y(_10914_)
);

AOI21X1 _20451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10110_),
    .B(_10202_),
    .C(_10198_),
    .Y(_10453_)
);

AOI21X1 _20031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9637_),
    .B(_9973_),
    .C(_9990_),
    .Y(_9992_)
);

NOR3X1 _19891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9519_),
    .B(_9520_),
    .C(_9518_),
    .Y(_9840_)
);

AOI21X1 _19471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9369_),
    .B(_9360_),
    .C(_9317_),
    .Y(_9379_)
);

NOR3X1 _19051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8916_),
    .B(_8912_),
    .C(_8915_),
    .Y(_8918_)
);

AOI21X1 _11978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3099_),
    .B(_3088_),
    .C(_3066_),
    .Y(_3110_)
);

OAI21X1 _21656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf1),
    .B(_7520__bF$buf1),
    .C(_11758_),
    .Y(_11773_)
);

AOI22X1 _21236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11301_),
    .B(_11306_),
    .C(_10993_),
    .D(_10997_),
    .Y(_11313_)
);

FILL SFILL64200x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4768_),
    .B(_4899_),
    .C(_4905_),
    .Y(_4907_)
);

AOI21X1 _13704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2806_),
    .B(_2808_),
    .C(_2816_),
    .Y(_3059_)
);

NAND2X1 _23802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2202_),
    .B(_2159_),
    .Y(_2208_)
);

OAI21X1 _16596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5856_),
    .B(_5847_),
    .C(_5851_),
    .Y(_6226_)
);

AOI21X1 _16176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5381_),
    .B(_5386_),
    .C(_5390_),
    .Y(_5766_)
);

OAI21X1 _14909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf2),
    .B(_3529__bF$buf0),
    .C(_4076_),
    .Y(_4377_)
);

XOR2X1 _12096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3635_),
    .B(_4390_),
    .Y(_4401_)
);

NOR2X1 _22194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_453_),
    .B(_454_),
    .Y(_455_)
);

AOI21X1 _18742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8565_),
    .B(_8560_),
    .C(_8528_),
    .Y(_8579_)
);

NAND3X1 _18322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8082_),
    .B(_8110_),
    .C(_8107_),
    .Y(_8119_)
);

FILL SFILL23720x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10969_),
    .B(_10967_),
    .C(_10970_),
    .Y(_10975_)
);

NAND3X1 _20507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10506_),
    .B(_10510_),
    .C(_10513_),
    .Y(_10514_)
);

NAND2X1 _23399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1763_),
    .B(_1769_),
    .Y(_1770_)
);

NAND3X1 _19947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9897_),
    .B(_9898_),
    .C(_9899_),
    .Y(_9900_)
);

OAI21X1 _19527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_4541__bF$buf0),
    .C(_9059_),
    .Y(_9440_)
);

NAND3X1 _19107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8974_),
    .B(_8978_),
    .C(_8934_),
    .Y(_8979_)
);

NAND2X1 _14662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4104_),
    .B(_4103_),
    .Y(_4107_)
);

NAND3X1 _14242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3642_),
    .B(_3647_),
    .C(_3645_),
    .Y(_3648_)
);

OAI21X1 _15867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf3),
    .B(_549__bF$buf1),
    .C(_5055_),
    .Y(_5427_)
);

INVX1 _15447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .Y(_4966_)
);

NAND3X1 _15027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4502_),
    .B(_4506_),
    .C(_4505_),
    .Y(_4507_)
);

INVX2 _20680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10702_),
    .Y(_10703_)
);

NAND3X1 _20260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10241_),
    .B(_10242_),
    .C(_10240_),
    .Y(_10243_)
);

FILL SFILL13720x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9151_),
    .B(_9155_),
    .C(_9164_),
    .Y(_9169_)
);

AOI21X1 _21885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11736_),
    .B(_11738_),
    .C(_11730_),
    .Y(_116_)
);

NAND3X1 _21465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11564_),
    .B(_11561_),
    .C(_11559_),
    .Y(_11565_)
);

AOI21X1 _21045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10742_),
    .B(_10779_),
    .C(_10783_),
    .Y(_11104_)
);

OAI21X1 _13933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3095_),
    .B(_3201_),
    .C(_3192_),
    .Y(_3310_)
);

OAI21X1 _13513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_9104__bF$buf1),
    .C(_2631_),
    .Y(_2850_)
);

NOR2X1 _23611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300__bF$buf2),
    .B(_7225__bF$buf2),
    .Y(_2002_)
);

FILL SFILL74200x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4166_),
    .B(_4167_),
    .Y(_4168_)
);

OAI21X1 _18971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8794_),
    .B(_8801_),
    .C(_8804_),
    .Y(_8831_)
);

NOR2X1 _18551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8368_),
    .B(_8369_),
    .Y(_8371_)
);

XNOR2X1 _18131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7885_),
    .B(_7882_),
    .Y(_7910_)
);

OAI21X1 _20736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10761_),
    .B(_10760_),
    .C(_10764_),
    .Y(_10765_)
);

NAND3X1 _20316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9996_),
    .B(_10304_),
    .C(_10298_),
    .Y(_10305_)
);

FILL SFILL33800x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_26_bF$buf3),
    .Y(_9691_)
);

NAND3X1 _19336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9002_),
    .B(_9218_),
    .C(_9212_),
    .Y(_9231_)
);

NAND2X1 _14891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4141_),
    .B(_4302_),
    .Y(_4358_)
);

OAI21X1 _14471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3881_),
    .B(_3885_),
    .C(_3888_),
    .Y(_3899_)
);

NAND3X1 _14051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3423_),
    .B(_3419_),
    .C(_3425_),
    .Y(_3439_)
);

NOR3X1 _15676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4868_),
    .B(_4867_),
    .C(_4869_),
    .Y(_5218_)
);

NOR3X1 _15256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4757_),
    .B(_4755_),
    .C(_4756_),
    .Y(_4758_)
);

FILL SFILL44040x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL58920x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11528_),
    .B(_11813_),
    .Y(_11815_)
);

OAI21X1 _21274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11349_),
    .B(_11351_),
    .C(_11346_),
    .Y(_11354_)
);

AOI21X1 _17822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7552_),
    .B(_7557_),
    .C(_7511_),
    .Y(_7571_)
);

AND2X2 _17402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf5),
    .B(areg_30_bF$buf5),
    .Y(_7111_)
);

FILL SFILL74120x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23720x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1223_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1226_)
);

NAND3X1 _22479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .B(_762_),
    .C(_763_),
    .Y(_766_)
);

INVX1 _22059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .Y(_306_)
);

NAND3X1 _18607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8079_),
    .B(_8181_),
    .C(_8182_),
    .Y(_8431_)
);

INVX1 _13742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3100_),
    .Y(_3101_)
);

AND2X2 _13322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2640_),
    .B(_2630_),
    .Y(_2641_)
);

OAI22X1 _23840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2139_),
    .B(_2179_),
    .C(_2247_),
    .D(_2224_),
    .Y(_2248_)
);

NAND2X1 _23420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_25_bF$buf1),
    .B(breg_29_bF$buf1),
    .Y(_1793_)
);

NAND3X1 _23000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1216_),
    .B(_1334_),
    .C(_1330_),
    .Y(_1335_)
);

FILL SFILL48920x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44200x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4414_),
    .B(_4418_),
    .C(_4389_),
    .Y(_4419_)
);

OAI21X1 _14527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_3958__bF$buf2),
    .C(_3959_),
    .Y(_3960_)
);

NAND2X1 _14107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .B(_2532_),
    .Y(_3499_)
);

OAI21X1 _18780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8616_),
    .B(_8619_),
    .C(_8608_),
    .Y(_8620_)
);

NAND3X1 _18360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8157_),
    .B(_8158_),
    .C(_8159_),
    .Y(_8160_)
);

NOR2X1 _20965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf2),
    .B(_7225__bF$buf4),
    .Y(_11016_)
);

NAND2X1 _20545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10229_),
    .B(_10238_),
    .Y(_10556_)
);

NAND3X1 _20125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10092_),
    .B(_10093_),
    .C(_10094_),
    .Y(_10095_)
);

AND2X2 _19985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9928_),
    .B(_9855_),
    .Y(_9942_)
);

OAI21X1 _19565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9141_),
    .B(_9201_),
    .C(_9194_),
    .Y(_9482_)
);

OAI21X1 _19145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf3),
    .B(_3529__bF$buf4),
    .C(_8624_),
    .Y(_9021_)
);

OAI21X1 _14280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .B(_3683_),
    .C(_3677_),
    .Y(_3689_)
);

FILL SFILL38920x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4921_),
    .B(_4919_),
    .C(_4907_),
    .Y(_5008_)
);

NAND3X1 _15065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4536_),
    .B(_4543_),
    .C(_4548_),
    .Y(_4549_)
);

AOI21X1 _21083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11142_),
    .B(_11145_),
    .C(_11140_),
    .Y(_11146_)
);

NOR3X1 _17631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7353_),
    .B(_7356_),
    .C(_7359_),
    .Y(_7361_)
);

OAI21X1 _17211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6899_),
    .B(_6898_),
    .C(_6897_),
    .Y(_6901_)
);

AOI21X1 _22288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .B(_556_),
    .C(_369_),
    .Y(_557_)
);

FILL SFILL33800x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8678_),
    .B(_8675_),
    .C(_8677_),
    .Y(_8682_)
);

OR2X2 _18416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8217_),
    .B(_8221_),
    .Y(_8222_)
);

OAI21X1 _13971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3349_),
    .B(_3345_),
    .C(_3311_),
    .Y(_3351_)
);

NOR3X1 _13551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2878_),
    .B(_2887_),
    .C(_2888_),
    .Y(_2891_)
);

NAND2X1 _13131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_11_bF$buf1),
    .Y(_2432_)
);

FILL SFILL13800x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_16_bF$buf2),
    .Y(_4210_)
);

OAI21X1 _14336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3736_),
    .B(_3742_),
    .C(_3744_),
    .Y(_3751_)
);

DFFPOSX1 _24014_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[4]),
    .CLK(clk_bF$buf10),
    .D(a[4])
);

FILL SFILL18840x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10443_),
    .B(_10435_),
    .Y(_10807_)
);

INVX2 _20354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10345_),
    .Y(_10346_)
);

AND2X2 _16902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5842_),
    .B(_6223_),
    .Y(_6562_)
);

AOI21X1 _19794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9732_),
    .B(_9731_),
    .C(_9724_),
    .Y(_9733_)
);

OAI21X1 _19374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9271_),
    .B(_8888_),
    .C(_9234_),
    .Y(_9272_)
);

NOR3X1 _21979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11838_),
    .B(_11840_),
    .C(_11831_),
    .Y(_219_)
);

NOR3X1 _21559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11650_),
    .B(_11654_),
    .C(_11653_),
    .Y(_11666_)
);

OAI21X1 _21139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11202_),
    .B(_11203_),
    .C(_11168_),
    .Y(_11207_)
);

AND2X2 _12822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_429_),
    .Y(_451_)
);

AND2X2 _12402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_7689_),
    .Y(_7755_)
);

AOI21X1 _22920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1236_),
    .B(_1237_),
    .C(_1101_),
    .Y(_1249_)
);

AOI21X1 _22500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_782_),
    .B(_784_),
    .C(_781_),
    .Y(_789_)
);

OAI21X1 _15294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4501_),
    .B(_4524_),
    .C(_4515_),
    .Y(_4800_)
);

FILL SFILL48920x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2757_),
    .B(_2947_),
    .C(_2952_),
    .Y(_2953_)
);

OR2X2 _23705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2102_),
    .B(_2056_),
    .Y(_2104_)
);

OAI21X1 _16499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5831_),
    .B(_5824_),
    .C(_5833_),
    .Y(_6119_)
);

NOR2X1 _16079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5284_),
    .B(_5656_),
    .Y(_5659_)
);

NOR3X1 _17860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7180_),
    .B(_7181_),
    .C(_7179_),
    .Y(_7612_)
);

AOI21X1 _17440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7147_),
    .B(_7146_),
    .C(_7145_),
    .Y(_7152_)
);

OAI21X1 _17020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6690_),
    .B(_6689_),
    .C(_6680_),
    .Y(_6691_)
);

NAND3X1 _22097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_340_),
    .B(_347_),
    .C(_293_),
    .Y(_348_)
);

AOI21X1 _18645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8450_),
    .B(_8451_),
    .C(_8074_),
    .Y(_8472_)
);

OAI21X1 _18225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7875_),
    .B(_7874_),
    .C(_7783_),
    .Y(_8013_)
);

FILL SFILL59080x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf3),
    .B(areg_16_bF$buf0),
    .Y(_3141_)
);

AOI21X1 _13360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2674_),
    .B(_2671_),
    .C(_2662_),
    .Y(_2682_)
);

NAND2X1 _14985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_13_bF$buf2),
    .Y(_4460_)
);

NAND3X1 _14565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3989_),
    .B(_3946_),
    .C(_3983_),
    .Y(_4002_)
);

INVX1 _14145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3540_),
    .Y(_3541_)
);

FILL SFILL3560x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10592_),
    .B(_10593_),
    .C(_10591_),
    .Y(_10598_)
);

XNOR2X1 _20163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10115_),
    .B(_10111_),
    .Y(_10137_)
);

FILL SFILL28920x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6347_),
    .B(_6346_),
    .C(_6345_),
    .Y(_6353_)
);

OAI21X1 _19183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9057_),
    .B(_9058_),
    .C(_9062_),
    .Y(_9063_)
);

OAI21X1 _21788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8_),
    .B(_2_),
    .C(_11894_),
    .Y(_9_)
);

AOI21X1 _21368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11457_),
    .B(_11456_),
    .C(_11455_),
    .Y(_11458_)
);

INVX2 _17916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7672_),
    .Y(_7673_)
);

INVX1 _12631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10035_),
    .Y(_10266_)
);

OAI21X1 _12211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5387_),
    .B(_5398_),
    .C(_5354_),
    .Y(_5661_)
);

AOI21X1 _13836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3195_),
    .B(_3203_),
    .C(_3047_),
    .Y(_3204_)
);

NAND3X1 _13416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2548_),
    .B(_2740_),
    .C(_2743_),
    .Y(_2744_)
);

BUFX2 _23934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[52]),
    .Y(y[52])
);

XNOR2X1 _23514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1891_),
    .Y(_1895_)
);

FILL SFILL18840x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _18874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8700_),
    .B(_8696_),
    .Y(_8724_)
);

NAND3X1 _18454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8223_),
    .B(_8256_),
    .C(_8259_),
    .Y(_8264_)
);

NOR2X1 _18034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7355_),
    .B(_7802_),
    .Y(_7803_)
);

NAND3X1 _20639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10657_),
    .B(_10658_),
    .C(_10656_),
    .Y(_10659_)
);

NOR3X1 _20219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10194_),
    .B(_10195_),
    .C(_10197_),
    .Y(_10198_)
);

NOR3X1 _19659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9188_),
    .B(_9196_),
    .C(_9198_),
    .Y(_9585_)
);

XNOR2X1 _19239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9101_),
    .B(_9098_),
    .Y(_9124_)
);

NOR2X1 _14794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3972_),
    .B(_4250_),
    .Y(_4251_)
);

AND2X2 _14374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3528_),
    .B(_3790_),
    .Y(_3792_)
);

DFFPOSX1 _24052_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[10]),
    .CLK(clk_bF$buf4),
    .D(b[10])
);

FILL SFILL69080x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(_5571_),
    .C(_5554_),
    .Y(_5572_)
);

INVX2 _15579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5110_),
    .Y(_5111_)
);

OAI21X1 _15159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4650_),
    .B(_4349_),
    .C(_4618_),
    .Y(_4651_)
);

OAI21X1 _20392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10384_),
    .B(_10383_),
    .C(_10382_),
    .Y(_10388_)
);

NAND2X1 _16940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6238_),
    .B(_6244_),
    .Y(_6603_)
);

AND2X2 _16520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_18_bF$buf0),
    .Y(_6142_)
);

OAI21X1 _16100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5315__bF$buf0),
    .C(_5681_),
    .Y(_5682_)
);

NAND3X1 _21597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11604_),
    .B(_11703_),
    .C(_11707_),
    .Y(_11708_)
);

NAND2X1 _21177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10927_),
    .B(_10932_),
    .Y(_11249_)
);

NAND3X1 _17725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7456_),
    .B(_7463_),
    .C(_7442_),
    .Y(_7464_)
);

NAND3X1 _17305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6997_),
    .B(_7003_),
    .C(_7002_),
    .Y(_7004_)
);

FILL SFILL59080x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11154_),
    .B(_11143_),
    .C(_11121_),
    .Y(_867_)
);

OAI21X1 _12440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8150_),
    .B(_8161_),
    .C(_8139_),
    .Y(_8172_)
);

NAND2X1 _12020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_5_bF$buf1),
    .Y(_3569_)
);

FILL SFILL3640x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _13645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2993_),
    .Y(_2994_)
);

NAND2X1 _13225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2532_),
    .B(_2533_),
    .Y(_2535_)
);

XNOR2X1 _23743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .B(_2135_),
    .Y(_2145_)
);

OAI21X1 _23323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1687_),
    .B(_1686_),
    .C(_1666_),
    .Y(_1688_)
);

FILL SFILL49080x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28920x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8487_),
    .B(_8512_),
    .C(_8513_),
    .Y(_8514_)
);

NAND3X1 _18263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7659_),
    .B(_8048_),
    .C(_8051_),
    .Y(_8055_)
);

FILL SFILL49000x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10574_),
    .B(_10579_),
    .Y(_10910_)
);

NAND3X1 _20448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10447_),
    .B(_10448_),
    .C(_10443_),
    .Y(_10449_)
);

INVX1 _20028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9987_),
    .Y(_9988_)
);

NAND3X1 _19888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9791_),
    .B(_9824_),
    .C(_9827_),
    .Y(_9836_)
);

OAI21X1 _19468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9090_),
    .B(_9091_),
    .C(_9088_),
    .Y(_9375_)
);

OAI21X1 _19048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf2),
    .B(_5668__bF$buf4),
    .C(_8901_),
    .Y(_8914_)
);

OAI21X1 _14183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3579_),
    .B(_3581_),
    .C(_3582_),
    .Y(_3583_)
);

FILL SFILL18920x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_),
    .B(_943_),
    .C(_856_),
    .Y(_1478_)
);

NOR3X1 _15388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4896_),
    .B(_4897_),
    .C(_4894_),
    .Y(_4903_)
);

FILL SFILL39000x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert130 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(breg_4_bF$buf0)
);

BUFX2 BUFX2_insert131 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf4)
);

BUFX2 BUFX2_insert132 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf3)
);

BUFX2 BUFX2_insert133 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf2)
);

AND2X2 _17954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7278_),
    .B(_7713_),
    .Y(_7715_)
);

BUFX2 BUFX2_insert134 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf1)
);

BUFX2 BUFX2_insert135 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(breg_13_bF$buf0)
);

NOR3X1 _17534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7253_),
    .B(_7248_),
    .C(_7252_),
    .Y(_7254_)
);

BUFX2 BUFX2_insert136 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921_),
    .Y(_5921__bF$buf3)
);

AOI21X1 _17114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6789_),
    .B(_6790_),
    .C(_6788_),
    .Y(_6795_)
);

BUFX2 BUFX2_insert137 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921_),
    .Y(_5921__bF$buf2)
);

BUFX2 BUFX2_insert138 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921_),
    .Y(_5921__bF$buf1)
);

BUFX2 BUFX2_insert139 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5921_),
    .Y(_5921__bF$buf0)
);

NAND3X1 _18739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8552_),
    .B(_8557_),
    .C(_8564_),
    .Y(_8575_)
);

NOR3X1 _18319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8112_),
    .B(_8113_),
    .C(_8114_),
    .Y(_8115_)
);

OAI21X1 _13874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3244_),
    .B(_2985_),
    .C(_3219_),
    .Y(_3245_)
);

NAND2X1 _13454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2784_),
    .B(_2783_),
    .Y(_2785_)
);

DFFPOSX1 _23972_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[26]),
    .CLK(clk_bF$buf7),
    .D(_0_[26])
);

AOI21X1 _13034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2324_),
    .C(_2323_),
    .Y(_2329_)
);

AOI21X1 _23552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1937_),
    .C(_1872_),
    .Y(_1938_)
);

NOR3X1 _23132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(_1471_),
    .C(_1475_),
    .Y(_1480_)
);

NAND2X1 _14659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4101_),
    .B(_4102_),
    .Y(_4103_)
);

AND2X2 _14239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_14_bF$buf4),
    .Y(_3644_)
);

FILL SFILL3720x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5132_),
    .B(_5133_),
    .C(_5131_),
    .Y(_5134_)
);

NOR2X1 _18492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7903_),
    .B(_8305_),
    .Y(_8306_)
);

NAND3X1 _18072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7827_),
    .B(_7830_),
    .C(_7840_),
    .Y(_7845_)
);

INVX1 _20677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10699_),
    .Y(_10700_)
);

XNOR2X1 _20257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10213_),
    .B(_10239_),
    .Y(_10240_)
);

NAND2X1 _16805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_22_bF$buf1),
    .Y(_6455_)
);

INVX1 _11940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2683_),
    .Y(_2694_)
);

NAND3X1 _19697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9270_),
    .B(_9610_),
    .C(_9617_),
    .Y(_9627_)
);

AOI21X1 _19277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9160_),
    .B(_9165_),
    .C(_9143_),
    .Y(_9166_)
);

FILL SFILL43880x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11242_),
    .B(_11286_),
    .C(_10024_),
    .Y(_11297_)
);

OAI21X1 _12305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6670_),
    .B(_6681_),
    .C(_6659_),
    .Y(_6692_)
);

NOR2X1 _22823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4541__bF$buf2),
    .B(_5676_),
    .Y(_1143_)
);

AOI21X1 _22403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_681_),
    .B(_682_),
    .C(_498_),
    .Y(_683_)
);

NAND3X1 _15197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4687_),
    .B(_4692_),
    .C(_4691_),
    .Y(_4693_)
);

OAI21X1 _23608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1829_),
    .B(_1924_),
    .C(_1927_),
    .Y(_1998_)
);

FILL SFILL49080x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7487_),
    .B(_7500_),
    .C(_7505_),
    .Y(_7506_)
);

XNOR2X1 _17343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7022_),
    .B(_7045_),
    .Y(_7046_)
);

FILL SFILL33880x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18600x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8688_),
    .B(_8685_),
    .C(_8681_),
    .Y(_8827_)
);

OAI21X1 _18548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8365_),
    .B(_8366_),
    .C(_8363_),
    .Y(_8367_)
);

OAI21X1 _18128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7905_),
    .B(_7904_),
    .C(_7889_),
    .Y(_7906_)
);

NAND3X1 _13683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3034_),
    .B(_3035_),
    .C(_3029_),
    .Y(_3036_)
);

XNOR2X1 _13263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2575_),
    .B(_2572_),
    .Y(_2576_)
);

NOR2X1 _23781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2170_),
    .Y(_2186_)
);

OAI21X1 _23361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1725_),
    .C(_1693_),
    .Y(_1730_)
);

NOR2X1 _14888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4353_),
    .B(_4095_),
    .Y(_4354_)
);

INVX1 _14468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3869_),
    .Y(_3895_)
);

FILL SFILL23800x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3430_),
    .B(_3434_),
    .C(_3358_),
    .Y(_3435_)
);

FILL SFILL23880x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8840x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54280x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53960x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53880x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _20486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10467_),
    .B(_10464_),
    .Y(_10491_)
);

NAND3X1 _20066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10004_),
    .B(_10028_),
    .C(_10029_),
    .Y(_10030_)
);

XNOR2X1 _16614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6224_),
    .B(_6245_),
    .Y(_6246_)
);

OAI21X1 _19086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf2),
    .B(_3781__bF$buf1),
    .C(_8541_),
    .Y(_8956_)
);

FILL SFILL8760x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _17819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7138_),
    .B(_7139_),
    .C(_7137_),
    .Y(_7567_)
);

OAI21X1 _12954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_385_),
    .C(_834_),
    .Y(_1902_)
);

NOR3X1 _12534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9049_),
    .B(_9148_),
    .C(_9159_),
    .Y(_9203_)
);

OAI21X1 _22632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9263_),
    .B(_10685_),
    .C(_933_),
    .Y(_934_)
);

AOI21X1 _12114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3547_),
    .B(_3745_),
    .C(_3810_),
    .Y(_4599_)
);

OAI21X1 _22212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_464_),
    .C(_468_),
    .Y(_475_)
);

FILL SFILL74440x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_2845_),
    .Y(_3097_)
);

NAND2X1 _13319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2634_),
    .Y(_2637_)
);

AND2X2 _23837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2186_),
    .B(_2231_),
    .Y(_2245_)
);

NOR2X1 _23417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1789_),
    .Y(_1790_)
);

FILL SFILL43960x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert510 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .Y(_3961__bF$buf2)
);

BUFX2 BUFX2_insert511 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .Y(_3961__bF$buf1)
);

BUFX2 BUFX2_insert512 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961_),
    .Y(_3961__bF$buf0)
);

BUFX2 BUFX2_insert513 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .Y(_3253__bF$buf3)
);

AOI21X1 _17992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7756_),
    .B(_7754_),
    .C(_7746_),
    .Y(_7757_)
);

BUFX2 BUFX2_insert514 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .Y(_3253__bF$buf2)
);

BUFX2 BUFX2_insert515 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .Y(_3253__bF$buf1)
);

INVX1 _17572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7275_),
    .Y(_7296_)
);

INVX1 _17152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6831_),
    .Y(_6836_)
);

BUFX2 BUFX2_insert516 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253_),
    .Y(_3253__bF$buf0)
);

BUFX2 BUFX2_insert517 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .Y(_3958__bF$buf3)
);

BUFX2 BUFX2_insert518 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .Y(_3958__bF$buf2)
);

BUFX2 BUFX2_insert519 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958_),
    .Y(_3958__bF$buf1)
);

FILL SFILL23960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8614_),
    .B(_8612_),
    .Y(_8617_)
);

AND2X2 _18357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7730_),
    .B(_7724_),
    .Y(_8157_)
);

OAI21X1 _13492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2826_),
    .B(_2646_),
    .C(_2637_),
    .Y(_2827_)
);

FILL FILL74120x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .B(_2366_),
    .Y(_2367_)
);

OAI21X1 _23590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1975_),
    .B(_488_),
    .C(_1977_),
    .Y(_1978_)
);

OAI21X1 _23170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_1267_),
    .C(_1376_),
    .Y(_1521_)
);

FILL SFILL64360x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .Y(_136_)
);

OAI21X1 _14697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4143_),
    .B(_4142_),
    .C(_4144_),
    .Y(_4145_)
);

NAND2X1 _14277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3400_),
    .B(_3685_),
    .Y(_3686_)
);

OAI21X1 _20295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10280_),
    .B(_10281_),
    .C(_10279_),
    .Y(_10282_)
);

AOI21X1 _16843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6130_),
    .B(_6214_),
    .C(_6211_),
    .Y(_6497_)
);

NAND2X1 _16423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(_5659_),
    .Y(_6036_)
);

NAND3X1 _16003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5573_),
    .B(_5576_),
    .C(_5575_),
    .Y(_5577_)
);

AND2X2 _17628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_19_bF$buf1),
    .Y(_7357_)
);

AOI21X1 _17208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6481_),
    .B(_6484_),
    .C(_6896_),
    .Y(_6897_)
);

NAND2X1 _12763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg_13_bF$buf0),
    .Y(_11712_)
);

NAND3X1 _12343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5914_),
    .B(_7098_),
    .C(_7054_),
    .Y(_7109_)
);

AND2X2 _22861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(_1010_),
    .Y(_1185_)
);

OAI21X1 _22441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_723_),
    .B(_495_),
    .C(_698_),
    .Y(_725_)
);

OAI21X1 _22021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf2),
    .B(_6050__bF$buf3),
    .C(_263_),
    .Y(_265_)
);

FILL SFILL18520x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59080x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8920x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3338_),
    .B(_3335_),
    .C(_3320_),
    .Y(_3347_)
);

FILL SFILL23800x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _13548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2881_),
    .B(_2882_),
    .Y(_2888_)
);

OAI21X1 _13128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_6582__bF$buf3),
    .C(_1936_),
    .Y(_2428_)
);

OR2X2 _23646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2027_),
    .B(_2039_),
    .Y(_2040_)
);

OAI21X1 _23226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686__bF$buf1),
    .B(_5676_),
    .C(_1580_),
    .Y(_1581_)
);

NOR3X1 _17381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7081_),
    .B(_7082_),
    .C(_7080_),
    .Y(_7088_)
);

OAI21X1 _18586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8400_),
    .B(_8407_),
    .C(_8281_),
    .Y(_8408_)
);

OAI21X1 _18166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7945_),
    .B(_7946_),
    .C(_7947_),
    .Y(_7948_)
);

FILL SFILL74120x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11832_),
    .B(_11834_),
    .Y(_11835_)
);

OAI21X1 _14086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3472_),
    .C(_3248_),
    .Y(_3477_)
);

INVX2 _12819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_407_),
    .Y(_418_)
);

AOI21X1 _22917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_946_),
    .B(_1080_),
    .C(_1245_),
    .Y(_1246_)
);

FILL SFILL8680x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6282_),
    .B(_6283_),
    .C(_6279_),
    .Y(_6288_)
);

AOI21X1 _16232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5465_),
    .B(_5507_),
    .C(_5504_),
    .Y(_5828_)
);

FILL SFILL19000x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7589_),
    .B(_7596_),
    .C(_7599_),
    .Y(_7609_)
);

NAND3X1 _17437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7141_),
    .B(_7148_),
    .C(_7064_),
    .Y(_7149_)
);

NAND3X1 _17017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6682_),
    .B(_6687_),
    .C(_6685_),
    .Y(_6688_)
);

INVX8 _12992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf4),
    .Y(_2287_)
);

NAND3X1 _12572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9477_),
    .B(_9521_),
    .C(_9554_),
    .Y(_9620_)
);

NOR2X1 _12152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_4258__bF$buf3),
    .Y(_5014_)
);

NAND2X1 _22670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_972_),
    .Y(_975_)
);

INVX1 _22250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_509_),
    .Y(_515_)
);

OAI21X1 _13777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3137_),
    .B(_3136_),
    .C(_3135_),
    .Y(_3138_)
);

NAND3X1 _13357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2675_),
    .B(_2659_),
    .C(_2678_),
    .Y(_2679_)
);

OAI21X1 _23875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2284_),
    .C(_2272_),
    .Y(_2285_)
);

NOR2X1 _23455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1823_),
    .Y(_1832_)
);

NAND3X1 _23035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(_1372_),
    .C(_1373_),
    .Y(_1374_)
);

OAI21X1 _17190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6868_),
    .B(_6869_),
    .C(_6865_),
    .Y(_6877_)
);

AOI21X1 _15923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5479_),
    .B(_5477_),
    .C(_5474_),
    .Y(_5489_)
);

OAI21X1 _15503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf0),
    .B(_3529__bF$buf3),
    .C(_4694_),
    .Y(_5028_)
);

OAI21X1 _18395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf3),
    .B(_3253__bF$buf1),
    .C(_8198_),
    .Y(_8199_)
);

NAND3X1 _16708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6265_),
    .B(_6342_),
    .C(_6348_),
    .Y(_6349_)
);

INVX2 _21941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_176_),
    .Y(_178_)
);

AOI21X1 _21521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11335_),
    .B(_11339_),
    .C(_11342_),
    .Y(_11626_)
);

AOI21X1 _21101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11164_),
    .B(_11163_),
    .C(_11162_),
    .Y(_11166_)
);

FILL SFILL44040x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10101_),
    .B(_10232_),
    .Y(_10233_)
);

NAND3X1 _12208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4094_),
    .B(_5607_),
    .C(_5618_),
    .Y(_5629_)
);

NOR2X1 _22726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5369_),
    .B(_6300__bF$buf2),
    .Y(_1037_)
);

AOI21X1 _22306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_397_),
    .C(_387_),
    .Y(_577_)
);

FILL SFILL8520x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6537_),
    .B(_6530_),
    .C(_6517_),
    .Y(_6539_)
);

NOR2X1 _16461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5688_),
    .B(_5750_),
    .Y(_6077_)
);

NAND3X1 _16041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5599_),
    .B(_5605_),
    .C(_5609_),
    .Y(_5619_)
);

AOI21X1 _17666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7045_),
    .B(_7398_),
    .C(_7019_),
    .Y(_7399_)
);

FILL SFILL74120x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _17246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6937_),
    .B(_6938_),
    .Y(_6939_)
);

NAND2X1 _12381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7393_),
    .B(_7459_),
    .Y(_7525_)
);

NOR2X1 _13586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2929_),
    .B(_2928_),
    .Y(_2930_)
);

NAND3X1 _13166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2467_),
    .C(_2458_),
    .Y(_2470_)
);

XOR2X1 _23684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_2068_),
    .Y(_2081_)
);

AOI21X1 _23264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1611_),
    .B(_1606_),
    .C(_1555_),
    .Y(_1624_)
);

NAND3X1 _19812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9750_),
    .B(_9752_),
    .C(_9749_),
    .Y(_9753_)
);

FILL SFILL64120x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24049_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[7]),
    .CLK(clk_bF$buf0),
    .D(b[7])
);

INVX2 _15732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4967_),
    .Y(_5280_)
);

AND2X2 _15312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_17_bF$buf5),
    .Y(_4820_)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[21]),
    .Y(areg_21_bF$buf0)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf5)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf4)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf3)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf2)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf1)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[18]),
    .Y(areg_18_bF$buf0)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf4)
);

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf3)
);

BUFX2 BUFX2_insert49 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf2)
);

NOR3X1 _20389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10369_),
    .B(_10355_),
    .C(_10376_),
    .Y(_10384_)
);

NAND2X1 _16937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6599_),
    .B(_6595_),
    .Y(_6600_)
);

NAND2X1 _16517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf2),
    .B(breg_18_bF$buf0),
    .Y(_6139_)
);

NAND2X1 _21750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11313_),
    .B(_11874_),
    .Y(_11875_)
);

AOI21X1 _21330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11400_),
    .B(_11404_),
    .C(_11370_),
    .Y(_11416_)
);

FILL SFILL54120x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_396_),
    .B(_680_),
    .C(_713_),
    .Y(_834_)
);

AOI21X1 _12437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6099_),
    .B(_6900_),
    .C(_6922_),
    .Y(_8139_)
);

XNOR2X1 _22955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(_1273_),
    .Y(_1287_)
);

XOR2X1 _12017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3514_),
    .B(_3525_),
    .Y(_3536_)
);

NAND3X1 _22535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_662_),
    .B(_827_),
    .C(_822_),
    .Y(_828_)
);

NOR2X1 _22115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf3),
    .B(_5369_),
    .Y(_367_)
);

FILL SFILL54040x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6322_),
    .B(_6328_),
    .C(_6306_),
    .Y(_6329_)
);

NAND3X1 _16270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5860_),
    .B(_5853_),
    .C(_5857_),
    .Y(_5869_)
);

FILL SFILL18680x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44520x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _17895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .B(_7644_),
    .Y(_7650_)
);

NAND3X1 _17475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7189_),
    .B(_7187_),
    .C(_7188_),
    .Y(_7190_)
);

OAI21X1 _17055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6671_),
    .B(_6666_),
    .C(_6673_),
    .Y(_6730_)
);

NOR2X1 _12190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf3),
    .B(_5420__bF$buf1),
    .Y(_5431_)
);

AOI21X1 _20601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10274_),
    .B(_10205_),
    .C(_10280_),
    .Y(_10618_)
);

FILL SFILL44040x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2576_),
    .B(_2719_),
    .C(_2720_),
    .Y(_2721_)
);

AOI21X1 _23493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1846_),
    .C(_1844_),
    .Y(_1873_)
);

OAI21X1 _23073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(_1275_),
    .C(_1280_),
    .Y(_1415_)
);

NAND3X1 _19621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9533_),
    .B(_9540_),
    .C(_9542_),
    .Y(_9544_)
);

AOI21X1 _19201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9080_),
    .B(_9081_),
    .C(_9079_),
    .Y(_9082_)
);

NAND2X1 _21806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf2),
    .B(breg_26_bF$buf4),
    .Y(_29_)
);

AOI21X1 _15961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5524_),
    .B(_5525_),
    .C(_5523_),
    .Y(_5531_)
);

FILL SFILL69240x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5051_),
    .B(_5054_),
    .C(_5057_),
    .Y(_5070_)
);

AOI21X1 _15121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4592_),
    .B(_4597_),
    .C(_4444_),
    .Y(_4611_)
);

NAND3X1 _20198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10165_),
    .B(_10152_),
    .C(_10155_),
    .Y(_10175_)
);

NAND3X1 _16746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6388_),
    .B(_6390_),
    .C(_6389_),
    .Y(_6391_)
);

INVX2 _16326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5930_),
    .Y(_5931_)
);

FILL SFILL69160x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10441_),
    .Y(_10650_)
);

INVX8 _12246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf3),
    .Y(_6044_)
);

NOR3X1 _22764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1076_),
    .B(_1077_),
    .C(_1078_),
    .Y(_1079_)
);

INVX2 _22344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_618_),
    .Y(_619_)
);

DFFPOSX1 _23969_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[23]),
    .CLK(clk_bF$buf2),
    .D(_0_[23])
);

FILL SFILL64120x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_1933_),
    .C(_1829_),
    .Y(_1934_)
);

OAI21X1 _23129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1474_),
    .B(_1475_),
    .C(_1471_),
    .Y(_1476_)
);

OAI21X1 _14812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4271_),
    .B(_4269_),
    .C(_4268_),
    .Y(_4272_)
);

NOR2X1 _17284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6561_),
    .B(_6974_),
    .Y(_6981_)
);

FILL SFILL59160x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10860_),
    .B(_10867_),
    .C(_10864_),
    .Y(_10868_)
);

AND2X2 _20410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10056_),
    .B(_10114_),
    .Y(_10407_)
);

AOI21X1 _18489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7895_),
    .B(_7897_),
    .C(_7904_),
    .Y(_8302_)
);

OAI21X1 _18069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7836_),
    .B(_7837_),
    .C(_7840_),
    .Y(_7841_)
);

NAND2X1 _19850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf1),
    .B(areg_20_bF$buf0),
    .Y(_9794_)
);

NAND2X1 _19430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_22_bF$buf0),
    .Y(_9333_)
);

NAND3X1 _19010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8475_),
    .B(_8864_),
    .C(_8858_),
    .Y(_8873_)
);

INVX8 _11937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .Y(_2661_)
);

NAND2X1 _21615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_20_bF$buf4),
    .B(areg_23_bF$buf0),
    .Y(_11728_)
);

OAI21X1 _15770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf0),
    .B(_5315__bF$buf1),
    .C(_5312_),
    .Y(_5320_)
);

NAND3X1 _15350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4856_),
    .B(_4860_),
    .C(_4858_),
    .Y(_4861_)
);

NOR3X1 _16975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6639_),
    .B(_6640_),
    .C(_6641_),
    .Y(_6642_)
);

AOI21X1 _16555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6173_),
    .B(_6174_),
    .C(_6166_),
    .Y(_6181_)
);

AOI21X1 _16135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4980_),
    .B(_5346_),
    .C(_5720_),
    .Y(_5721_)
);

FILL SFILL54200x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8391_),
    .B(_1239_),
    .C(_9904_),
    .Y(_1250_)
);

INVX4 _12475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf3),
    .Y(_8555_)
);

AOI21X1 _22993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1318_),
    .B(_1316_),
    .C(_1298_),
    .Y(_1328_)
);

AOI21X1 _12055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3909_),
    .B(_3942_),
    .C(_3372_),
    .Y(_3953_)
);

NOR2X1 _22573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .B(_868_),
    .Y(_870_)
);

NOR3X1 _22153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_408_),
    .C(_406_),
    .Y(_410_)
);

NOR2X1 _18701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8531_),
    .B(_8532_),
    .Y(_8534_)
);

XNOR2X1 _23778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2181_),
    .B(_2177_),
    .Y(_2182_)
);

OAI21X1 _23358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .B(_1725_),
    .C(_1692_),
    .Y(_1726_)
);

AND2X2 _19906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9509_),
    .B(_9502_),
    .Y(_9856_)
);

FILL SFILL69240x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3855_),
    .B(_3860_),
    .Y(_4062_)
);

AND2X2 _14201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_11_bF$buf0),
    .Y(_3602_)
);

NAND3X1 _17093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6424_),
    .B(_6507_),
    .C(_6506_),
    .Y(_6772_)
);

AND2X2 _15826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg_19_bF$buf1),
    .Y(_5382_)
);

NAND3X1 _15406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4676_),
    .B(_4915_),
    .C(_4922_),
    .Y(_4923_)
);

OAI22X1 _18298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf4),
    .B(_6050__bF$buf0),
    .C(_3646__bF$buf0),
    .D(_5668__bF$buf3),
    .Y(_8092_)
);

FILL SFILL59240x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11648_),
    .B(_11684_),
    .C(_70_),
    .Y(_71_)
);

NAND3X1 _21424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11514_),
    .B(_11515_),
    .C(_11513_),
    .Y(_11520_)
);

NAND2X1 _21004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10758_),
    .B(_10766_),
    .Y(_11059_)
);

FILL SFILL64360x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3800x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64040x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _22629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10680_),
    .Y(_930_)
);

NAND3X1 _22209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(_470_),
    .C(_468_),
    .Y(_471_)
);

OAI21X1 _16784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6051_),
    .B(_6430_),
    .C(_6431_),
    .Y(_6432_)
);

AOI21X1 _16364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5954_),
    .B(_5960_),
    .C(_5912_),
    .Y(_5973_)
);

BUFX2 BUFX2_insert480 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf1)
);

BUFX2 BUFX2_insert481 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(breg_5_bF$buf0)
);

BUFX2 BUFX2_insert482 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf3)
);

BUFX2 BUFX2_insert483 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf2)
);

BUFX2 BUFX2_insert484 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf1)
);

AOI21X1 _17989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7274_),
    .B(_7308_),
    .C(_7752_),
    .Y(_7753_)
);

BUFX2 BUFX2_insert485 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(breg_14_bF$buf0)
);

AOI21X1 _17569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6926_),
    .B(_7291_),
    .C(_6928_),
    .Y(_7292_)
);

BUFX2 BUFX2_insert486 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(breg_2_bF$buf4)
);

NOR3X1 _17149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6819_),
    .B(_6831_),
    .C(_6827_),
    .Y(_6832_)
);

BUFX2 BUFX2_insert487 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(breg_2_bF$buf3)
);

BUFX2 BUFX2_insert488 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(breg_2_bF$buf2)
);

BUFX2 BUFX2_insert489 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .Y(breg_2_bF$buf1)
);

FILL SFILL33880x50 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6450_),
    .Y(_6461_)
);

OAI21X1 _22382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_660_),
    .B(_657_),
    .C(_656_),
    .Y(_661_)
);

OAI21X1 _18930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8767_),
    .B(_8768_),
    .C(_8744_),
    .Y(_8785_)
);

AND2X2 _18510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7916_),
    .B(_7911_),
    .Y(_8325_)
);

FILL SFILL33960x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2804_),
    .B(_2810_),
    .Y(_2823_)
);

NOR2X1 _13069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_2362__bF$buf0),
    .Y(_2363_)
);

INVX1 _23587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_920_),
    .Y(_1975_)
);

NOR3X1 _23167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1364_),
    .B(_1504_),
    .C(_1508_),
    .Y(_1518_)
);

NOR2X1 _19715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf0),
    .B(_7225__bF$buf3),
    .Y(_9646_)
);

FILL SFILL18760x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4295_),
    .B(_4300_),
    .C(_4152_),
    .Y(_4313_)
);

OAI21X1 _14430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3633_),
    .B(_3634_),
    .C(_3631_),
    .Y(_3853_)
);

AOI21X1 _14010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3389_),
    .B(_3391_),
    .C(_3392_),
    .Y(_3393_)
);

NAND3X1 _15635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5152_),
    .B(_5166_),
    .C(_5172_),
    .Y(_5173_)
);

INVX1 _15215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4712_),
    .Y(_4713_)
);

FILL SFILL23960x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _11975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf4),
    .B(areg_2_bF$buf2),
    .C(breg_1_bF$buf3),
    .D(areg_1_bF$buf3),
    .Y(_3077_)
);

NAND3X1 _21653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11763_),
    .B(_11769_),
    .C(_11766_),
    .Y(_11770_)
);

NAND3X1 _21233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11005_),
    .B(_11304_),
    .C(_11305_),
    .Y(_11310_)
);

FILL SFILL69320x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1172_),
    .C(_1132_),
    .Y(_1181_)
);

AOI21X1 _22438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_720_),
    .C(_709_),
    .Y(_721_)
);

AND2X2 _22018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf2),
    .B(breg_27_bF$buf4),
    .Y(_261_)
);

AND2X2 _13701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2796_),
    .B(_3053_),
    .Y(_3056_)
);

NAND2X1 _16593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_16_bF$buf4),
    .Y(_6223_)
);

OAI22X1 _16173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf3),
    .B(_3253__bF$buf3),
    .C(_6582__bF$buf2),
    .D(_3529__bF$buf1),
    .Y(_5763_)
);

NOR3X1 _14906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4370_),
    .B(_4372_),
    .C(_4373_),
    .Y(_4374_)
);

FILL SFILL29000x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7534_),
    .B(_7532_),
    .C(_7530_),
    .Y(_7544_)
);

NAND3X1 _17378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7066_),
    .B(_7079_),
    .C(_7083_),
    .Y(_7084_)
);

INVX1 _12093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4357_),
    .Y(_4368_)
);

AOI21X1 _22191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_193_),
    .C(_209_),
    .Y(_452_)
);

FILL SFILL8600x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10964_),
    .B(_10971_),
    .C(_10697_),
    .Y(_10972_)
);

NAND2X1 _20504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_26_bF$buf4),
    .Y(_10511_)
);

AOI21X1 _13298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2608_),
    .B(_2607_),
    .C(_2606_),
    .Y(_2613_)
);

NAND2X1 _23396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .B(_1763_),
    .Y(_1768_)
);

NAND2X1 _19944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9502_),
    .B(_9509_),
    .Y(_9897_)
);

OAI21X1 _19524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_3961__bF$buf0),
    .C(_9426_),
    .Y(_9437_)
);

NAND3X1 _19104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8959_),
    .B(_8964_),
    .C(_8971_),
    .Y(_8976_)
);

NOR3X1 _21709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11830_),
    .B(_11827_),
    .C(_11715_),
    .Y(_11831_)
);

FILL FILL74200x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5416_),
    .B(_5417_),
    .C(_5408_),
    .Y(_5424_)
);

OAI21X1 _15444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4962_),
    .B(_4961_),
    .C(_4957_),
    .Y(_4963_)
);

AND2X2 _15024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_17_bF$buf5),
    .Y(_4504_)
);

FILL SFILL33640x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _16649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6283_),
    .B(_6279_),
    .C(_6282_),
    .Y(_6284_)
);

AOI21X1 _16229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5822_),
    .C(_5823_),
    .Y(_5824_)
);

OAI21X1 _21882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_6686__bF$buf2),
    .C(_11729_),
    .Y(_113_)
);

AOI21X1 _21462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11547_),
    .B(_11548_),
    .C(_11258_),
    .Y(_11562_)
);

AOI21X1 _21042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11083_),
    .B(_11087_),
    .C(_11090_),
    .Y(_11101_)
);

FILL SFILL13880x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2259_),
    .Y(_2270_)
);

OAI21X1 _12569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9565_),
    .B(_9576_),
    .C(_9554_),
    .Y(_9587_)
);

OAI21X1 _12149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4818_),
    .B(_3449_),
    .C(_4697_),
    .Y(_4981_)
);

XOR2X1 _22667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_969_),
    .B(_957_),
    .Y(_972_)
);

NAND2X1 _22247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf1),
    .B(breg_27_bF$buf4),
    .Y(_512_)
);

OAI21X1 _13930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3299_),
    .B(_3300_),
    .C(_3297_),
    .Y(_3306_)
);

XOR2X1 _13510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2631_),
    .B(_2845_),
    .Y(_2846_)
);

INVX2 _14715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4164_),
    .Y(_4165_)
);

NAND3X1 _17187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6850_),
    .B(_6873_),
    .C(_6866_),
    .Y(_6874_)
);

FILL SFILL23960x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10406_),
    .B(_10466_),
    .Y(_10762_)
);

AOI21X1 _20313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10296_),
    .B(_10295_),
    .C(_10294_),
    .Y(_10302_)
);

OAI21X1 _19753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9355_),
    .B(_9358_),
    .C(_9349_),
    .Y(_9688_)
);

NOR3X1 _19333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8825_),
    .B(_8832_),
    .C(_8835_),
    .Y(_9228_)
);

FILL SFILL69320x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_160_),
    .C(_11818_),
    .Y(_174_)
);

NOR2X1 _21518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11613_),
    .B(_11615_),
    .Y(_11622_)
);

NAND3X1 _15673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5205_),
    .B(_5207_),
    .C(_5202_),
    .Y(_5215_)
);

AOI21X1 _15253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .B(_4750_),
    .C(_4748_),
    .Y(_4755_)
);

NOR2X1 _16878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6523_),
    .B(_6521_),
    .Y(_6535_)
);

NAND3X1 _16458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6066_),
    .B(_6069_),
    .C(_6072_),
    .Y(_6073_)
);

OAI21X1 _16038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5455_),
    .B(_5450_),
    .C(_5457_),
    .Y(_5615_)
);

FILL SFILL59320x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_9153_),
    .Y(_11812_)
);

AOI21X1 _21271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11339_),
    .B(_11338_),
    .C(_11335_),
    .Y(_11351_)
);

OAI21X1 _12798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_4434__bF$buf3),
    .C(_10452_),
    .Y(_188_)
);

NAND3X1 _12378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7316_),
    .B(_7404_),
    .C(_7481_),
    .Y(_7492_)
);

INVX1 _22896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .Y(_1223_)
);

NAND3X1 _22476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_759_),
    .C(_758_),
    .Y(_763_)
);

NAND2X1 _22056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_24_bF$buf2),
    .Y(_303_)
);

NAND3X1 _18604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8426_),
    .B(_8427_),
    .C(_8425_),
    .Y(_8428_)
);

FILL FILL74200x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33720x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9370_),
    .B(_9360_),
    .Y(_9749_)
);

NOR3X1 _14944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4411_),
    .B(_4407_),
    .C(_4410_),
    .Y(_4416_)
);

NAND2X1 _14524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf1),
    .B(areg_19_bF$buf0),
    .Y(_3957_)
);

OAI21X1 _14104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3494_),
    .B(_3496_),
    .C(_3492_),
    .Y(_3497_)
);

AOI21X1 _15729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5263_),
    .B(_5257_),
    .C(_5007_),
    .Y(_5276_)
);

OAI21X1 _15309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4498_),
    .B(_4815_),
    .C(_4507_),
    .Y(_4816_)
);

AOI21X1 _20962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10962_),
    .B(_10955_),
    .C(_10813_),
    .Y(_11013_)
);

AOI21X1 _20542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10535_),
    .B(_10539_),
    .C(_10542_),
    .Y(_10553_)
);

NAND2X1 _20122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10040_),
    .B(_10037_),
    .Y(_10092_)
);

NOR3X1 _19982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9570_),
    .B(_9569_),
    .C(_9572_),
    .Y(_9939_)
);

NOR3X1 _19562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9468_),
    .B(_9463_),
    .C(_9469_),
    .Y(_9479_)
);

AND2X2 _19142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_19_bF$buf5),
    .Y(_9018_)
);

FILL SFILL58840x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11869_),
    .B(_11871_),
    .Y(_11872_)
);

NAND3X1 _21327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11398_),
    .B(_11393_),
    .C(_11403_),
    .Y(_11413_)
);

NAND2X1 _15482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5000_),
    .B(_4998_),
    .Y(_5005_)
);

NOR2X1 _15062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4250_),
    .B(_4545_),
    .Y(_4546_)
);

AOI21X1 _16687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6324_),
    .B(_6325_),
    .C(_6309_),
    .Y(_6326_)
);

NAND3X1 _16267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5858_),
    .B(_5865_),
    .C(_5845_),
    .Y(_5866_)
);

FILL SFILL69000x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3253__bF$buf0),
    .B(_4551__bF$buf4),
    .C(_11141_),
    .Y(_11142_)
);

FILL SFILL69400x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5244_),
    .B(_5278_),
    .C(_5091_),
    .Y(_5398_)
);

OAI21X1 _22285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_553_),
    .C(_551_),
    .Y(_554_)
);

AOI21X1 _18833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8678_),
    .B(_8677_),
    .C(_8675_),
    .Y(_8679_)
);

NAND3X1 _18413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8210_),
    .B(_8196_),
    .C(_8214_),
    .Y(_8219_)
);

FILL SFILL74280x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_30_bF$buf3),
    .C(_9537_),
    .Y(_9540_)
);

FILL SFILL74600x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_14_bF$buf0),
    .Y(_4207_)
);

NAND3X1 _14333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3746_),
    .B(_3747_),
    .C(_3744_),
    .Y(_3748_)
);

DFFPOSX1 _24011_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[1]),
    .CLK(clk_bF$buf10),
    .D(a[1])
);

FILL SFILL74200x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .B(_5186_),
    .C(_5189_),
    .Y(_5527_)
);

NAND3X1 _15538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5043_),
    .B(_5059_),
    .C(_5065_),
    .Y(_5066_)
);

NOR3X1 _15118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4298_),
    .B(_4299_),
    .C(_4297_),
    .Y(_4607_)
);

AOI21X1 _20771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10462_),
    .B(_10548_),
    .C(_10552_),
    .Y(_10804_)
);

AOI21X1 _20351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10291_),
    .B(_10297_),
    .C(_9998_),
    .Y(_10343_)
);

AOI21X1 _19791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9320_),
    .B(_9353_),
    .C(_9357_),
    .Y(_9730_)
);

OAI21X1 _19371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8923_),
    .B(_8893_),
    .C(_8931_),
    .Y(_9269_)
);

OAI21X1 _21976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_196_),
    .C(_198_),
    .Y(_216_)
);

OAI22X1 _21556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11383_),
    .B(_11442_),
    .C(_11662_),
    .D(_11441_),
    .Y(_11663_)
);

OAI21X1 _21136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11202_),
    .B(_11203_),
    .C(_11199_),
    .Y(_11204_)
);

OAI21X1 _15291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4790_),
    .B(_4791_),
    .C(_4775_),
    .Y(_4797_)
);

AOI21X1 _13604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2943_),
    .B(_2944_),
    .C(_2942_),
    .Y(_2950_)
);

NAND2X1 _23702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2098_),
    .B(_2100_),
    .Y(_2101_)
);

NAND3X1 _16496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6111_),
    .B(_6115_),
    .C(_6114_),
    .Y(_6116_)
);

NAND2X1 _16076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5655_),
    .B(_5656_),
    .Y(_5657_)
);

AOI21X1 _14809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3981_),
    .B(_3979_),
    .C(_4267_),
    .Y(_4268_)
);

AOI21X1 _22094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_337_),
    .C(_336_),
    .Y(_345_)
);

AOI21X1 _18642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8464_),
    .B(_8465_),
    .C(_8468_),
    .Y(_8469_)
);

NAND3X1 _18222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7991_),
    .B(_7996_),
    .C(_7926_),
    .Y(_8010_)
);

FILL SFILL23720x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf2),
    .B(areg_27_bF$buf3),
    .Y(_10865_)
);

OAI21X1 _20407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf2),
    .B(_5315__bF$buf4),
    .C(_10396_),
    .Y(_10404_)
);

INVX2 _23299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .Y(_1661_)
);

OAI21X1 _19847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9460_),
    .B(_9427_),
    .C(_9452_),
    .Y(_9791_)
);

OR2X2 _19427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9324_),
    .B(_9325_),
    .Y(_9330_)
);

NOR3X1 _19007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8443_),
    .B(_8447_),
    .C(_8449_),
    .Y(_8870_)
);

AND2X2 _14982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_13_bF$buf2),
    .Y(_4457_)
);

NOR3X1 _14562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3699_),
    .B(_3695_),
    .C(_3703_),
    .Y(_3999_)
);

OAI21X1 _14142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3283_),
    .B(_3281_),
    .C(_3273_),
    .Y(_3538_)
);

FILL SFILL8680x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5311_),
    .B(_5316_),
    .C(_5314_),
    .Y(_5317_)
);

NAND2X1 _15347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4539_),
    .B(_4857_),
    .Y(_4858_)
);

NAND3X1 _20580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10592_),
    .B(_10591_),
    .C(_10593_),
    .Y(_10594_)
);

OAI21X1 _20160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10124_),
    .B(_10120_),
    .C(_10118_),
    .Y(_10133_)
);

FILL SFILL48840x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_22_bF$buf3),
    .Y(_9059_)
);

AOI21X1 _21785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_5_),
    .C(_11896_),
    .Y(_6_)
);

INVX2 _21365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11447_),
    .Y(_11455_)
);

INVX2 _17913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7669_),
    .Y(_7670_)
);

FILL SFILL74280x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3184_),
    .B(_3188_),
    .C(_3096_),
    .Y(_3201_)
);

OAI21X1 _13413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2737_),
    .C(_2552_),
    .Y(_2741_)
);

BUFX2 _23931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[49]),
    .Y(y[49])
);

XOR2X1 _23511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_1891_),
    .Y(_1892_)
);

FILL SFILL34120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43800x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74200x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4057_),
    .Y(_4058_)
);

FILL SFILL69560x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8719_),
    .B(_8718_),
    .C(_8703_),
    .Y(_8721_)
);

NAND3X1 _18451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8255_),
    .B(_8256_),
    .C(_8259_),
    .Y(_8261_)
);

FILL SFILL64280x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _18031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf2),
    .B(_3253__bF$buf1),
    .C(_2287__bF$buf3),
    .D(_3529__bF$buf4),
    .Y(_7800_)
);

AOI21X1 _20636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9993_),
    .B(_10316_),
    .C(_10655_),
    .Y(_10656_)
);

AOI21X1 _20216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10180_),
    .B(_10173_),
    .C(_10141_),
    .Y(_10195_)
);

FILL SFILL28840x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9570_),
    .B(_9569_),
    .C(_9572_),
    .Y(_9582_)
);

FILL SFILL64200x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9111_),
    .B(_9108_),
    .C(_9106_),
    .Y(_9121_)
);

INVX2 _14791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4247_),
    .Y(_4248_)
);

NAND2X1 _14371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg_20_bF$buf1),
    .Y(_3789_)
);

NOR3X1 _15996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5556_),
    .B(_5560_),
    .C(_5565_),
    .Y(_5569_)
);

XNOR2X1 _15576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5107_),
    .B(_5105_),
    .Y(_5108_)
);

NAND3X1 _15156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4643_),
    .B(_4646_),
    .C(_4647_),
    .Y(_4648_)
);

FILL SFILL54200x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11691_),
    .B(_11695_),
    .C(_11646_),
    .Y(_11705_)
);

XNOR2X1 _21174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11236_),
    .B(_11240_),
    .Y(_11246_)
);

AOI21X1 _17722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7458_),
    .B(_7460_),
    .C(_7444_),
    .Y(_7461_)
);

NAND3X1 _17302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6989_),
    .B(_6984_),
    .C(_6991_),
    .Y(_7001_)
);

FILL SFILL74120x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf0),
    .B(_6427_),
    .C(_1115_),
    .Y(_1116_)
);

NOR2X1 _22379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_653_),
    .Y(_657_)
);

NAND3X1 _18927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8779_),
    .B(_8374_),
    .C(_8781_),
    .Y(_8782_)
);

OAI21X1 _18507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8321_),
    .B(_7950_),
    .C(_7944_),
    .Y(_8322_)
);

OAI21X1 _13642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2765_),
    .C(_2767_),
    .Y(_2991_)
);

NAND2X1 _13222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .B(_2531_),
    .Y(_2532_)
);

OAI21X1 _23740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2139_),
    .C(_2140_),
    .Y(_2141_)
);

XOR2X1 _23320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1683_),
    .B(_1672_),
    .Y(_1684_)
);

FILL SFILL48920x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4004_),
    .B(_4011_),
    .C(_4013_),
    .Y(_4310_)
);

OAI21X1 _14427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3846_),
    .B(_3845_),
    .C(_3808_),
    .Y(_3850_)
);

NAND2X1 _14007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf3),
    .B(areg_16_bF$buf2),
    .Y(_3390_)
);

FILL SFILL13720x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8509_),
    .B(_8503_),
    .C(_8488_),
    .Y(_8510_)
);

OAI21X1 _18260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8049_),
    .B(_8050_),
    .C(_7661_),
    .Y(_8051_)
);

OAI21X1 _20865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10898_),
    .B(_10899_),
    .C(_10896_),
    .Y(_10907_)
);

NAND3X1 _20445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10429_),
    .B(_10434_),
    .C(_10436_),
    .Y(_10446_)
);

OAI21X1 _20025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9971_),
    .B(_9974_),
    .C(_9977_),
    .Y(_9985_)
);

AOI21X1 _19885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9831_),
    .B(_9832_),
    .C(_9786_),
    .Y(_9833_)
);

OAI21X1 _19465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9366_),
    .B(_9368_),
    .C(_9319_),
    .Y(_9372_)
);

AOI21X1 _19045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8905_),
    .B(_8910_),
    .C(_8898_),
    .Y(_8911_)
);

AOI21X1 _14180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3574_),
    .B(_3575_),
    .C(_3573_),
    .Y(_3579_)
);

FILL SFILL38920x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1434_),
    .B(_11701_),
    .C(_34_),
    .Y(_1445_)
);

FILL SFILL38840x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34120x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4769_),
    .B(_4810_),
    .C(_4809_),
    .Y(_4900_)
);

BUFX2 BUFX2_insert100 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf0)
);

BUFX2 BUFX2_insert101 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf5)
);

BUFX2 BUFX2_insert102 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf4)
);

BUFX2 BUFX2_insert103 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf3)
);

NAND2X1 _17951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_26_bF$buf2),
    .Y(_7712_)
);

BUFX2 BUFX2_insert104 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf2)
);

BUFX2 BUFX2_insert105 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf1)
);

OAI21X1 _17531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf1),
    .B(_5668__bF$buf0),
    .C(_7237_),
    .Y(_7251_)
);

BUFX2 BUFX2_insert106 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(breg_7_bF$buf0)
);

NAND3X1 _17111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6788_),
    .B(_6789_),
    .C(_6790_),
    .Y(_6792_)
);

BUFX2 BUFX2_insert107 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434_),
    .Y(_4434__bF$buf3)
);

BUFX2 BUFX2_insert108 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434_),
    .Y(_4434__bF$buf2)
);

BUFX2 BUFX2_insert109 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434_),
    .Y(_4434__bF$buf1)
);

FILL SFILL28840x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _22188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_203_),
    .Y(_448_)
);

NAND3X1 _18736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8527_),
    .B(_8567_),
    .C(_8571_),
    .Y(_8572_)
);

AOI21X1 _18316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7669_),
    .B(_7693_),
    .C(_7691_),
    .Y(_8112_)
);

AOI21X1 _13871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3238_),
    .B(_2980_),
    .C(_3240_),
    .Y(_3242_)
);

NAND2X1 _13451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2780_),
    .B(_2762_),
    .Y(_2782_)
);

NAND3X1 _13031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2325_),
    .B(_2324_),
    .C(_2323_),
    .Y(_2326_)
);

FILL SFILL13800x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf2),
    .B(_2763_),
    .Y(_4100_)
);

OAI21X1 _14236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3359_),
    .B(_3640_),
    .C(_3368_),
    .Y(_3641_)
);

FILL SFILL13400x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18840x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10460_),
    .B(_10696_),
    .C(_10626_),
    .Y(_10697_)
);

OAI21X1 _20254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10235_),
    .B(_10236_),
    .C(_10230_),
    .Y(_10237_)
);

OAI21X1 _16802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf1),
    .B(_5318_),
    .C(_6447_),
    .Y(_6452_)
);

NOR3X1 _19694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9233_),
    .B(_9237_),
    .C(_9240_),
    .Y(_9624_)
);

AND2X2 _19274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8369_),
    .B(_9156_),
    .Y(_9163_)
);

INVX2 _21879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .Y(_109_)
);

OAI21X1 _21459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11551_),
    .B(_11557_),
    .C(_11325_),
    .Y(_11558_)
);

NAND3X1 _21039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11059_),
    .B(_11096_),
    .C(_11091_),
    .Y(_11097_)
);

OAI21X1 _12722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11220_),
    .B(_11209_),
    .C(_11198_),
    .Y(_11264_)
);

XNOR2X1 _12302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6417_),
    .B(_6363_),
    .Y(_6659_)
);

NAND2X1 _22820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_25_bF$buf1),
    .B(breg_25_bF$buf1),
    .Y(_1139_)
);

AOI21X1 _22400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_678_),
    .C(_499_),
    .Y(_679_)
);

NOR2X1 _15194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4688_),
    .B(_4689_),
    .Y(_4690_)
);

FILL SFILL48920x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3299_),
    .B(_3300_),
    .C(_3302_),
    .Y(_3303_)
);

OAI21X1 _13507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2631_),
    .C(_2842_),
    .Y(_2843_)
);

OAI21X1 _23605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1940_),
    .B(_1939_),
    .C(_1937_),
    .Y(_1995_)
);

NAND3X1 _16399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6003_),
    .B(_5667_),
    .C(_6009_),
    .Y(_6010_)
);

AOI21X1 _17760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7494_),
    .B(_7491_),
    .C(_7489_),
    .Y(_7502_)
);

OAI21X1 _17340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7040_),
    .B(_7041_),
    .C(_7039_),
    .Y(_7042_)
);

FILL SFILL34200x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8805_),
    .B(_8823_),
    .C(_8804_),
    .Y(_8824_)
);

NAND2X1 _18545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_30_bF$buf3),
    .Y(_8364_)
);

NAND2X1 _18125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_23_bF$buf2),
    .Y(_7903_)
);

FILL SFILL59080x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3019_),
    .B(_3010_),
    .C(_3018_),
    .Y(_3032_)
);

AND2X2 _13260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2569_),
    .Y(_2572_)
);

FILL SFILL38920x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4301_),
    .B(_4308_),
    .C(_4065_),
    .Y(_4351_)
);

OAI21X1 _14465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3890_),
    .B(_3891_),
    .C(_3875_),
    .Y(_3892_)
);

NOR3X1 _14045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3428_),
    .B(_3426_),
    .C(_3425_),
    .Y(_3432_)
);

OAI21X1 _20483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10487_),
    .B(_10486_),
    .C(_10470_),
    .Y(_10488_)
);

OAI21X1 _20063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10026_),
    .B(_10019_),
    .C(_10005_),
    .Y(_10027_)
);

FILL SFILL28920x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6240_),
    .B(_6241_),
    .C(_6239_),
    .Y(_6243_)
);

AOI21X1 _19083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8946_),
    .B(_8945_),
    .C(_8944_),
    .Y(_8953_)
);

NOR3X1 _21688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11805_),
    .B(_11807_),
    .C(_11806_),
    .Y(_11808_)
);

OAI21X1 _21268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf1),
    .B(_6050__bF$buf3),
    .C(_11337_),
    .Y(_11347_)
);

NAND3X1 _17816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7551_),
    .B(_7546_),
    .C(_7554_),
    .Y(_7564_)
);

OAI21X1 _12951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1772_),
    .B(_1783_),
    .C(_1751_),
    .Y(_1860_)
);

OAI21X1 _12531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9159_),
    .B(_9148_),
    .C(_9049_),
    .Y(_9170_)
);

AOI21X1 _12111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4477_),
    .B(_4412_),
    .C(_4368_),
    .Y(_4566_)
);

FILL SFILL18920x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3091_),
    .B(_3092_),
    .C(_3093_),
    .Y(_3094_)
);

XNOR2X1 _13316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2633_),
    .B(_2630_),
    .Y(_2634_)
);

AOI22X1 _23834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2241_),
    .B(_2231_),
    .C(_2233_),
    .D(_2219_),
    .Y(_2242_)
);

NAND2X1 _23414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(_1786_),
    .Y(_1787_)
);

FILL SFILL18840x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _18774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_19_bF$buf5),
    .Y(_8614_)
);

AOI21X1 _18354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7809_),
    .B(_7791_),
    .C(_7813_),
    .Y(_8154_)
);

OAI21X1 _20959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11008_),
    .B(_10695_),
    .C(_10980_),
    .Y(_11009_)
);

NAND3X1 _20539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10462_),
    .B(_10543_),
    .C(_10548_),
    .Y(_10549_)
);

AOI21X1 _20119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10076_),
    .B(_10072_),
    .C(_10043_),
    .Y(_10088_)
);

AND2X2 _21900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11764_),
    .B(_131_),
    .Y(_132_)
);

OAI21X1 _19979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9917_),
    .B(_9922_),
    .C(_9927_),
    .Y(_9935_)
);

NAND3X1 _19559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9391_),
    .B(_9474_),
    .C(_9470_),
    .Y(_9475_)
);

OAI21X1 _19139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8611_),
    .B(_8626_),
    .C(_8617_),
    .Y(_9014_)
);

AOI21X1 _14694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4137_),
    .B(_4136_),
    .C(_4135_),
    .Y(_4142_)
);

NOR3X1 _14274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3678_),
    .B(_3682_),
    .C(_3681_),
    .Y(_3683_)
);

AOI21X1 _15899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5223_),
    .B(_5227_),
    .C(_5150_),
    .Y(_5462_)
);

NAND3X1 _15479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4764_),
    .B(_5000_),
    .C(_4916_),
    .Y(_5001_)
);

OAI21X1 _15059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_4541__bF$buf4),
    .C(_4250_),
    .Y(_4542_)
);

FILL SFILL3720x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10276_),
    .B(_10278_),
    .Y(_10279_)
);

NAND3X1 _16840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6488_),
    .B(_6489_),
    .C(_6440_),
    .Y(_6493_)
);

NAND2X1 _16420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6032_),
    .B(_6029_),
    .Y(_6033_)
);

NAND2X1 _16000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5553_),
    .B(_5549_),
    .Y(_5573_)
);

OAI21X1 _21497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11576_),
    .B(_11324_),
    .C(_11567_),
    .Y(_11599_)
);

AOI21X1 _21077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10829_),
    .B(_10832_),
    .C(_10839_),
    .Y(_11139_)
);

NAND2X1 _17625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_19_bF$buf5),
    .Y(_7354_)
);

NAND3X1 _17205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6847_),
    .B(_6888_),
    .C(_6893_),
    .Y(_6894_)
);

FILL SFILL59080x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10419_),
    .B(_11187_),
    .C(_11275_),
    .Y(_11679_)
);

NOR2X1 _12340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5826_),
    .B(_5837_),
    .Y(_7076_)
);

FILL SFILL3640x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3098_),
    .B(_3124_),
    .C(_3114_),
    .Y(_3344_)
);

OAI21X1 _13545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf0),
    .B(_2884__bF$buf0),
    .C(_2881_),
    .Y(_2885_)
);

OR2X2 _13125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2034_),
    .B(_2424_),
    .Y(_2425_)
);

NOR2X1 _23643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2033_),
    .B(_2030_),
    .Y(_2037_)
);

NAND2X1 _23223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .B(areg_28_bF$buf4),
    .Y(_1578_)
);

DFFPOSX1 _24008_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[62]),
    .CLK(clk_bF$buf3),
    .D(_0_[62])
);

FILL SFILL49080x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8332_),
    .B(_8398_),
    .C(_8395_),
    .Y(_8405_)
);

AOI21X1 _18163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7939_),
    .B(_7940_),
    .C(_7932_),
    .Y(_7945_)
);

FILL SFILL49000x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10798_),
    .B(_10799_),
    .C(_10794_),
    .Y(_10800_)
);

OAI21X1 _20348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10338_),
    .B(_10318_),
    .C(_10311_),
    .Y(_10339_)
);

AOI21X1 _19788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9711_),
    .B(_9715_),
    .C(_9716_),
    .Y(_9726_)
);

OAI21X1 _19368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7651_),
    .B(_9264_),
    .C(_9263_),
    .Y(_9265_)
);

OAI21X1 _14083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3473_),
    .B(_3472_),
    .C(_3468_),
    .Y(_3474_)
);

FILL SFILL18920x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_374_),
    .Y(_385_)
);

AOI21X1 _22914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1242_),
    .C(_1099_),
    .Y(_1243_)
);

NAND3X1 _15288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4788_),
    .B(_4792_),
    .C(_4773_),
    .Y(_4793_)
);

NAND3X1 _17854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7224_),
    .B(_7339_),
    .C(_7337_),
    .Y(_7606_)
);

OAI21X1 _17434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7138_),
    .B(_7139_),
    .C(_7093_),
    .Y(_7146_)
);

OR2X2 _17014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6683_),
    .B(_6684_),
    .Y(_6685_)
);

FILL SFILL74440x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8460_),
    .B(_8461_),
    .C(_8070_),
    .Y(_8465_)
);

NOR3X1 _18219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7570_),
    .B(_7571_),
    .C(_7568_),
    .Y(_8006_)
);

INVX1 _13774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3129_),
    .Y(_3135_)
);

NOR3X1 _13354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2663_),
    .B(_2667_),
    .C(_2673_),
    .Y(_2676_)
);

AOI21X1 _23872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2279_),
    .B(_2278_),
    .C(_2281_),
    .Y(_2282_)
);

NAND3X1 _23452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1824_),
    .B(_1828_),
    .C(_1781_),
    .Y(_1829_)
);

NOR3X1 _23032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .B(_1219_),
    .C(_1222_),
    .Y(_1371_)
);

FILL SFILL53880x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4173_),
    .B(_4164_),
    .C(_4168_),
    .Y(_4454_)
);

OAI21X1 _14559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3978_),
    .B(_3982_),
    .C(_3985_),
    .Y(_3995_)
);

NAND2X1 _14139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3524_),
    .B(_3532_),
    .Y(_3534_)
);

FILL SFILL3720x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43960x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .B(_5484_),
    .C(_5472_),
    .Y(_5485_)
);

NOR3X1 _15500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5020_),
    .B(_5022_),
    .C(_5023_),
    .Y(_5024_)
);

OAI21X1 _18392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7804_),
    .B(_7794_),
    .C(_7798_),
    .Y(_8196_)
);

NOR3X1 _20997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11048_),
    .B(_11049_),
    .C(_11050_),
    .Y(_11051_)
);

AND2X2 _20577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10238_),
    .B(_10229_),
    .Y(_10591_)
);

OAI21X1 _20157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10125_),
    .B(_10129_),
    .C(_10117_),
    .Y(_10130_)
);

OAI21X1 _16705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6338_),
    .B(_6339_),
    .C(_6293_),
    .Y(_6346_)
);

NAND3X1 _19597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9516_),
    .B(_9509_),
    .C(_9515_),
    .Y(_9517_)
);

NAND3X1 _19177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9055_),
    .B(_9048_),
    .C(_9052_),
    .Y(_9056_)
);

FILL SFILL43880x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43800x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_10_bF$buf5),
    .Y(_10200_)
);

NAND3X1 _12205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4105_),
    .B(_5508_),
    .C(_5585_),
    .Y(_5596_)
);

NOR2X1 _22723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_1033_),
    .Y(_1034_)
);

NAND3X1 _22303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_572_),
    .C(_573_),
    .Y(_574_)
);

NAND3X1 _15097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4578_),
    .B(_4583_),
    .C(_4495_),
    .Y(_4584_)
);

BUFX2 _23928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[46]),
    .Y(y[46])
);

XOR2X1 _23508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1888_),
    .B(_1885_),
    .Y(_1889_)
);

FILL SFILL49080x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7389_),
    .B(_7390_),
    .C(_7381_),
    .Y(_7396_)
);

NOR2X1 _17243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6533_),
    .B(_6935_),
    .Y(_6936_)
);

FILL SFILL33880x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_25_bF$buf4),
    .Y(_8717_)
);

NOR3X1 _18448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8242_),
    .B(_8239_),
    .C(_8241_),
    .Y(_8257_)
);

AND2X2 _18028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_19_bF$buf5),
    .Y(_7796_)
);

OAI21X1 _13583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2829_),
    .B(_2830_),
    .C(_2827_),
    .Y(_2927_)
);

NAND3X1 _13163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2460_),
    .B(_2466_),
    .C(_2463_),
    .Y(_2467_)
);

NAND3X1 _23681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_28_bF$buf3),
    .B(breg_29_bF$buf2),
    .C(_2076_),
    .Y(_2078_)
);

XOR2X1 _23261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1619_),
    .B(_1617_),
    .Y(_1621_)
);

FILL SFILL39080x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf2),
    .B(areg_22_bF$buf1),
    .Y(_4245_)
);

NOR2X1 _14368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3254_),
    .B(_3528_),
    .Y(_3784_)
);

FILL SFILL23800x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24046_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[4]),
    .CLK(clk_bF$buf10),
    .D(b[4])
);

FILL SFILL8840x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53960x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[24]),
    .Y(areg_24_bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[24]),
    .Y(areg_24_bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[24]),
    .Y(areg_24_bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[24]),
    .Y(areg_24_bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[24]),
    .Y(areg_24_bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258_),
    .Y(_4258__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258_),
    .Y(_4258__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258_),
    .Y(_4258__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258_),
    .Y(_4258__bF$buf0)
);

AOI21X1 _20386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10380_),
    .B(_10377_),
    .C(_10352_),
    .Y(_10381_)
);

OAI21X1 _16934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6590_),
    .B(_6591_),
    .C(_6592_),
    .Y(_6597_)
);

XNOR2X1 _16514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6135_),
    .B(_6133_),
    .Y(_6136_)
);

FILL SFILL53960x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74120x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48920x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7026_),
    .B(_7030_),
    .C(_7035_),
    .Y(_7457_)
);

OAI21X1 _12854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_724_),
    .C(_385_),
    .Y(_801_)
);

NAND3X1 _12434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7931_),
    .B(_7997_),
    .C(_8029_),
    .Y(_8106_)
);

XOR2X1 _22952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1283_),
    .B(_1273_),
    .Y(_1284_)
);

NAND2X1 _12014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg_5_bF$buf0),
    .Y(_3503_)
);

OAI21X1 _22532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_820_),
    .C(_772_),
    .Y(_825_)
);

NAND3X1 _22112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_361_),
    .B(_362_),
    .C(_363_),
    .Y(_364_)
);

OAI21X1 _13639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2986_),
    .B(_2942_),
    .C(_2934_),
    .Y(_2987_)
);

NAND3X1 _13219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .B(_2517_),
    .C(_2522_),
    .Y(_2528_)
);

NAND2X1 _23737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_27_bF$buf3),
    .B(areg_30_bF$buf0),
    .Y(_2138_)
);

OAI21X1 _23317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(_1679_),
    .C(_1680_),
    .Y(_1681_)
);

FILL SFILL74360x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7642_),
    .B(_7209_),
    .C(_7633_),
    .Y(_7647_)
);

NAND2X1 _17472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7184_),
    .B(_7186_),
    .Y(_7187_)
);

OAI21X1 _17052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6724_),
    .B(_6726_),
    .C(_6723_),
    .Y(_6727_)
);

FILL SFILL23960x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8505_),
    .B(_8506_),
    .C(_8491_),
    .Y(_8507_)
);

NAND3X1 _18257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7660_),
    .B(_8042_),
    .C(_8043_),
    .Y(_8048_)
);

NAND3X1 _13392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2711_),
    .B(_2577_),
    .C(_2717_),
    .Y(_2718_)
);

FILL FILL74120x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1787_),
    .B(_1868_),
    .Y(_1869_)
);

NOR2X1 _23070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1274_),
    .B(_1281_),
    .Y(_1411_)
);

OAI21X1 _21803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11686_),
    .B(_25_),
    .C(_11678_),
    .Y(_26_)
);

AOI21X1 _14597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3520_),
    .B(_3751_),
    .C(_3758_),
    .Y(_4037_)
);

NAND3X1 _14177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3574_),
    .B(_3575_),
    .C(_3573_),
    .Y(_3576_)
);

OAI21X1 _20195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10170_),
    .B(_10171_),
    .C(_10169_),
    .Y(_10172_)
);

NAND2X1 _16743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6386_),
    .B(_6387_),
    .Y(_6388_)
);

AND2X2 _16323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5923_),
    .B(_5927_),
    .Y(_5928_)
);

OAI21X1 _17948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7707_),
    .B(_7310_),
    .C(_7302_),
    .Y(_7708_)
);

AOI21X1 _17528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7242_),
    .B(_7246_),
    .C(_7234_),
    .Y(_7247_)
);

INVX1 _17108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6421_),
    .Y(_6788_)
);

FILL SFILL18600x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8961_),
    .B(_10606_),
    .C(_8994_),
    .Y(_10617_)
);

AOI21X1 _12243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6001_),
    .B(_5990_),
    .C(_5870_),
    .Y(_6012_)
);

INVX2 _22761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .Y(_1076_)
);

XNOR2X1 _22341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_614_),
    .B(_609_),
    .Y(_616_)
);

FILL SFILL59080x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8920x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _13868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2980_),
    .B(_3238_),
    .Y(_0_[18])
);

FILL SFILL23800x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2775_),
    .B(_2777_),
    .Y(_2778_)
);

DFFPOSX1 _23966_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[20]),
    .CLK(clk_bF$buf2),
    .D(_0_[20])
);

AND2X2 _13028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1870_),
    .Y(_2323_)
);

OAI21X1 _23546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1841_),
    .B(_1727_),
    .C(_1847_),
    .Y(_1931_)
);

NAND2X1 _23126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1461_),
    .Y(_1473_)
);

NAND3X1 _17281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6969_),
    .B(_6973_),
    .C(_6976_),
    .Y(_6978_)
);

FILL SFILL13880x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _18486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_5921__bF$buf2),
    .C(_7217__bF$buf4),
    .D(_4541__bF$buf1),
    .Y(_8299_)
);

NAND2X1 _18066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_19_bF$buf5),
    .Y(_7838_)
);

FILL SFILL74120x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2617_),
    .Y(_2628_)
);

NOR2X1 _21612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11722_),
    .B(_11724_),
    .Y(_11725_)
);

FILL SFILL29000x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11198_),
    .B(_11209_),
    .C(_11220_),
    .Y(_11231_)
);

NAND2X1 _22817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1134_),
    .B(_1135_),
    .Y(_1136_)
);

AOI21X1 _16972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6633_),
    .B(_6634_),
    .C(_6632_),
    .Y(_6639_)
);

AND2X2 _16552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .B(_6177_),
    .Y(_6178_)
);

NAND3X1 _16132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5712_),
    .B(_5671_),
    .C(_5717_),
    .Y(_5718_)
);

OAI21X1 _17757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7104_),
    .B(_7094_),
    .C(_7099_),
    .Y(_7499_)
);

AOI21X1 _17337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6612_),
    .B(_6616_),
    .C(_6619_),
    .Y(_7039_)
);

AOI21X1 _12892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9948_),
    .B(_11527_),
    .C(_11549_),
    .Y(_1217_)
);

INVX2 _12472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8511_),
    .Y(_8522_)
);

NAND3X1 _22990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1319_),
    .B(_1323_),
    .C(_1295_),
    .Y(_1324_)
);

AOI21X1 _12052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2431_),
    .B(_2989_),
    .C(_3011_),
    .Y(_3920_)
);

NAND2X1 _22570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf2),
    .B(areg_31_bF$buf2),
    .Y(_866_)
);

NOR2X1 _22150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(_405_),
    .Y(_406_)
);

OAI21X1 _13677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3028_),
    .B(_3020_),
    .C(_2990_),
    .Y(_3029_)
);

OAI21X1 _13257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2567_),
    .B(_2568_),
    .C(_2368_),
    .Y(_2569_)
);

NAND2X1 _23775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_29_bF$buf2),
    .B(areg_30_bF$buf0),
    .Y(_2179_)
);

AND2X2 _23355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1719_),
    .B(_1716_),
    .Y(_1723_)
);

OAI21X1 _19903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9852_),
    .B(_9851_),
    .C(_9849_),
    .Y(_9853_)
);

AOI21X1 _17090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6750_),
    .B(_6755_),
    .C(_6600_),
    .Y(_6768_)
);

OAI21X1 _15823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5020_),
    .B(_5023_),
    .C(_5027_),
    .Y(_5379_)
);

NOR3X1 _15403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4912_),
    .B(_4913_),
    .C(_4909_),
    .Y(_4920_)
);

AND2X2 _18295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_28_bF$buf0),
    .Y(_8089_)
);

AOI21X1 _16608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5849_),
    .B(_5852_),
    .C(_5855_),
    .Y(_6239_)
);

NAND3X1 _21841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_66_),
    .B(_65_),
    .C(_64_),
    .Y(_68_)
);

AOI21X1 _21421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11514_),
    .B(_11515_),
    .C(_11513_),
    .Y(_11517_)
);

NAND3X1 _21001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11016_),
    .B(_11054_),
    .C(_11053_),
    .Y(_11056_)
);

FILL SFILL44040x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1489_),
    .B(_1816_),
    .C(_1762_),
    .Y(_1827_)
);

NAND2X1 _12528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_11_bF$buf1),
    .Y(_9137_)
);

INVX1 _22626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9985_),
    .Y(_927_)
);

NAND3X1 _12108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4325_),
    .B(_4478_),
    .C(_4522_),
    .Y(_4533_)
);

AOI21X1 _22206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11885_),
    .B(_216_),
    .C(_467_),
    .Y(_468_)
);

NOR2X1 _16781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf2),
    .B(_6427_),
    .Y(_6429_)
);

NOR3X1 _16361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5582_),
    .C(_5580_),
    .Y(_5970_)
);

BUFX2 BUFX2_insert450 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420_),
    .Y(_5420__bF$buf3)
);

BUFX2 BUFX2_insert451 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420_),
    .Y(_5420__bF$buf2)
);

BUFX2 BUFX2_insert452 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420_),
    .Y(_5420__bF$buf1)
);

BUFX2 BUFX2_insert453 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420_),
    .Y(_5420__bF$buf0)
);

BUFX2 BUFX2_insert454 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf4)
);

NAND3X1 _17986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7708_),
    .B(_7745_),
    .C(_7749_),
    .Y(_7750_)
);

AOI21X1 _17566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7282_),
    .B(_7284_),
    .C(_7281_),
    .Y(_7289_)
);

BUFX2 BUFX2_insert455 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf3)
);

NAND2X1 _17146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6824_),
    .B(_6825_),
    .Y(_6829_)
);

BUFX2 BUFX2_insert456 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf2)
);

BUFX2 BUFX2_insert457 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf1)
);

BUFX2 BUFX2_insert458 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[13]),
    .Y(areg_13_bF$buf0)
);

BUFX2 BUFX2_insert459 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[23]),
    .Y(breg_23_bF$buf3)
);

XNOR2X1 _12281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6417_),
    .B(_6374_),
    .Y(_6428_)
);

NAND3X1 _13486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2800_),
    .B(_2819_),
    .C(_2811_),
    .Y(_2820_)
);

INVX2 _13066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .Y(_2360_)
);

AOI21X1 _23584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1956_),
    .B(_1971_),
    .C(_924_),
    .Y(_1972_)
);

AOI21X1 _23164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1509_),
    .B(_1514_),
    .C(_1407_),
    .Y(_1515_)
);

AOI21X1 _19712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9588_),
    .B(_9589_),
    .C(_9390_),
    .Y(_9643_)
);

FILL SFILL64120x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4850_),
    .Y(_5170_)
);

OAI21X1 _15212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4415_),
    .B(_4417_),
    .C(_4409_),
    .Y(_4710_)
);

NAND3X1 _20289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10271_),
    .B(_10274_),
    .C(_10205_),
    .Y(_10275_)
);

NAND3X1 _16837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6488_),
    .B(_6489_),
    .C(_6487_),
    .Y(_6490_)
);

NOR3X1 _16417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6026_),
    .B(_6027_),
    .C(_6022_),
    .Y(_6030_)
);

NAND2X1 _11972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3033_),
    .B(_3000_),
    .Y(_3044_)
);

OAI21X1 _21650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2763_),
    .B(_6686__bF$buf2),
    .C(_11765_),
    .Y(_11766_)
);

NAND2X1 _21230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11306_),
    .B(_11301_),
    .Y(_11307_)
);

XNOR2X1 _12757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9937_),
    .B(_11636_),
    .Y(_0_[12])
);

NAND3X1 _12337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7032_),
    .B(_7031_),
    .C(_5804_),
    .Y(_7043_)
);

NAND3X1 _22855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1176_),
    .C(_1177_),
    .Y(_1178_)
);

OAI21X1 _22435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_237_),
    .B(_717_),
    .C(_716_),
    .Y(_718_)
);

NAND2X1 _22015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf5),
    .B(breg_29_bF$buf4),
    .Y(_258_)
);

OAI21X1 _16590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5978_),
    .B(_6218_),
    .C(_5968_),
    .Y(_6219_)
);

AOI21X1 _16170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5756_),
    .B(_5758_),
    .C(_5754_),
    .Y(_5759_)
);

NAND2X1 _14903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_18_bF$buf5),
    .Y(_4371_)
);

NAND3X1 _17795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7528_),
    .B(_7540_),
    .C(_7535_),
    .Y(_7541_)
);

AOI21X1 _17375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7072_),
    .B(_7071_),
    .C(_7068_),
    .Y(_7081_)
);

NAND2X1 _12090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_6_bF$buf4),
    .Y(_4336_)
);

NAND3X1 _20921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10962_),
    .B(_10955_),
    .C(_10813_),
    .Y(_10969_)
);

OAI21X1 _20501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf2),
    .B(_4541__bF$buf0),
    .C(_10503_),
    .Y(_10508_)
);

FILL SFILL44040x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(_2430_),
    .Y(_2610_)
);

OAI21X1 _23393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1760_),
    .B(_1759_),
    .C(_1660_),
    .Y(_1765_)
);

AOI21X1 _19941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9550_),
    .B(_9552_),
    .C(_9558_),
    .Y(_9894_)
);

OAI21X1 _19521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf4),
    .B(_3961__bF$buf0),
    .C(_9432_),
    .Y(_9434_)
);

OAI21X1 _19101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8969_),
    .B(_8968_),
    .C(_8971_),
    .Y(_8973_)
);

AOI21X1 _21706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11824_),
    .B(_11823_),
    .C(_11825_),
    .Y(_11828_)
);

AND2X2 _15861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5055_),
    .B(_5106_),
    .Y(_5421_)
);

NAND2X1 _15441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4960_),
    .B(_4957_),
    .Y(_4961_)
);

INVX2 _15021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4499_),
    .Y(_4501_)
);

NAND3X1 _20098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10044_),
    .B(_10059_),
    .C(_10064_),
    .Y(_10065_)
);

AOI21X1 _16646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6273_),
    .B(_6278_),
    .C(_6280_),
    .Y(_6281_)
);

NAND3X1 _16226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5811_),
    .B(_5805_),
    .C(_5809_),
    .Y(_5821_)
);

AOI21X1 _12986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(_560_),
    .C(_2228_),
    .Y(_2238_)
);

AOI21X1 _12566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7283_),
    .B(_8073_),
    .C(_9543_),
    .Y(_9554_)
);

NOR2X1 _12146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4939_),
    .B(_4019_),
    .Y(_4950_)
);

XNOR2X1 _22664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_958_),
    .B(_968_),
    .Y(_969_)
);

NAND2X1 _22244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf5),
    .B(breg_29_bF$buf4),
    .Y(_509_)
);

OAI21X1 _23869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2236_),
    .B(_2211_),
    .C(_2257_),
    .Y(_2278_)
);

FILL SFILL64120x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _23449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1801_),
    .B(_1782_),
    .Y(_1825_)
);

INVX2 _23029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .Y(_1367_)
);

XNOR2X1 _14712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4161_),
    .B(_4157_),
    .Y(_4162_)
);

OAI21X1 _17184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf3),
    .B(_3781__bF$buf2),
    .C(_6455_),
    .Y(_6871_)
);

FILL SFILL59160x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5478_),
    .B(_5481_),
    .Y(_5482_)
);

NAND3X1 _20730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10750_),
    .B(_10754_),
    .C(_10757_),
    .Y(_10758_)
);

NAND3X1 _20310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10291_),
    .B(_10297_),
    .C(_9998_),
    .Y(_10298_)
);

NAND2X1 _18389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_21_bF$buf4),
    .Y(_8192_)
);

FILL SFILL49160x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9648_),
    .B(_9676_),
    .C(_9672_),
    .Y(_9684_)
);

OAI21X1 _19330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9205_),
    .B(_9211_),
    .C(_9215_),
    .Y(_9224_)
);

FILL SFILL54120x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_170_),
    .C(_94_),
    .Y(_171_)
);

NAND3X1 _21515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11612_),
    .B(_11618_),
    .C(_11616_),
    .Y(_11619_)
);

NAND3X1 _15670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5206_),
    .B(_5210_),
    .C(_5193_),
    .Y(_5211_)
);

NAND3X1 _15250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4749_),
    .B(_4750_),
    .C(_4748_),
    .Y(_4751_)
);

NAND3X1 _16875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6519_),
    .B(_6528_),
    .C(_6526_),
    .Y(_6532_)
);

NAND2X1 _16455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_22_bF$buf1),
    .Y(_6070_)
);

OAI21X1 _16035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5610_),
    .B(_5611_),
    .C(_5609_),
    .Y(_5612_)
);

OAI21X1 _12795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10518_),
    .B(_10463_),
    .C(_10540_),
    .Y(_155_)
);

NAND2X1 _12375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7448_),
    .B(_7415_),
    .Y(_7459_)
);

NAND3X1 _22893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1219_),
    .B(_1183_),
    .C(_1188_),
    .Y(_1220_)
);

NAND3X1 _22473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_759_),
    .C(_758_),
    .Y(_760_)
);

NAND2X1 _22053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_25_bF$buf1),
    .Y(_300_)
);

AOI21X1 _18601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8015_),
    .B(_8017_),
    .C(_8423_),
    .Y(_8425_)
);

AOI22X1 _23678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_27_bF$buf3),
    .B(areg_30_bF$buf5),
    .C(breg_28_bF$buf5),
    .D(areg_29_bF$buf4),
    .Y(_2074_)
);

NOR2X1 _23258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5369_),
    .B(_9153_),
    .Y(_1617_)
);

AOI21X1 _19806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9391_),
    .B(_9470_),
    .C(_9479_),
    .Y(_9746_)
);

FILL SFILL69240x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4410_),
    .B(_4411_),
    .C(_4407_),
    .Y(_4413_)
);

AOI21X1 _14521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3930_),
    .B(_3951_),
    .C(_3952_),
    .Y(_3954_)
);

AOI21X1 _14101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3488_),
    .B(_3489_),
    .C(_3230_),
    .Y(_3494_)
);

FILL SFILL34040x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5261_),
    .B(_5262_),
    .C(_5008_),
    .Y(_5273_)
);

AOI21X1 _15306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4558_),
    .B(_4562_),
    .C(_4528_),
    .Y(_4813_)
);

OAI21X1 _18198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7971_),
    .B(_7972_),
    .C(_7965_),
    .Y(_7983_)
);

OAI21X1 _21744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11854_),
    .B(_11858_),
    .C(_11861_),
    .Y(_11869_)
);

OAI21X1 _21324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11408_),
    .B(_11409_),
    .C(_11407_),
    .Y(_11410_)
);

FILL SFILL3800x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _22949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(_1279_),
    .Y(_1280_)
);

OAI21X1 _22529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_819_),
    .B(_820_),
    .C(_818_),
    .Y(_821_)
);

AND2X2 _22109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_69_),
    .Y(_361_)
);

AOI21X1 _16684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5931_),
    .B(_5935_),
    .C(_5939_),
    .Y(_6323_)
);

AOI21X1 _16264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5861_),
    .B(_5862_),
    .C(_5847_),
    .Y(_5863_)
);

NOR2X1 _17889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7641_),
    .B(_7642_),
    .Y(_7643_)
);

NAND3X1 _17469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7177_),
    .B(_6919_),
    .C(_7182_),
    .Y(_7183_)
);

AOI21X1 _17049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6306_),
    .B(_6328_),
    .C(_6722_),
    .Y(_6723_)
);

OAI21X1 _12184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5267_),
    .B(_5256_),
    .C(_5124_),
    .Y(_5365_)
);

OAI21X1 _22282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf3),
    .B(_5315__bF$buf2),
    .C(_300_),
    .Y(_551_)
);

NOR2X1 _18830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8634_),
    .B(_8629_),
    .Y(_8675_)
);

NAND3X1 _18410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8209_),
    .B(_8210_),
    .C(_8214_),
    .Y(_8215_)
);

FILL SFILL33960x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2709_),
    .B(_2708_),
    .C(_2707_),
    .Y(_2714_)
);

AOI21X1 _23487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1864_),
    .B(_1774_),
    .C(_1865_),
    .Y(_1866_)
);

NAND2X1 _23067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(_1330_),
    .Y(_1408_)
);

NAND2X1 _19615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_29_bF$buf3),
    .Y(_9537_)
);

FILL SFILL18760x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3921_),
    .Y(_4203_)
);

AOI21X1 _14330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3457_),
    .B(_3309_),
    .C(_3463_),
    .Y(_3744_)
);

FILL SFILL18680x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33720x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf3),
    .B(_3402__bF$buf2),
    .C(_5518_),
    .Y(_5524_)
);

OAI21X1 _15535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf2),
    .B(_2586__bF$buf3),
    .C(_4723_),
    .Y(_5063_)
);

NAND3X1 _15115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4584_),
    .B(_4591_),
    .C(_4594_),
    .Y(_4604_)
);

NAND3X1 _21973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_212_),
    .C(_198_),
    .Y(_213_)
);

NAND3X1 _21553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11656_),
    .B(_11659_),
    .C(_11658_),
    .Y(_11660_)
);

OAI21X1 _21133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11185_),
    .B(_11186_),
    .C(_11183_),
    .Y(_11201_)
);

NAND3X1 _22758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1063_),
    .B(_1027_),
    .C(_1032_),
    .Y(_1072_)
);

OR2X2 _22338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_610_),
    .B(_611_),
    .Y(_612_)
);

NAND3X1 _13601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2941_),
    .B(_2945_),
    .C(_2760_),
    .Y(_2947_)
);

NAND3X1 _16493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6096_),
    .B(_6101_),
    .C(_6104_),
    .Y(_6113_)
);

NAND3X1 _16073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5653_),
    .B(_5646_),
    .C(_5284_),
    .Y(_5654_)
);

NAND3X1 _14806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4262_),
    .B(_4264_),
    .C(_4263_),
    .Y(_4265_)
);

FILL SFILL29000x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7433_),
    .B(_7429_),
    .Y(_7434_)
);

NAND2X1 _17278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_17_bF$buf4),
    .Y(_6974_)
);

FILL SFILL69160x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59320x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_53_),
    .Y(_342_)
);

FILL SFILL8600x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8520x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10851_),
    .B(_10861_),
    .Y(_10862_)
);

OAI21X1 _20404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10400_),
    .B(_10399_),
    .C(_10395_),
    .Y(_10401_)
);

NAND3X1 _13198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2503_),
    .B(_2504_),
    .C(_2502_),
    .Y(_2505_)
);

AOI21X1 _23296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1558_),
    .C(_1570_),
    .Y(_1658_)
);

AOI21X1 _19844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9772_),
    .B(_9777_),
    .C(_9765_),
    .Y(_9788_)
);

FILL SFILL3800x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9324_),
    .B(_9325_),
    .Y(_9327_)
);

OAI21X1 _19004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8854_),
    .B(_8857_),
    .C(_8860_),
    .Y(_8867_)
);

NAND2X1 _21609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf2),
    .B(areg_22_bF$buf2),
    .Y(_11721_)
);

FILL FILL74200x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5312_),
    .B(_5313_),
    .Y(_5314_)
);

NAND2X1 _15344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf0),
    .B(areg_22_bF$buf1),
    .Y(_4855_)
);

FILL SFILL49240x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6633_),
    .B(_6634_),
    .C(_6632_),
    .Y(_6635_)
);

OAI21X1 _16549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf0),
    .B(_2362__bF$buf3),
    .C(_6168_),
    .Y(_6174_)
);

NAND3X1 _16129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5700_),
    .B(_5704_),
    .C(_5710_),
    .Y(_5714_)
);

AOI21X1 _21782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11612_),
    .B(_11618_),
    .C(_11621_),
    .Y(_3_)
);

AND2X2 _21362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf4),
    .B(areg_24_bF$buf4),
    .Y(_11452_)
);

INVX1 _17910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7665_),
    .Y(_7666_)
);

FILL SFILL39160x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_1086_),
    .C(_11657_),
    .Y(_1184_)
);

AOI21X1 _12469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8084_),
    .B(_8117_),
    .C(_7196_),
    .Y(_8489_)
);

NOR2X1 _22987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1317_),
    .Y(_1321_)
);

OAI21X1 _12049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3865_),
    .B(_3876_),
    .C(_3471_),
    .Y(_3887_)
);

XNOR2X1 _22567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(_848_),
    .Y(_863_)
);

NOR2X1 _22147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11528_),
    .B(_178_),
    .Y(_403_)
);

AOI21X1 _13830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2923_),
    .B(_2840_),
    .C(_3196_),
    .Y(_3197_)
);

AOI21X1 _13410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2722_),
    .B(_2728_),
    .C(_2554_),
    .Y(_2737_)
);

OAI21X1 _14615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3516_),
    .B(_4054_),
    .C(_4053_),
    .Y(_4055_)
);

NOR3X1 _17087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6367_),
    .B(_6368_),
    .C(_6366_),
    .Y(_6765_)
);

FILL SFILL23960x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10652_),
    .B(_10651_),
    .C(_10340_),
    .Y(_10653_)
);

OAI21X1 _20213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10191_),
    .B(_9856_),
    .C(_9891_),
    .Y(_10192_)
);

NAND3X1 _19653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9474_),
    .B(_9470_),
    .C(_9476_),
    .Y(_9579_)
);

OAI21X1 _19233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9112_),
    .B(_9117_),
    .C(_9105_),
    .Y(_9118_)
);

FILL SFILL69320x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _21838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .Y(_64_)
);

NOR3X1 _21418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11225_),
    .B(_11247_),
    .C(_11245_),
    .Y(_11513_)
);

OAI21X1 _15993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5565_),
    .B(_5560_),
    .C(_5556_),
    .Y(_5566_)
);

NAND2X1 _15573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_14_bF$buf2),
    .Y(_5105_)
);

OAI21X1 _15153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4640_),
    .B(_4335_),
    .C(_4636_),
    .Y(_4645_)
);

FILL SFILL13960x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6049_),
    .Y(_6425_)
);

NAND3X1 _16358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5949_),
    .B(_5953_),
    .C(_5956_),
    .Y(_5966_)
);

OAI21X1 _21591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11517_),
    .B(_11440_),
    .C(_11520_),
    .Y(_11702_)
);

AND2X2 _21171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11236_),
    .B(_11240_),
    .Y(_11243_)
);

NAND3X1 _12698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10946_),
    .B(_10990_),
    .C(_10792_),
    .Y(_11000_)
);

NOR2X1 _12278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6187_),
    .B(_6385_),
    .Y(_6396_)
);

NAND2X1 _22796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf2),
    .B(breg_28_bF$buf3),
    .Y(_1113_)
);

NAND2X1 _22376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_653_),
    .Y(_654_)
);

INVX2 _18924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7968_),
    .Y(_8779_)
);

NAND3X1 _18504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8312_),
    .B(_8313_),
    .C(_8311_),
    .Y(_8319_)
);

FILL FILL74200x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9615_),
    .B(_9274_),
    .C(_9606_),
    .Y(_9639_)
);

NAND3X1 _14844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4287_),
    .B(_4294_),
    .C(_4297_),
    .Y(_4307_)
);

OAI21X1 _14424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3846_),
    .B(_3845_),
    .C(_3841_),
    .Y(_3847_)
);

NOR2X1 _14004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf3),
    .B(_2287__bF$buf2),
    .Y(_3387_)
);

NAND3X1 _15629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5165_),
    .B(_5160_),
    .C(_5163_),
    .Y(_5166_)
);

NAND3X1 _15209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4684_),
    .B(_4693_),
    .C(_4696_),
    .Y(_4706_)
);

NAND3X1 _20862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10815_),
    .B(_10897_),
    .C(_10903_),
    .Y(_10904_)
);

NAND3X1 _20442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10435_),
    .B(_10442_),
    .C(_10391_),
    .Y(_10443_)
);

XOR2X1 _20022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9634_),
    .B(_9982_),
    .Y(_0_[37])
);

AOI21X1 _19882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9822_),
    .B(_9829_),
    .C(_9790_),
    .Y(_9830_)
);

OAI21X1 _19462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9366_),
    .B(_9368_),
    .C(_9363_),
    .Y(_9369_)
);

NOR2X1 _19042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8498_),
    .B(_8907_),
    .Y(_8908_)
);

NOR2X1 _11969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2705_),
    .B(_2968_),
    .Y(_3011_)
);

NAND3X1 _21647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11757_),
    .B(_11762_),
    .C(_11760_),
    .Y(_11763_)
);

NAND3X1 _21227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11006_),
    .B(_11298_),
    .C(_11299_),
    .Y(_11304_)
);

OAI21X1 _12910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9937_),
    .B(_1380_),
    .C(_1401_),
    .Y(_1412_)
);

AOI21X1 _15382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4878_),
    .B(_4883_),
    .C(_4845_),
    .Y(_4897_)
);

FILL SFILL8680x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6214_),
    .B(_6215_),
    .C(_6213_),
    .Y(_6216_)
);

OAI21X1 _16167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf3),
    .B(_3253__bF$buf3),
    .C(_5755_),
    .Y(_5756_)
);

AND2X2 _12087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4160_),
    .B(_4281_),
    .Y(_4303_)
);

XNOR2X1 _22185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_203_),
    .Y(_445_)
);

NOR3X1 _18733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8562_),
    .B(_8561_),
    .C(_8564_),
    .Y(_8569_)
);

NAND3X1 _18313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8093_),
    .B(_8086_),
    .C(_8098_),
    .Y(_8109_)
);

FILL SFILL13560x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10800_),
    .B(_10805_),
    .C(_10807_),
    .Y(_10965_)
);

FILL SFILL74280x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9890_),
    .B(_9884_),
    .C(_9889_),
    .Y(_9891_)
);

AND2X2 _19518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf4),
    .B(areg_21_bF$buf3),
    .Y(_9430_)
);

AND2X2 _14653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4091_),
    .B(_4096_),
    .Y(_4097_)
);

NAND2X1 _14233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3632_),
    .B(_3637_),
    .Y(_3638_)
);

FILL SFILL74200x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf3),
    .B(_2362__bF$buf5),
    .C(_5411_),
    .Y(_5417_)
);

OAI21X1 _15438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4955_),
    .B(_4954_),
    .C(_4651_),
    .Y(_4958_)
);

OAI21X1 _15018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4496_),
    .B(_4276_),
    .C(_4266_),
    .Y(_4497_)
);

NAND2X1 _20671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10449_),
    .B(_10455_),
    .Y(_10694_)
);

OAI21X1 _20251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_9153_),
    .C(_10218_),
    .Y(_10234_)
);

OAI21X1 _19691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9605_),
    .B(_9608_),
    .C(_9612_),
    .Y(_9621_)
);

NAND3X1 _19271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9158_),
    .B(_9151_),
    .C(_9155_),
    .Y(_9160_)
);

FILL SFILL64280x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11729_),
    .B(_105_),
    .Y(_106_)
);

NAND3X1 _21456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11541_),
    .B(_11546_),
    .C(_11544_),
    .Y(_11555_)
);

NOR3X1 _21036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10833_),
    .B(_10835_),
    .C(_10828_),
    .Y(_11094_)
);

NOR2X1 _15191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_3526_),
    .Y(_4687_)
);

AOI21X1 _13924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3286_),
    .B(_3290_),
    .C(_3257_),
    .Y(_3300_)
);

NAND2X1 _13504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2834_),
    .B(_2839_),
    .Y(_2840_)
);

OAI21X1 _23602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(_1770_),
    .C(_1991_),
    .Y(_1992_)
);

OAI21X1 _16396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5999_),
    .B(_6000_),
    .C(_5745_),
    .Y(_6007_)
);

NAND2X1 _14709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_13_bF$buf3),
    .Y(_4158_)
);

NOR2X1 _18962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8791_),
    .B(_8820_),
    .Y(_8821_)
);

NOR2X1 _18542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7967_),
    .B(_7111_),
    .Y(_8361_)
);

OAI21X1 _18122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7894_),
    .B(_7899_),
    .C(_7888_),
    .Y(_7900_)
);

NAND2X1 _20727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .B(breg_22_bF$buf2),
    .Y(_10755_)
);

OAI21X1 _20307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10287_),
    .B(_10289_),
    .C(_10109_),
    .Y(_10295_)
);

NAND2X1 _23199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1483_),
    .B(_1490_),
    .Y(_1552_)
);

NOR3X1 _19747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9678_),
    .B(_9679_),
    .C(_9680_),
    .Y(_9681_)
);

AOI21X1 _19327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8991_),
    .B(_8996_),
    .C(_8891_),
    .Y(_9221_)
);

OAI21X1 _14882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4347_),
    .B(_4057_),
    .C(_4321_),
    .Y(_4348_)
);

NAND3X1 _14462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3882_),
    .B(_3884_),
    .C(_3883_),
    .Y(_3889_)
);

OAI21X1 _14042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3428_),
    .B(_3426_),
    .C(_3425_),
    .Y(_3429_)
);

NOR3X1 _15667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5195_),
    .B(_5199_),
    .C(_5204_),
    .Y(_5208_)
);

NAND2X1 _15247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4703_),
    .B(_4707_),
    .Y(_4748_)
);

NAND2X1 _20480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf4),
    .B(areg_21_bF$buf0),
    .Y(_10484_)
);

AOI21X1 _20060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10021_),
    .B(_10022_),
    .C(_10007_),
    .Y(_10023_)
);

FILL SFILL8600x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8541_),
    .B(_8605_),
    .Y(_8949_)
);

FILL SFILL13640x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11514_),
    .B(_11509_),
    .Y(_11805_)
);

OAI21X1 _21265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11343_),
    .B(_11342_),
    .C(_11334_),
    .Y(_11344_)
);

OAI21X1 _17813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7508_),
    .B(_7509_),
    .C(_7487_),
    .Y(_7561_)
);

FILL SFILL74280x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2811_),
    .B(_2820_),
    .Y(_3091_)
);

NAND2X1 _13313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_10_bF$buf0),
    .Y(_2631_)
);

NAND2X1 _23831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2215_),
    .Y(_2239_)
);

INVX1 _23411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .Y(_1784_)
);

FILL SFILL74200x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4399_),
    .B(_4404_),
    .C(_4408_),
    .Y(_4409_)
);

NAND2X1 _14518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf4),
    .B(areg_18_bF$buf4),
    .Y(_3950_)
);

INVX2 _18771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8609_),
    .Y(_8611_)
);

NAND3X1 _18351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8144_),
    .B(_8148_),
    .C(_8149_),
    .Y(_8151_)
);

FILL SFILL64280x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10730_),
    .B(_10700_),
    .C(_10738_),
    .Y(_11006_)
);

NOR3X1 _20536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10248_),
    .B(_10210_),
    .C(_10247_),
    .Y(_10546_)
);

NAND3X1 _20116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10065_),
    .B(_10070_),
    .C(_10075_),
    .Y(_10085_)
);

NAND3X1 _19976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9842_),
    .B(_9847_),
    .C(_9849_),
    .Y(_9932_)
);

NAND3X1 _19556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9456_),
    .B(_9424_),
    .C(_9462_),
    .Y(_9472_)
);

FILL SFILL64200x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8948_),
    .B(_9009_),
    .Y(_9011_)
);

NAND3X1 _14691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4135_),
    .B(_4137_),
    .C(_4136_),
    .Y(_4139_)
);

NAND2X1 _14271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf2),
    .B(areg_20_bF$buf3),
    .Y(_3680_)
);

NAND3X1 _15896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5448_),
    .B(_5449_),
    .C(_5444_),
    .Y(_5459_)
);

OAI21X1 _15476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4754_),
    .B(_4761_),
    .C(_4764_),
    .Y(_4998_)
);

AND2X2 _15056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_23_bF$buf3),
    .Y(_4539_)
);

FILL SFILL54200x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11595_),
    .B(_11320_),
    .C(_11580_),
    .Y(_11596_)
);

OAI21X1 _21074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3958__bF$buf2),
    .B(_3781__bF$buf3),
    .C(_11072_),
    .Y(_11136_)
);

XNOR2X1 _17622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7350_),
    .B(_7345_),
    .Y(_7351_)
);

NAND3X1 _17202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6874_),
    .B(_6879_),
    .C(_6886_),
    .Y(_6891_)
);

FILL SFILL74120x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .B(_995_),
    .Y(_1007_)
);

NAND2X1 _22279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf2),
    .B(breg_24_bF$buf2),
    .Y(_547_)
);

OAI21X1 _18827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8670_),
    .B(_8671_),
    .C(_8638_),
    .Y(_8672_)
);

NOR2X1 _18407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7802_),
    .B(_8211_),
    .Y(_8212_)
);

OAI21X1 _13962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3336_),
    .B(_3337_),
    .C(_3322_),
    .Y(_3341_)
);

NAND2X1 _13542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_17_bF$buf2),
    .Y(_2882_)
);

NAND2X1 _13122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2421_),
    .Y(_2422_)
);

AOI21X1 _23640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1906_),
    .B(_2031_),
    .C(_2032_),
    .Y(_2033_)
);

NAND2X1 _23220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1441_),
    .B(_1454_),
    .Y(_1575_)
);

NAND2X1 _14747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4199_),
    .B(_4195_),
    .Y(_4200_)
);

OAI21X1 _14327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3720_),
    .B(_3727_),
    .C(_3592_),
    .Y(_3741_)
);

DFFPOSX1 _24005_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[59]),
    .CLK(clk_bF$buf9),
    .D(_0_[59])
);

FILL SFILL13720x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8328_),
    .B(_8327_),
    .C(_8283_),
    .Y(_8401_)
);

NAND3X1 _18160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7932_),
    .B(_7939_),
    .C(_7940_),
    .Y(_7941_)
);

NAND3X1 _20765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10787_),
    .B(_10780_),
    .C(_10785_),
    .Y(_10797_)
);

NAND2X1 _20345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10317_),
    .B(_10322_),
    .Y(_10336_)
);

NAND3X1 _19785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9689_),
    .B(_9722_),
    .C(_9717_),
    .Y(_9723_)
);

NAND2X1 _19365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9259_),
    .B(_9261_),
    .Y(_9262_)
);

NAND3X1 _14080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3443_),
    .B(_3450_),
    .C(_3452_),
    .Y(_3470_)
);

FILL SFILL44120x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_210_),
    .Y(_352_)
);

AOI21X1 _22911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .B(_1234_),
    .C(_1100_),
    .Y(_1240_)
);

NOR3X1 _15285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4776_),
    .B(_4784_),
    .C(_4786_),
    .Y(_4790_)
);

FILL SFILL3880x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7600_),
    .B(_7601_),
    .C(_7599_),
    .Y(_7603_)
);

NAND3X1 _17431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7086_),
    .B(_7079_),
    .C(_7083_),
    .Y(_7143_)
);

INVX1 _17011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6680_),
    .Y(_6682_)
);

FILL SFILL28840x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_328_),
    .B(_329_),
    .C(_326_),
    .Y(_338_)
);

NAND2X1 _18636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8458_),
    .B(_8462_),
    .Y(_8463_)
);

OAI21X1 _18216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7985_),
    .B(_7990_),
    .C(_7993_),
    .Y(_8003_)
);

OR2X2 _13771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3111_),
    .B(_3130_),
    .Y(_3132_)
);

AND2X2 _13351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2665_),
    .B(_2666_),
    .Y(_2673_)
);

NAND2X1 _14976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_12_bF$buf4),
    .Y(_4451_)
);

OAI21X1 _14556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3943_),
    .B(_3944_),
    .C(_3917_),
    .Y(_3992_)
);

OAI21X1 _14136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3254_),
    .B(_3528_),
    .C(_3530_),
    .Y(_3531_)
);

FILL SFILL18840x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10702_),
    .B(_10727_),
    .C(_10724_),
    .Y(_11048_)
);

AOI21X1 _20574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10574_),
    .B(_10578_),
    .C(_10560_),
    .Y(_10588_)
);

NAND2X1 _20154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10121_),
    .B(_10122_),
    .Y(_10127_)
);

NAND3X1 _16702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6267_),
    .B(_6288_),
    .C(_6289_),
    .Y(_6343_)
);

NAND3X1 _19594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9503_),
    .B(_9496_),
    .C(_9501_),
    .Y(_9514_)
);

NOR2X1 _19174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8657_),
    .B(_8699_),
    .Y(_9053_)
);

NOR2X1 _21779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11899_),
    .B(_11900_),
    .Y(_11907_)
);

NAND2X1 _21359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_24_bF$buf4),
    .Y(_11448_)
);

OAI21X1 _17907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7607_),
    .B(_7662_),
    .C(_7597_),
    .Y(_7663_)
);

NAND2X1 _12622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10090_),
    .B(_10156_),
    .Y(_10167_)
);

NAND2X1 _12202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5552_),
    .B(_5519_),
    .Y(_5563_)
);

OAI21X1 _22720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1025_),
    .C(_951_),
    .Y(_1030_)
);

OAI21X1 _22300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(_565_),
    .C(_558_),
    .Y(_570_)
);

AOI21X1 _15094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4575_),
    .B(_4574_),
    .C(_4573_),
    .Y(_4581_)
);

AOI21X1 _13827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3192_),
    .B(_3193_),
    .C(_3191_),
    .Y(_3194_)
);

NOR3X1 _13407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_2521_),
    .C(_2518_),
    .Y(_2734_)
);

BUFX2 _23925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[43]),
    .Y(y[43])
);

NAND2X1 _23505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_28_bF$buf4),
    .B(breg_28_bF$buf5),
    .Y(_1886_)
);

AOI21X1 _16299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5896_),
    .B(_5899_),
    .C(_5900_),
    .Y(_5901_)
);

NAND2X1 _17660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_18_bF$buf0),
    .Y(_7392_)
);

OAI21X1 _17240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6520_),
    .B(_6535_),
    .C(_6526_),
    .Y(_6932_)
);

OAI21X1 _18865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8708_),
    .B(_8713_),
    .C(_8702_),
    .Y(_8714_)
);

OAI21X1 _18445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8247_),
    .B(_8253_),
    .C(_8223_),
    .Y(_8254_)
);

INVX2 _18025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7792_),
    .Y(_7793_)
);

OAI21X1 _13580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2922_),
    .B(_2921_),
    .C(_2920_),
    .Y(_2923_)
);

INVX1 _13160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .Y(_2463_)
);

FILL SFILL38920x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_3957_),
    .C(_3966_),
    .Y(_4242_)
);

INVX8 _14365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf0),
    .Y(_3781_)
);

DFFPOSX1 _24043_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[1]),
    .CLK(clk_bF$buf1),
    .D(b[1])
);

FILL SFILL3560x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10373_),
    .B(_10374_),
    .C(_10370_),
    .Y(_10378_)
);

NOR3X1 _16931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6590_),
    .B(_6591_),
    .C(_6592_),
    .Y(_6594_)
);

INVX2 _16511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6131_),
    .Y(_6133_)
);

FILL SFILL28840x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11693_),
    .B(_11694_),
    .C(_11647_),
    .Y(_11698_)
);

AOI22X1 _21168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_31_bF$buf3),
    .C(breg_11_bF$buf1),
    .D(areg_30_bF$buf2),
    .Y(_11239_)
);

NOR2X1 _17716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7446_),
    .B(_7447_),
    .Y(_7454_)
);

AOI21X1 _12851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_757_),
    .B(_746_),
    .C(_691_),
    .Y(_768_)
);

OAI21X1 _12431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8052_),
    .B(_8063_),
    .C(_8029_),
    .Y(_8073_)
);

OR2X2 _12011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3460_),
    .B(_3438_),
    .Y(_3471_)
);

OAI21X1 _13636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2783_),
    .B(_2784_),
    .C(_2786_),
    .Y(_2984_)
);

NAND3X1 _13216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2516_),
    .C(_2518_),
    .Y(_2525_)
);

NOR2X1 _23734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7520__bF$buf2),
    .B(_6815__bF$buf3),
    .Y(_2135_)
);

NAND2X1 _23314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf0),
    .B(breg_29_bF$buf1),
    .Y(_1678_)
);

AOI21X1 _18674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8088_),
    .B(_8092_),
    .C(_8096_),
    .Y(_8504_)
);

OAI21X1 _18254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8039_),
    .B(_8044_),
    .C(_7659_),
    .Y(_8045_)
);

NOR3X1 _20859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10588_),
    .B(_10262_),
    .C(_10587_),
    .Y(_10900_)
);

AOI21X1 _20439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10438_),
    .B(_10437_),
    .C(_10431_),
    .Y(_10439_)
);

NAND3X1 _20019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9638_),
    .B(_9965_),
    .C(_9969_),
    .Y(_9979_)
);

NAND3X1 _21800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11890_),
    .B(_21_),
    .C(_20_),
    .Y(_22_)
);

AOI21X1 _19879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9800_),
    .B(_9803_),
    .C(_9813_),
    .Y(_9826_)
);

OAI21X1 _19459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9351_),
    .B(_9350_),
    .C(_9348_),
    .Y(_9365_)
);

OAI22X1 _19039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_5190__bF$buf2),
    .D(_5668__bF$buf4),
    .Y(_8904_)
);

OAI21X1 _14594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4017_),
    .B(_4024_),
    .C(_3779_),
    .Y(_4034_)
);

OR2X2 _14174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3535_),
    .B(_3533_),
    .Y(_3573_)
);

FILL SFILL69080x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _12907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1358_),
    .C(_1314_),
    .D(_1325_),
    .Y(_1380_)
);

NAND3X1 _15799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5350_),
    .B(_5349_),
    .C(_5351_),
    .Y(_5352_)
);

NOR3X1 _15379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4567_),
    .B(_4568_),
    .C(_4565_),
    .Y(_4893_)
);

AOI21X1 _20192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9430_),
    .B(_10148_),
    .C(_9809_),
    .Y(_10169_)
);

NAND3X1 _16740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6378_),
    .B(_6383_),
    .C(_6127_),
    .Y(_6384_)
);

NOR2X1 _16320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5918_),
    .B(_5919_),
    .Y(_5924_)
);

AOI21X1 _21397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11484_),
    .B(_11485_),
    .C(_11476_),
    .Y(_11490_)
);

NAND3X1 _17945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7665_),
    .B(_7704_),
    .C(_7703_),
    .Y(_7705_)
);

NOR2X1 _17525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6821_),
    .B(_7243_),
    .Y(_7244_)
);

AOI21X1 _17105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6764_),
    .B(_6770_),
    .C(_6509_),
    .Y(_6785_)
);

FILL SFILL59080x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10507_),
    .B(_10529_),
    .Y(_10584_)
);

NOR2X1 _12240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5969_),
    .B(_5958_),
    .Y(_0_[8])
);

FILL SFILL3640x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3232_),
    .C(_2981_),
    .Y(_3236_)
);

DFFPOSX1 _23963_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[17]),
    .CLK(clk_bF$buf0),
    .D(_0_[17])
);

NAND3X1 _13445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2772_),
    .B(_2774_),
    .C(_2767_),
    .Y(_2775_)
);

NOR3X1 _13025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2305_),
    .B(_2131_),
    .C(_2311_),
    .Y(_2320_)
);

AOI21X1 _23543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1926_),
    .B(_1927_),
    .C(_1837_),
    .Y(_1928_)
);

NAND3X1 _23123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1464_),
    .B(_1437_),
    .C(_1469_),
    .Y(_1470_)
);

FILL SFILL3560x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28920x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8292_),
    .B(_8295_),
    .C(_8290_),
    .Y(_8296_)
);

NAND3X1 _18063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7834_),
    .B(_7827_),
    .C(_7830_),
    .Y(_7835_)
);

OAI21X1 _20668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10381_),
    .B(_10351_),
    .C(_10389_),
    .Y(_10690_)
);

NAND3X1 _20248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10224_),
    .B(_10215_),
    .C(_10228_),
    .Y(_10229_)
);

OAI21X1 _11931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2453_),
    .B(_2540_),
    .C(_2584_),
    .Y(_2605_)
);

NAND3X1 _19688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9612_),
    .B(_9613_),
    .C(_9616_),
    .Y(_9617_)
);

NAND2X1 _19268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_31_bF$buf0),
    .Y(_9156_)
);

FILL SFILL18920x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9389_),
    .B(_9378_),
    .C(_9356_),
    .Y(_11198_)
);

OAI21X1 _22814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1007_),
    .B(_1005_),
    .C(_997_),
    .Y(_1133_)
);

XNOR2X1 _15188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4682_),
    .B(_4678_),
    .Y(_4683_)
);

OAI21X1 _17754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf2),
    .B(_5921__bF$buf0),
    .C(_7490_),
    .Y(_7496_)
);

NOR2X1 _17334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7027_),
    .B(_7028_),
    .Y(_7036_)
);

NOR3X1 _18959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8770_),
    .B(_7968_),
    .C(_8781_),
    .Y(_8817_)
);

AOI21X1 _18539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8342_),
    .B(_8345_),
    .C(_8347_),
    .Y(_8357_)
);

NAND2X1 _18119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7892_),
    .B(_7890_),
    .Y(_7896_)
);

NOR3X1 _13674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3014_),
    .B(_2773_),
    .C(_3025_),
    .Y(_3026_)
);

NAND2X1 _13254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2565_),
    .Y(_2566_)
);

NAND2X1 _23772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2175_),
    .Y(_2176_)
);

NAND2X1 _23352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1716_),
    .B(_1719_),
    .Y(_1720_)
);

AND2X2 _19900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9471_),
    .B(_9465_),
    .Y(_9849_)
);

NAND2X1 _14879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4343_),
    .B(_4055_),
    .Y(_4344_)
);

AOI21X1 _14459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3884_),
    .B(_3883_),
    .C(_3882_),
    .Y(_3885_)
);

AOI21X1 _14039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3168_),
    .B(_3166_),
    .C(_3173_),
    .Y(_3425_)
);

FILL SFILL43960x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5372_),
    .B(_5373_),
    .Y(_5375_)
);

NAND3X1 _15400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4677_),
    .B(_4764_),
    .C(_4762_),
    .Y(_4916_)
);

OAI21X1 _18292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7682_),
    .B(_7672_),
    .C(_7676_),
    .Y(_8086_)
);

AOI21X1 _20897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10927_),
    .B(_10931_),
    .C(_10915_),
    .Y(_10942_)
);

OAI21X1 _20477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10476_),
    .B(_10480_),
    .C(_10469_),
    .Y(_10481_)
);

AOI21X1 _20057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9654_),
    .B(_9658_),
    .C(_9661_),
    .Y(_10020_)
);

AND2X2 _16605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5854_),
    .B(_6234_),
    .Y(_6236_)
);

NAND3X1 _19497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9402_),
    .B(_9406_),
    .C(_9405_),
    .Y(_9407_)
);

OAI21X1 _19077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf0),
    .B(_5315__bF$buf4),
    .C(_8938_),
    .Y(_8946_)
);

FILL SFILL43880x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_232_),
    .Y(_1794_)
);

INVX8 _12525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf0),
    .Y(_9104_)
);

NOR2X1 _12105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4489_),
    .B(_4466_),
    .Y(_4500_)
);

NAND2X1 _22623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_10686_),
    .Y(_924_)
);

OAI21X1 _22203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_464_),
    .C(_246_),
    .Y(_465_)
);

XNOR2X1 _23828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2213_),
    .B(_2235_),
    .Y(_0_[60])
);

INVX1 _23408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1725_),
    .Y(_1780_)
);

BUFX2 BUFX2_insert420 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf3)
);

BUFX2 BUFX2_insert421 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf2)
);

BUFX2 BUFX2_insert422 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf1)
);

BUFX2 BUFX2_insert423 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(areg_2_bF$buf0)
);

NOR3X1 _17983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7740_),
    .B(_7739_),
    .C(_7742_),
    .Y(_7747_)
);

BUFX2 BUFX2_insert424 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[29]),
    .Y(breg_29_bF$buf4)
);

BUFX2 BUFX2_insert425 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[29]),
    .Y(breg_29_bF$buf3)
);

NAND2X1 _17563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_22_bF$buf1),
    .Y(_7286_)
);

BUFX2 BUFX2_insert426 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[29]),
    .Y(breg_29_bF$buf2)
);

NOR2X1 _17143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6824_),
    .B(_6825_),
    .Y(_6826_)
);

BUFX2 BUFX2_insert427 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[29]),
    .Y(breg_29_bF$buf1)
);

BUFX2 BUFX2_insert428 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[29]),
    .Y(breg_29_bF$buf0)
);

BUFX2 BUFX2_insert429 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .Y(_2586__bF$buf4)
);

FILL SFILL33880x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _18768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8606_),
    .B(_8604_),
    .Y(_8607_)
);

OAI21X1 _18348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8142_),
    .B(_8141_),
    .C(_8138_),
    .Y(_8147_)
);

INVX1 _13483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2816_),
    .Y(_2817_)
);

NAND2X1 _23581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1961_),
    .B(_1967_),
    .Y(_1969_)
);

NAND2X1 _13063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .B(_2335_),
    .Y(_2357_)
);

FILL SFILL23880x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1505_),
    .B(_1506_),
    .C(_1507_),
    .Y(_1512_)
);

NAND2X1 _14688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4091_),
    .Y(_4135_)
);

XNOR2X1 _14268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3675_),
    .B(_3670_),
    .Y(_3676_)
);

FILL SFILL53960x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9555_),
    .B(_9912_),
    .C(_9917_),
    .Y(_10272_)
);

FILL SFILL13880x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6058_),
    .B(_6095_),
    .C(_6098_),
    .Y(_6487_)
);

AOI21X1 _16414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6010_),
    .B(_6015_),
    .C(_5666_),
    .Y(_6027_)
);

FILL SFILL8760x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _17619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7286_),
    .B(_7346_),
    .Y(_7347_)
);

OAI21X1 _12754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11549_),
    .B(_11560_),
    .C(_9948_),
    .Y(_11614_)
);

NAND3X1 _12334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6955_),
    .B(_6999_),
    .C(_6023_),
    .Y(_7020_)
);

NAND2X1 _22852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1127_),
    .B(_1131_),
    .Y(_1175_)
);

OAI21X1 _22432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_702_),
    .B(_472_),
    .C(_714_),
    .Y(_715_)
);

NOR2X1 _22012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf4),
    .B(_6815__bF$buf0),
    .Y(_255_)
);

FILL SFILL29000x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3336_),
    .B(_3337_),
    .C(_3321_),
    .Y(_3338_)
);

NAND2X1 _13539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf3),
    .B(areg_15_bF$buf3),
    .Y(_2878_)
);

FILL SFILL3720x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2402_),
    .B(_2406_),
    .C(_2413_),
    .Y(_2417_)
);

OAI21X1 _23637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(_1903_),
    .C(_2029_),
    .Y(_2030_)
);

XOR2X1 _23217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1571_),
    .B(_1556_),
    .Y(_1572_)
);

FILL SFILL43960x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4366_),
    .Y(_4367_)
);

NAND2X1 _17792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_31_bF$buf4),
    .Y(_7538_)
);

OAI21X1 _17372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6690_),
    .B(_6680_),
    .C(_6685_),
    .Y(_7078_)
);

FILL SFILL23960x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8429_),
    .B(_8436_),
    .C(_8439_),
    .Y(_8859_)
);

OAI21X1 _18577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8397_),
    .B(_8396_),
    .C(_8360_),
    .Y(_8398_)
);

NAND3X1 _18157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7933_),
    .B(_7937_),
    .C(_7936_),
    .Y(_7938_)
);

NAND2X1 _13292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(_2602_),
    .Y(_2607_)
);

FILL FILL74120x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _23390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1759_),
    .B(_1660_),
    .C(_1760_),
    .Y(_1761_)
);

INVX1 _21703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11820_),
    .Y(_11825_)
);

OAI21X1 _14497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_2465__bF$buf0),
    .C(_3919_),
    .Y(_3927_)
);

NOR3X1 _14077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(_3194_),
    .C(_3197_),
    .Y(_3467_)
);

NAND3X1 _22908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .B(_1232_),
    .C(_1231_),
    .Y(_1236_)
);

OAI21X1 _20095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf1),
    .B(_3781__bF$buf1),
    .C(_9702_),
    .Y(_10062_)
);

NAND3X1 _16643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6276_),
    .B(_6277_),
    .C(_6274_),
    .Y(_6278_)
);

NAND3X1 _16223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5779_),
    .B(_5817_),
    .C(_5810_),
    .Y(_5818_)
);

FILL SFILL18920x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7169_),
    .B(_7013_),
    .C(_7598_),
    .Y(_7599_)
);

AOI21X1 _17428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7119_),
    .B(_7128_),
    .C(_7106_),
    .Y(_7139_)
);

AOI21X1 _17008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6321_),
    .B(_6316_),
    .C(_6307_),
    .Y(_6678_)
);

NOR2X1 _12983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2196_),
    .Y(_2207_)
);

NAND3X1 _12563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9488_),
    .B(_9510_),
    .C(_9499_),
    .Y(_9521_)
);

FILL SFILL23880x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3953_),
    .B(_4840_),
    .C(_4884_),
    .Y(_4917_)
);

OR2X2 _22661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_742_),
    .B(_964_),
    .Y(_966_)
);

NOR2X1 _22241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf3),
    .B(_6815__bF$buf0),
    .Y(_506_)
);

FILL SFILL18520x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2898_),
    .B(_2896_),
    .C(_2890_),
    .Y(_3128_)
);

AND2X2 _23866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2265_),
    .B(_2274_),
    .Y(_2276_)
);

INVX8 _13348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf0),
    .Y(_2669_)
);

NAND3X1 _23446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1698_),
    .B(_1717_),
    .C(_1821_),
    .Y(_1822_)
);

NAND3X1 _23026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1340_),
    .C(_1344_),
    .Y(_1364_)
);

FILL SFILL39000x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _17181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6851_),
    .B(_6860_),
    .C(_6861_),
    .Y(_6868_)
);

FILL SFILL13880x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf1),
    .B(_2884__bF$buf1),
    .C(_5478_),
    .Y(_5479_)
);

NAND2X1 _18386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_8189_)
);

FILL SFILL13800x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_161_),
    .B(_163_),
    .C(_162_),
    .Y(_168_)
);

NAND2X1 _21512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11613_),
    .B(_11615_),
    .Y(_11616_)
);

FILL SFILL28680x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg_9_bF$buf3),
    .C(areg_2_bF$buf1),
    .D(breg_10_bF$buf3),
    .Y(_10134_)
);

NAND3X1 _22717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(_1023_),
    .C(_1026_),
    .Y(_1027_)
);

AOI21X1 _16872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6528_),
    .B(_6526_),
    .C(_6519_),
    .Y(_6529_)
);

OAI21X1 _16452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_5318_),
    .C(_6063_),
    .Y(_6067_)
);

AOI21X1 _16032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5148_),
    .B(_5234_),
    .C(_5608_),
    .Y(_5609_)
);

OAI21X1 _17657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf1),
    .B(_2560__bF$buf0),
    .C(_7385_),
    .Y(_7389_)
);

AND2X2 _17237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6863_),
    .B(_6927_),
    .Y(_6929_)
);

NAND3X1 _12792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11690_),
    .B(_111_),
    .C(_100_),
    .Y(_122_)
);

NAND2X1 _12372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg_6_bF$buf2),
    .Y(_7426_)
);

NOR2X1 _22890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_1190_),
    .Y(_1216_)
);

NAND3X1 _22470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_750_),
    .C(_755_),
    .Y(_756_)
);

NAND2X1 _22050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_42_),
    .B(_49_),
    .Y(_296_)
);

NAND3X1 _13997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3360_),
    .B(_3378_),
    .C(_3374_),
    .Y(_3379_)
);

AOI21X1 _13577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2695_),
    .B(_2693_),
    .C(_2691_),
    .Y(_2920_)
);

INVX2 _13157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .Y(_2460_)
);

NAND2X1 _23675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_28_bF$buf3),
    .B(breg_29_bF$buf2),
    .Y(_2071_)
);

OAI21X1 _23255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1610_),
    .B(_1608_),
    .C(_1572_),
    .Y(_1614_)
);

NAND3X1 _19803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9742_),
    .B(_9741_),
    .C(_9736_),
    .Y(_9743_)
);

FILL SFILL54040x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5264_),
    .B(_4969_),
    .C(_5269_),
    .Y(_5270_)
);

NAND3X1 _15303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4793_),
    .B(_4799_),
    .C(_4800_),
    .Y(_4810_)
);

NOR3X1 _18195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7543_),
    .B(_7542_),
    .C(_7544_),
    .Y(_7980_)
);

AOI21X1 _16928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6585_),
    .B(_6586_),
    .C(_6584_),
    .Y(_6590_)
);

OAI21X1 _16508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5992_),
    .B(_6128_),
    .C(_5982_),
    .Y(_6129_)
);

XOR2X1 _21741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11594_),
    .B(_11865_),
    .Y(_0_[43])
);

AND2X2 _21321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11083_),
    .B(_11075_),
    .Y(_11407_)
);

FILL SFILL44040x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10990_),
    .B(_10792_),
    .C(_11022_),
    .Y(_735_)
);

NAND3X1 _12428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7821_),
    .B(_7865_),
    .C(_7887_),
    .Y(_8041_)
);

OAI21X1 _22946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1119_),
    .B(_1275_),
    .C(_1276_),
    .Y(_1277_)
);

NOR2X1 _12008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3405_),
    .B(_3427_),
    .Y(_3438_)
);

AOI21X1 _22526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_578_),
    .C(_817_),
    .Y(_818_)
);

AOI21X1 _22106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_172_),
    .B(_174_),
    .C(_165_),
    .Y(_358_)
);

FILL SFILL8520x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6317_),
    .B(_6318_),
    .Y(_6320_)
);

AOI21X1 _16261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5474_),
    .B(_5479_),
    .C(_5482_),
    .Y(_5860_)
);

FILL SFILL8440x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6039_),
    .B(_5300_),
    .C(_7639_),
    .Y(_7640_)
);

AOI21X1 _17466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7175_),
    .B(_7174_),
    .C(_7173_),
    .Y(_7180_)
);

NAND3X1 _17046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6717_),
    .B(_6719_),
    .C(_6718_),
    .Y(_6720_)
);

OAI21X1 _12181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5310_),
    .B(_5321_),
    .C(_5299_),
    .Y(_5332_)
);

NAND3X1 _13386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2710_),
    .C(_2579_),
    .Y(_2711_)
);

NAND2X1 _23484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1863_),
    .B(_1862_),
    .Y(_1864_)
);

OAI21X1 _23064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1286_),
    .B(_1287_),
    .C(_1292_),
    .Y(_1405_)
);

INVX1 _19612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9533_),
    .Y(_9534_)
);

FILL SFILL38680x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64120x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _15952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3958__bF$buf2),
    .C(_4116__bF$buf3),
    .D(_3402__bF$buf2),
    .Y(_5521_)
);

AOI21X1 _15532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5052_),
    .B(_5053_),
    .C(_5044_),
    .Y(_5060_)
);

NAND3X1 _15112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4362_),
    .B(_4441_),
    .C(_4442_),
    .Y(_4601_)
);

FILL SFILL64040x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9885_),
    .B(_10164_),
    .C(_10163_),
    .Y(_10165_)
);

AOI21X1 _16737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6376_),
    .B(_6375_),
    .C(_6373_),
    .Y(_6381_)
);

INVX8 _16317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf3),
    .Y(_5921_)
);

AOI21X1 _21970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_185_),
    .C(_11826_),
    .Y(_209_)
);

INVX1 _21550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11650_),
    .Y(_11656_)
);

NAND3X1 _21130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11168_),
    .B(_11192_),
    .C(_11196_),
    .Y(_11197_)
);

FILL SFILL28680x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x50 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8994_),
    .Y(_10551_)
);

NAND3X1 _12237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4928_),
    .B(_5859_),
    .C(_5936_),
    .Y(_5947_)
);

OAI21X1 _22755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1068_),
    .B(_1065_),
    .C(_885_),
    .Y(_1069_)
);

NAND2X1 _22335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf4),
    .B(breg_23_bF$buf2),
    .Y(_609_)
);

FILL SFILL54040x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6108_),
    .B(_6107_),
    .C(_6104_),
    .Y(_6109_)
);

AOI21X1 _16070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5648_),
    .B(_5649_),
    .C(_5305_),
    .Y(_5650_)
);

XNOR2X1 _14803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4240_),
    .B(_4261_),
    .Y(_4262_)
);

NAND3X1 _17695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7414_),
    .B(_7419_),
    .C(_7427_),
    .Y(_7431_)
);

NOR2X1 _17275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6967_),
    .B(_6970_),
    .Y(_6971_)
);

OAI21X1 _20821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf3),
    .B(_6300__bF$buf1),
    .C(_10851_),
    .Y(_10859_)
);

NAND2X1 _20401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf3),
    .B(breg_24_bF$buf1),
    .Y(_10398_)
);

AND2X2 _13195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2421_),
    .Y(_2502_)
);

INVX1 _23293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1652_),
    .Y(_1655_)
);

INVX2 _19841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9758_),
    .Y(_9785_)
);

NAND2X1 _19421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_25_bF$buf5),
    .Y(_9324_)
);

NAND3X1 _19001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8861_),
    .B(_8862_),
    .C(_8860_),
    .Y(_8864_)
);

FILL SFILL8920x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _11928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .Y(_2562_)
);

NOR2X1 _21606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11535_),
    .B(_11524_),
    .Y(_11718_)
);

INVX1 _15761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5309_),
    .Y(_5311_)
);

AOI21X1 _15341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4831_),
    .B(_4849_),
    .C(_4850_),
    .Y(_4852_)
);

FILL SFILL34040x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _16966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6608_),
    .B(_6631_),
    .Y(_6632_)
);

OAI22X1 _16546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf0),
    .B(_2560__bF$buf1),
    .C(_549__bF$buf0),
    .D(_2362__bF$buf3),
    .Y(_6171_)
);

OAI21X1 _16126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5708_),
    .B(_5709_),
    .C(_5710_),
    .Y(_5711_)
);

FILL SFILL38760x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_1140_),
    .C(_11417_),
    .Y(_1151_)
);

NAND2X1 _12466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8435_),
    .B(_8446_),
    .Y(_8457_)
);

NAND2X1 _22984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1317_),
    .Y(_1318_)
);

AOI21X1 _12046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3776_),
    .B(_3843_),
    .C(_3471_),
    .Y(_3854_)
);

OR2X2 _22564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_850_),
    .Y(_860_)
);

INVX1 _22144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_151_),
    .Y(_400_)
);

FILL SFILL59160x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _23769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2143_),
    .Y(_2172_)
);

OAI21X1 _23349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(_1715_),
    .C(_1699_),
    .Y(_1716_)
);

OAI21X1 _14612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4050_),
    .B(_3771_),
    .C(_4045_),
    .Y(_4052_)
);

NAND3X1 _17084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6742_),
    .B(_6749_),
    .C(_6752_),
    .Y(_6762_)
);

NAND2X1 _15817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg_22_bF$buf3),
    .Y(_5372_)
);

AOI21X1 _20630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10641_),
    .B(_10648_),
    .C(_10341_),
    .Y(_10649_)
);

NAND3X1 _20210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10174_),
    .B(_10168_),
    .C(_10172_),
    .Y(_10188_)
);

OAI21X1 _18289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7684_),
    .B(_7670_),
    .C(_7694_),
    .Y(_8082_)
);

FILL SFILL49160x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _19650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9574_),
    .B(_9573_),
    .C(_9572_),
    .Y(_9575_)
);

NAND2X1 _19230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .B(_9110_),
    .Y(_9114_)
);

FILL FILL74200x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11749_),
    .B(_11747_),
    .C(_60_),
    .Y(_61_)
);

OAI21X1 _21415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11496_),
    .B(_11500_),
    .C(_11502_),
    .Y(_11510_)
);

NAND3X1 _15990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5557_),
    .B(_5561_),
    .C(_5559_),
    .Y(_5562_)
);

NAND2X1 _15570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5100_),
    .B(_5096_),
    .Y(_5101_)
);

NOR3X1 _15150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4342_),
    .B(_4640_),
    .C(_4054_),
    .Y(_4641_)
);

AOI21X1 _16775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6370_),
    .B(_6377_),
    .C(_6129_),
    .Y(_6422_)
);

FILL SFILL39160x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5906_),
    .B(_5901_),
    .C(_5908_),
    .Y(_5963_)
);

BUFX2 BUFX2_insert390 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[25]),
    .Y(areg_25_bF$buf3)
);

BUFX2 BUFX2_insert391 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[25]),
    .Y(areg_25_bF$buf2)
);

BUFX2 BUFX2_insert392 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[25]),
    .Y(areg_25_bF$buf1)
);

BUFX2 BUFX2_insert393 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[25]),
    .Y(areg_25_bF$buf0)
);

BUFX2 BUFX2_insert394 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf4)
);

FILL SFILL54120x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert395 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf3)
);

BUFX2 BUFX2_insert396 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf2)
);

BUFX2 BUFX2_insert397 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf1)
);

BUFX2 BUFX2_insert398 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(areg_5_bF$buf0)
);

NOR3X1 _12695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10814_),
    .B(_10913_),
    .C(_10924_),
    .Y(_10968_)
);

BUFX2 BUFX2_insert399 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[22]),
    .Y(areg_22_bF$buf4)
);

NOR2X1 _12275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf0),
    .B(_4258__bF$buf3),
    .Y(_6363_)
);

NAND2X1 _22793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1108_),
    .B(_1109_),
    .Y(_1110_)
);

OAI21X1 _22373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_419_),
    .C(_650_),
    .Y(_651_)
);

OAI21X1 _18921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8364_),
    .B(_8772_),
    .C(_8774_),
    .Y(_8776_)
);

NOR3X1 _18501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7946_),
    .B(_7947_),
    .C(_7945_),
    .Y(_8316_)
);

DFFPOSX1 _23998_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[52]),
    .CLK(clk_bF$buf6),
    .D(_0_[52])
);

NAND3X1 _23578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4343_),
    .B(_1964_),
    .C(_1963_),
    .Y(_1965_)
);

NOR3X1 _23158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1506_),
    .B(_1507_),
    .C(_1505_),
    .Y(_1508_)
);

OAI21X1 _19706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9635_),
    .B(_9270_),
    .C(_9619_),
    .Y(_9636_)
);

FILL SFILL69240x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4067_),
    .B(_4148_),
    .C(_4150_),
    .Y(_4304_)
);

OAI21X1 _14421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3829_),
    .B(_3830_),
    .C(_3824_),
    .Y(_3844_)
);

OAI21X1 _14001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3381_),
    .B(_3382_),
    .C(_3380_),
    .Y(_3384_)
);

FILL SFILL34040x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5153_),
    .B(_5161_),
    .C(_5162_),
    .Y(_5163_)
);

NAND3X1 _15206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4683_),
    .B(_4698_),
    .C(_4702_),
    .Y(_4703_)
);

AND2X2 _18098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7414_),
    .B(_7407_),
    .Y(_7873_)
);

OR2X2 _11966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2968_),
    .B(_2705_),
    .Y(_2978_)
);

NAND2X1 _21644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11758_),
    .B(_11759_),
    .Y(_11760_)
);

OAI21X1 _21224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11296_),
    .B(_11300_),
    .C(_11005_),
    .Y(_11301_)
);

FILL SFILL64360x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1155_),
    .C(_1136_),
    .Y(_1171_)
);

NOR2X1 _22429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_710_),
    .Y(_712_)
);

NOR2X1 _22009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf1),
    .B(_7225__bF$buf4),
    .Y(_251_)
);

INVX2 _16584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6130_),
    .Y(_6213_)
);

OAI21X1 _16164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5391_),
    .B(_5380_),
    .C(_5384_),
    .Y(_5753_)
);

INVX1 _17789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7533_),
    .Y(_7534_)
);

OAI21X1 _17369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf2),
    .B(_4541__bF$buf1),
    .C(_7070_),
    .Y(_7074_)
);

INVX2 _12084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4259_),
    .Y(_4270_)
);

AOI21X1 _22182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_432_),
    .C(_366_),
    .Y(_442_)
);

OAI21X1 _18730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8562_),
    .B(_8561_),
    .C(_8564_),
    .Y(_8565_)
);

NOR3X1 _18310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8104_),
    .B(_8100_),
    .C(_8103_),
    .Y(_8105_)
);

NAND3X1 _20915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10904_),
    .B(_10908_),
    .C(_10961_),
    .Y(_10962_)
);

FILL SFILL33960x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .B(_2602_),
    .Y(_2603_)
);

AOI21X1 _23387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1753_),
    .B(_1757_),
    .C(_1661_),
    .Y(_1758_)
);

NAND3X1 _19935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9877_),
    .B(_9870_),
    .C(_9875_),
    .Y(_9888_)
);

AOI21X1 _19515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8641_),
    .B(_9426_),
    .C(_9057_),
    .Y(_9427_)
);

FILL SFILL18760x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4089_),
    .B(_4088_),
    .C(_4073_),
    .Y(_4093_)
);

AOI21X1 _14230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3629_),
    .B(_3628_),
    .C(_3630_),
    .Y(_3634_)
);

FILL SFILL33720x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _15855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf2),
    .B(_2560__bF$buf4),
    .C(_9104__bF$buf3),
    .D(_2362__bF$buf5),
    .Y(_5414_)
);

AOI21X1 _15435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4937_),
    .B(_4943_),
    .C(_4654_),
    .Y(_4955_)
);

NAND3X1 _15015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4491_),
    .B(_4492_),
    .C(_4493_),
    .Y(_4494_)
);

OAI21X1 _21873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11733_),
    .B(_11728_),
    .C(_11737_),
    .Y(_103_)
);

NAND3X1 _21453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11426_),
    .B(_11432_),
    .C(_11434_),
    .Y(_11552_)
);

NAND3X1 _21033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11083_),
    .B(_11087_),
    .C(_11090_),
    .Y(_11091_)
);

OAI21X1 _22658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf3),
    .B(_6427_),
    .C(_961_),
    .Y(_962_)
);

NOR2X1 _22238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf4),
    .B(_7225__bF$buf4),
    .Y(_502_)
);

FILL SFILL69240x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3295_),
    .B(_3050_),
    .C(_3084_),
    .Y(_3297_)
);

NOR3X1 _13501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2829_),
    .B(_2830_),
    .C(_2832_),
    .Y(_2837_)
);

NAND3X1 _16393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5739_),
    .B(_5732_),
    .C(_5736_),
    .Y(_6004_)
);

NAND2X1 _14706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3897_),
    .B(_3903_),
    .Y(_4155_)
);

FILL SFILL29000x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7309_),
    .B(_7313_),
    .C(_7317_),
    .Y(_7324_)
);

AND2X2 _17178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6455_),
    .B(_6514_),
    .Y(_6864_)
);

FILL SFILL59240x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _20724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10745_),
    .B(_10746_),
    .Y(_10752_)
);

NAND3X1 _20304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10104_),
    .B(_10097_),
    .C(_10102_),
    .Y(_10292_)
);

OAI21X1 _13098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2388_),
    .B(_2393_),
    .C(_2394_),
    .Y(_2395_)
);

OAI21X1 _23196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1430_),
    .B(_1410_),
    .C(_1432_),
    .Y(_1549_)
);

AOI21X1 _19744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9282_),
    .B(_9304_),
    .C(_9302_),
    .Y(_9678_)
);

NAND3X1 _19324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9216_),
    .B(_9217_),
    .C(_9215_),
    .Y(_9218_)
);

AOI21X1 _21929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_162_),
    .C(_161_),
    .Y(_164_)
);

INVX2 _21509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11611_),
    .Y(_11612_)
);

FILL FILL74200x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5204_),
    .B(_5199_),
    .C(_5195_),
    .Y(_5205_)
);

AOI21X1 _15244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4726_),
    .B(_4733_),
    .C(_4711_),
    .Y(_4745_)
);

FILL FILL74120x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6522_),
    .B(_6524_),
    .C(_6520_),
    .Y(_6525_)
);

NAND2X1 _16449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6062_),
    .B(_6063_),
    .Y(_6064_)
);

NAND3X1 _16029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5604_),
    .B(_5602_),
    .C(_5603_),
    .Y(_5605_)
);

AOI21X1 _21682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11785_),
    .B(_11793_),
    .C(_11751_),
    .Y(_11802_)
);

NAND2X1 _21262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_27_bF$buf5),
    .Y(_11341_)
);

OAI21X1 _17810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7555_),
    .B(_7556_),
    .C(_7554_),
    .Y(_7557_)
);

FILL SFILL13880x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11701_),
    .B(_34_),
    .C(_78_),
    .Y(_89_)
);

OAI22X1 _12369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5047_),
    .B(_7382_),
    .C(_6374_),
    .D(_6407_),
    .Y(_7393_)
);

XOR2X1 _22887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1212_),
    .B(_1199_),
    .Y(_1213_)
);

INVX1 _22467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_745_),
    .Y(_753_)
);

AND2X2 _22047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_289_),
    .B(_292_),
    .Y(_293_)
);

AOI21X1 _13730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2843_),
    .B(_2861_),
    .C(_2865_),
    .Y(_3087_)
);

NOR2X1 _13310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1936_),
    .B(_2435_),
    .Y(_2627_)
);

OAI21X1 _14935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf2),
    .B(_2586__bF$buf3),
    .C(_4158_),
    .Y(_4406_)
);

AOI21X1 _14515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3693_),
    .B(_3692_),
    .C(_3677_),
    .Y(_3947_)
);

FILL SFILL23960x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10998_),
    .B(_10688_),
    .C(_11002_),
    .Y(_11003_)
);

NAND3X1 _20533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10535_),
    .B(_10539_),
    .C(_10542_),
    .Y(_10543_)
);

OAI21X1 _20113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10080_),
    .B(_10081_),
    .C(_10078_),
    .Y(_10082_)
);

NAND2X1 _19973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9928_),
    .B(_9927_),
    .Y(_9929_)
);

AOI21X1 _19553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9097_),
    .B(_9130_),
    .C(_9139_),
    .Y(_9469_)
);

INVX2 _19133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9007_),
    .Y(_9008_)
);

FILL SFILL69320x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13560x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11598_),
    .B(_11853_),
    .C(_11849_),
    .Y(_11863_)
);

AOI21X1 _21318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11164_),
    .B(_11162_),
    .C(_11151_),
    .Y(_11403_)
);

OAI21X1 _15893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5455_),
    .B(_5450_),
    .C(_5368_),
    .Y(_5456_)
);

OAI21X1 _15473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4985_),
    .B(_4986_),
    .C(_4972_),
    .Y(_4995_)
);

OAI21X1 _15053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4243_),
    .B(_4247_),
    .C(_4246_),
    .Y(_4536_)
);

FILL SFILL13960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6310_),
    .B(_6315_),
    .C(_6313_),
    .Y(_6316_)
);

NOR2X1 _16258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5476_),
    .B(_5850_),
    .Y(_5856_)
);

INVX1 _21491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11590_),
    .Y(_11593_)
);

AND2X2 _21071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10889_),
    .B(_10882_),
    .Y(_11133_)
);

NAND3X1 _12598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8467_),
    .B(_9850_),
    .C(_9861_),
    .Y(_9904_)
);

XNOR2X1 _12178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5080_),
    .B(_5014_),
    .Y(_5299_)
);

NAND3X1 _22696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_981_),
    .B(_1003_),
    .C(_997_),
    .Y(_1004_)
);

OAI21X1 _22276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_299_),
    .C(_307_),
    .Y(_544_)
);

NAND3X1 _18824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8662_),
    .B(_8663_),
    .C(_8664_),
    .Y(_8669_)
);

AOI21X1 _18404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7795_),
    .B(_7800_),
    .C(_7803_),
    .Y(_8209_)
);

FILL FILL74200x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8369_),
    .B(_9173_),
    .Y(_9530_)
);

OAI21X1 _14744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4190_),
    .B(_4191_),
    .C(_4192_),
    .Y(_4197_)
);

NAND3X1 _14324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3587_),
    .B(_3523_),
    .C(_3588_),
    .Y(_3738_)
);

DFFPOSX1 _24002_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[56]),
    .CLK(clk_bF$buf9),
    .D(_0_[56])
);

FILL SFILL74200x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_19_bF$buf3),
    .Y(_5517_)
);

AND2X2 _15529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4723_),
    .B(_4771_),
    .Y(_5056_)
);

OAI21X1 _15109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4595_),
    .B(_4596_),
    .C(_4594_),
    .Y(_4597_)
);

NAND3X1 _20762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10786_),
    .B(_10793_),
    .C(_10740_),
    .Y(_10794_)
);

NAND2X1 _20342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10331_),
    .B(_10333_),
    .Y(_10334_)
);

AOI21X1 _19782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9710_),
    .B(_9704_),
    .C(_9690_),
    .Y(_9720_)
);

OR2X2 _19362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9258_),
    .B(_9251_),
    .Y(_9259_)
);

OAI22X1 _21967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_201_),
    .C(_202_),
    .D(_205_),
    .Y(_206_)
);

NOR2X1 _21547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11651_),
    .B(_11652_),
    .Y(_11653_)
);

NOR3X1 _21127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11186_),
    .B(_11190_),
    .C(_11185_),
    .Y(_11194_)
);

NAND3X1 _12810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_308_),
    .C(_242_),
    .Y(_319_)
);

FILL SFILL23640x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4786_),
    .B(_4784_),
    .C(_4776_),
    .Y(_4787_)
);

OAI21X1 _16487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6091_),
    .B(_6092_),
    .C(_6089_),
    .Y(_6106_)
);

AOI21X1 _16067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5277_),
    .B(_4967_),
    .C(_5281_),
    .Y(_5647_)
);

FILL SFILL23960x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(_334_),
    .C(_327_),
    .Y(_335_)
);

NAND3X1 _18633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8071_),
    .B(_8454_),
    .C(_8455_),
    .Y(_8460_)
);

NAND3X1 _18213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7919_),
    .B(_7922_),
    .C(_7915_),
    .Y(_8000_)
);

AND2X2 _20818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_10855_)
);

FILL SFILL74280x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9771_),
    .B(_9770_),
    .C(_9767_),
    .Y(_9781_)
);

NAND2X1 _19418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8952_),
    .B(_8959_),
    .Y(_9320_)
);

NAND2X1 _14973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4175_),
    .B(_4183_),
    .Y(_4448_)
);

NAND3X1 _14553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3988_),
    .B(_3987_),
    .C(_3985_),
    .Y(_3989_)
);

FILL SFILL13960x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf4),
    .B(breg_19_bF$buf3),
    .Y(_3528_)
);

OAI21X1 _15758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5265_),
    .B(_5268_),
    .C(_5257_),
    .Y(_5307_)
);

NAND2X1 _15338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg_19_bF$buf0),
    .Y(_4848_)
);

NAND3X1 _20991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11029_),
    .B(_11021_),
    .C(_11033_),
    .Y(_11045_)
);

NAND3X1 _20571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10582_),
    .B(_10583_),
    .C(_10581_),
    .Y(_10585_)
);

NOR2X1 _20151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10121_),
    .B(_10122_),
    .Y(_10124_)
);

INVX2 _19591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9484_),
    .Y(_9511_)
);

OAI21X1 _19171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf0),
    .B(_3402__bF$buf1),
    .C(_9045_),
    .Y(_9050_)
);

NAND3X1 _21776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11897_),
    .B(_11903_),
    .C(_11901_),
    .Y(_11904_)
);

XNOR2X1 _21356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11444_),
    .B(_11441_),
    .Y(_11445_)
);

NAND2X1 _17904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7329_),
    .B(_7605_),
    .Y(_7660_)
);

NAND3X1 _15091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4497_),
    .B(_4570_),
    .C(_4576_),
    .Y(_4578_)
);

NAND2X1 _13824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3094_),
    .B(_3090_),
    .Y(_3191_)
);

NAND3X1 _13404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2718_),
    .B(_2721_),
    .C(_2724_),
    .Y(_2731_)
);

BUFX2 _23922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[40]),
    .Y(y[40])
);

NOR2X1 _23502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1793_),
    .B(_1797_),
    .Y(_1883_)
);

OAI21X1 _16296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3961__bF$buf4),
    .C(_5891_),
    .Y(_5898_)
);

OAI21X1 _14609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4047_),
    .B(_4048_),
    .C(_4046_),
    .Y(_4049_)
);

NAND2X1 _18862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8706_),
    .B(_8704_),
    .Y(_8711_)
);

NAND3X1 _18442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8232_),
    .B(_8235_),
    .C(_8245_),
    .Y(_8251_)
);

NOR2X1 _18022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7787_),
    .B(_7789_),
    .Y(_7790_)
);

AOI21X1 _20627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10633_),
    .B(_10634_),
    .C(_10348_),
    .Y(_10646_)
);

OAI21X1 _20207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10183_),
    .B(_10184_),
    .C(_10116_),
    .Y(_10185_)
);

NAND2X1 _23099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .B(areg_27_bF$buf4),
    .Y(_1443_)
);

AOI21X1 _19647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9195_),
    .B(_9191_),
    .C(_9200_),
    .Y(_9572_)
);

NOR2X1 _19227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9109_),
    .B(_9110_),
    .Y(_9111_)
);

FILL SFILL23640x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _14782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_19_bF$buf0),
    .C(breg_4_bF$buf4),
    .D(areg_18_bF$buf4),
    .Y(_4239_)
);

XNOR2X1 _14362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3777_),
    .B(_3535_),
    .Y(_3778_)
);

DFFPOSX1 _24040_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[30]),
    .CLK(clk_bF$buf3),
    .D(a[30])
);

NAND2X1 _15987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5197_),
    .B(_5558_),
    .Y(_5559_)
);

OAI21X1 _15567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5093_),
    .B(_5092_),
    .C(_5094_),
    .Y(_5098_)
);

NAND3X1 _15147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4331_),
    .B(_4638_),
    .C(_4637_),
    .Y(_4639_)
);

AOI21X1 _20380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10362_),
    .B(_10361_),
    .C(_10358_),
    .Y(_10374_)
);

FILL SFILL8600x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11693_),
    .B(_11694_),
    .C(_11692_),
    .Y(_11695_)
);

NAND2X1 _21165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10920_),
    .B(_10922_),
    .Y(_11236_)
);

NAND3X1 _17713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7445_),
    .B(_7450_),
    .C(_7449_),
    .Y(_7451_)
);

FILL SFILL74280x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _18918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_31_bF$buf0),
    .Y(_8772_)
);

NOR3X1 _13633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2961_),
    .B(_2962_),
    .C(_2960_),
    .Y(_2981_)
);

OAI21X1 _13213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_2521_),
    .C(_2518_),
    .Y(_2522_)
);

NAND3X1 _23731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2070_),
    .B(_2075_),
    .C(_2078_),
    .Y(_2132_)
);

NAND2X1 _23311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_25_bF$buf1),
    .B(breg_27_bF$buf1),
    .Y(_1675_)
);

FILL SFILL74200x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4298_),
    .B(_4299_),
    .C(_4297_),
    .Y(_4300_)
);

NOR2X1 _14418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .B(_3839_),
    .Y(_3840_)
);

NOR2X1 _18671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8493_),
    .B(_8494_),
    .Y(_8501_)
);

NAND3X1 _18251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8036_),
    .B(_8037_),
    .C(_7663_),
    .Y(_8042_)
);

FILL SFILL64280x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10896_),
    .B(_10889_),
    .C(_10894_),
    .Y(_10897_)
);

AOI21X1 _20436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10043_),
    .B(_10076_),
    .C(_10080_),
    .Y(_10436_)
);

NOR3X1 _20016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9605_),
    .B(_9608_),
    .C(_9612_),
    .Y(_9976_)
);

AOI21X1 _19876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9451_),
    .B(_9453_),
    .C(_9459_),
    .Y(_9823_)
);

NOR2X1 _19456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8971_),
    .B(_9361_),
    .Y(_9362_)
);

FILL SFILL64200x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _19036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_8901_)
);

NOR3X1 _14591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4029_),
    .B(_3778_),
    .C(_4025_),
    .Y(_4031_)
);

AOI21X1 _14171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3553_),
    .B(_3559_),
    .C(_3539_),
    .Y(_3570_)
);

OAI21X1 _12904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11560_),
    .B(_9707_),
    .C(_11494_),
    .Y(_1347_)
);

OAI21X1 _15796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4986_),
    .B(_4972_),
    .C(_4988_),
    .Y(_5349_)
);

NAND3X1 _15376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4871_),
    .B(_4877_),
    .C(_4880_),
    .Y(_4890_)
);

FILL SFILL58920x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54200x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11181_),
    .B(_11230_),
    .Y(_11487_)
);

OAI21X1 _17942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7701_),
    .B(_7696_),
    .C(_7666_),
    .Y(_7702_)
);

OAI22X1 _17522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf1),
    .B(_5668__bF$buf3),
    .C(_2792_),
    .D(_6050__bF$buf0),
    .Y(_7241_)
);

OAI21X1 _17102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6767_),
    .B(_6768_),
    .C(_6511_),
    .Y(_6782_)
);

FILL SFILL44200x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_897_),
    .C(_728_),
    .Y(_898_)
);

NAND3X1 _22179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_435_),
    .C(_436_),
    .Y(_438_)
);

AOI21X1 _18727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8545_),
    .B(_8551_),
    .C(_8529_),
    .Y(_8562_)
);

OAI21X1 _18307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf0),
    .B(_5668__bF$buf3),
    .C(_8089_),
    .Y(_8102_)
);

AOI21X1 _13862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3230_),
    .B(_3232_),
    .C(_2958_),
    .Y(_3233_)
);

DFFPOSX1 _23960_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[14]),
    .CLK(clk_bF$buf10),
    .D(_0_[14])
);

OAI21X1 _13442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_2763_),
    .C(_2771_),
    .Y(_2772_)
);

NAND3X1 _13022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1902_),
    .B(_2312_),
    .C(_2316_),
    .Y(_2317_)
);

NAND2X1 _23540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1923_),
    .Y(_1924_)
);

NOR2X1 _23120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1462_),
    .B(_1461_),
    .Y(_1466_)
);

NOR3X1 _14647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4088_),
    .B(_4073_),
    .C(_4089_),
    .Y(_4090_)
);

NAND3X1 _14227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3629_),
    .B(_3628_),
    .C(_3630_),
    .Y(_3631_)
);

FILL SFILL13720x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf4),
    .B(_4541__bF$buf1),
    .C(_8291_),
    .Y(_8292_)
);

NOR2X1 _18060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7392_),
    .B(_7440_),
    .Y(_7831_)
);

INVX1 _20665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10686_),
    .Y(_10687_)
);

NOR2X1 _20245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9871_),
    .B(_10225_),
    .Y(_10226_)
);

NOR3X1 _19685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9591_),
    .B(_9597_),
    .C(_9601_),
    .Y(_9614_)
);

INVX4 _19265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_29_bF$buf5),
    .Y(_9153_)
);

FILL SFILL3960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11000_),
    .B(_11044_),
    .C(_10704_),
    .Y(_11165_)
);

OR2X2 _22811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1110_),
    .B(_1124_),
    .Y(_1130_)
);

NOR2X1 _15185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4364_),
    .B(_4679_),
    .Y(_4680_)
);

FILL SFILL3880x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3279_),
    .B(_3284_),
    .C(_3287_),
    .Y(_3293_)
);

NAND2X1 _17751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_24_bF$buf3),
    .Y(_7493_)
);

NAND3X1 _17331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7026_),
    .B(_7030_),
    .C(_7029_),
    .Y(_7033_)
);

FILL SFILL28840x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33800x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8806_),
    .B(_8807_),
    .C(_8744_),
    .Y(_8814_)
);

NAND3X1 _18536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8334_),
    .B(_8349_),
    .C(_8353_),
    .Y(_8354_)
);

OAI21X1 _18116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_4541__bF$buf1),
    .C(_7892_),
    .Y(_7893_)
);

AOI21X1 _13671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3005_),
    .B(_3009_),
    .C(_2991_),
    .Y(_3023_)
);

OAI21X1 _13251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf1),
    .B(_2560__bF$buf4),
    .C(_2561_),
    .Y(_2563_)
);

NAND2X1 _14876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4335_),
    .B(_4341_),
    .Y(_4342_)
);

FILL SFILL13800x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3875_),
    .Y(_3882_)
);

NAND3X1 _14036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3412_),
    .B(_3406_),
    .C(_3410_),
    .Y(_3422_)
);

FILL SFILL18840x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10258_),
    .B(_10932_),
    .C(_10938_),
    .Y(_10939_)
);

NAND2X1 _20474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10473_),
    .B(_10471_),
    .Y(_10478_)
);

NOR2X1 _20054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10009_),
    .B(_10010_),
    .Y(_10017_)
);

NAND3X1 _16602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6228_),
    .B(_6232_),
    .C(_6230_),
    .Y(_6233_)
);

AND2X2 _19494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf5),
    .B(breg_18_bF$buf2),
    .Y(_9404_)
);

OAI21X1 _19074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8942_),
    .B(_8941_),
    .C(_8937_),
    .Y(_8943_)
);

NAND3X1 _21679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11796_),
    .B(_11797_),
    .C(_11795_),
    .Y(_11798_)
);

NAND2X1 _21259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11336_),
    .B(_11337_),
    .Y(_11338_)
);

AOI21X1 _17807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7128_),
    .B(_7106_),
    .C(_7553_),
    .Y(_7554_)
);

NAND3X1 _12942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1685_),
    .B(_1729_),
    .C(_1751_),
    .Y(_1762_)
);

AND2X2 _12522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_10_bF$buf4),
    .Y(_9071_)
);

OAI21X1 _12102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf2),
    .B(_2508_),
    .C(_4466_),
    .Y(_4477_)
);

AOI22X1 _22620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_908_),
    .C(_701_),
    .D(_707_),
    .Y(_920_)
);

NAND3X1 _22200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_457_),
    .C(_249_),
    .Y(_461_)
);

FILL SFILL48920x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3083_),
    .B(_3078_),
    .C(_3082_),
    .Y(_3084_)
);

OAI21X1 _13307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2622_),
    .B(_2623_),
    .C(_2621_),
    .Y(_2624_)
);

XOR2X1 _23825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2232_),
    .B(_2231_),
    .Y(_2233_)
);

OAI21X1 _23405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_),
    .B(_1666_),
    .C(_1690_),
    .Y(_1777_)
);

OAI21X1 _16199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf3),
    .B(_2560__bF$buf1),
    .C(_5786_),
    .Y(_5790_)
);

FILL SFILL13720x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7740_),
    .B(_7739_),
    .C(_7742_),
    .Y(_7743_)
);

INVX1 _17560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7277_),
    .Y(_7282_)
);

NOR2X1 _17140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6430_),
    .B(_6821_),
    .Y(_6822_)
);

INVX2 _18765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8603_),
    .Y(_8604_)
);

NAND3X1 _18345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8124_),
    .B(_8143_),
    .C(_8140_),
    .Y(_8144_)
);

NOR2X1 _13480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2812_),
    .B(_2809_),
    .Y(_2813_)
);

NAND2X1 _13060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11549_),
    .B(_1206_),
    .Y(_2354_)
);

FILL SFILL38920x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4120_),
    .B(_4113_),
    .C(_4099_),
    .Y(_4132_)
);

INVX2 _14265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3672_),
    .Y(_3673_)
);

FILL SFILL3480x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10245_),
    .B(_10209_),
    .C(_10249_),
    .Y(_10269_)
);

FILL SFILL28920x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6475_),
    .B(_6476_),
    .C(_6473_),
    .Y(_6484_)
);

OAI21X1 _16411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6013_),
    .B(_6014_),
    .C(_5667_),
    .Y(_6024_)
);

NAND2X1 _21488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11589_),
    .B(_11584_),
    .Y(_11590_)
);

NAND3X1 _21068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11128_),
    .B(_11127_),
    .C(_11126_),
    .Y(_11129_)
);

AND2X2 _17616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6997_),
    .B(_6990_),
    .Y(_7344_)
);

NAND3X1 _12751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9762_),
    .B(_11538_),
    .C(_11571_),
    .Y(_11582_)
);

NOR3X1 _12331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6933_),
    .B(_6088_),
    .C(_6922_),
    .Y(_6977_)
);

NAND3X1 _13956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3330_),
    .B(_3334_),
    .C(_3322_),
    .Y(_3335_)
);

XNOR2X1 _13536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2874_),
    .B(_2871_),
    .Y(_2875_)
);

OAI21X1 _13116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2411_),
    .C(_2413_),
    .Y(_2414_)
);

AOI21X1 _23634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1898_),
    .B(_1899_),
    .C(_1910_),
    .Y(_2027_)
);

XNOR2X1 _23214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(_1568_),
    .Y(_1569_)
);

FILL SFILL18840x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8839_),
    .B(_8845_),
    .C(_8848_),
    .Y(_8856_)
);

NAND3X1 _18574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8389_),
    .B(_8388_),
    .C(_8387_),
    .Y(_8395_)
);

AND2X2 _18154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_26_bF$buf3),
    .Y(_7935_)
);

AOI21X1 _20759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10789_),
    .B(_10788_),
    .C(_10782_),
    .Y(_10790_)
);

INVX1 _20339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10329_),
    .Y(_10330_)
);

OAI21X1 _21700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11808_),
    .B(_11804_),
    .C(_11820_),
    .Y(_11821_)
);

OAI21X1 _19779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9419_),
    .B(_9421_),
    .C(_9413_),
    .Y(_9716_)
);

XNOR2X1 _19359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8879_),
    .B(_9255_),
    .Y(_0_[35])
);

NAND3X1 _14494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3918_),
    .B(_3923_),
    .C(_3922_),
    .Y(_3924_)
);

AOI21X1 _14074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3443_),
    .B(_3450_),
    .C(_3310_),
    .Y(_3464_)
);

AND2X2 _12807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_166_),
    .Y(_286_)
);

AOI21X1 _22905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(_1231_),
    .C(_1102_),
    .Y(_1233_)
);

NAND3X1 _15699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5235_),
    .B(_5241_),
    .C(_5103_),
    .Y(_5242_)
);

NAND2X1 _15279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_15_bF$buf1),
    .Y(_4783_)
);

NAND3X1 _20092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10051_),
    .B(_10055_),
    .C(_10058_),
    .Y(_10059_)
);

INVX1 _16640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6268_),
    .Y(_6274_)
);

AOI21X1 _16220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5812_),
    .B(_5813_),
    .C(_5806_),
    .Y(_5814_)
);

OR2X2 _21297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11374_),
    .B(_11375_),
    .Y(_11380_)
);

NAND3X1 _17845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7593_),
    .B(_7595_),
    .C(_7594_),
    .Y(_7596_)
);

NOR3X1 _17425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6712_),
    .B(_6709_),
    .C(_6713_),
    .Y(_7136_)
);

NAND3X1 _17005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6665_),
    .B(_6660_),
    .C(_6664_),
    .Y(_6675_)
);

FILL SFILL59080x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf2),
    .B(areg_11_bF$buf1),
    .Y(_2174_)
);

XOR2X1 _12560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8687_),
    .B(_8676_),
    .Y(_9488_)
);

NAND3X1 _12140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4862_),
    .B(_4851_),
    .C(_4873_),
    .Y(_4884_)
);

FILL SFILL38920x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3123_),
    .B(_3124_),
    .C(_3122_),
    .Y(_3125_)
);

NOR2X1 _23863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .B(_2268_),
    .Y(_2273_)
);

NAND2X1 _13345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_16_bF$buf0),
    .Y(_2666_)
);

XNOR2X1 _23443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1818_),
    .B(_1806_),
    .Y(_1819_)
);

NOR2X1 _23023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1345_),
    .Y(_1361_)
);

FILL SFILL3560x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28840x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf1),
    .B(areg_17_bF$buf4),
    .Y(_5476_)
);

AOI21X1 _18383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8009_),
    .B(_8010_),
    .C(_7880_),
    .Y(_8186_)
);

NOR3X1 _20988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11039_),
    .B(_11035_),
    .C(_11038_),
    .Y(_11040_)
);

XNOR2X1 _20568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10559_),
    .B(_10580_),
    .Y(_10581_)
);

NOR2X1 _20148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9774_),
    .B(_10119_),
    .Y(_10120_)
);

AOI21X1 _19588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9495_),
    .B(_9494_),
    .C(_9491_),
    .Y(_9507_)
);

NAND2X1 _19168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9041_),
    .B(_9045_),
    .Y(_9046_)
);

FILL SFILL63960x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10090_),
    .Y(_10101_)
);

AOI21X1 _22714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(_1021_),
    .C(_1018_),
    .Y(_1024_)
);

OAI21X1 _15088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4567_),
    .B(_4568_),
    .C(_4528_),
    .Y(_4574_)
);

BUFX2 _23919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[37]),
    .Y(y[37])
);

NAND2X1 _17654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7384_),
    .B(_7385_),
    .Y(_7386_)
);

INVX2 _17234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6925_),
    .Y(_6926_)
);

FILL SFILL53960x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf4),
    .B(_6300__bF$buf0),
    .C(_8706_),
    .Y(_8707_)
);

AOI21X1 _18439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8240_),
    .B(_8246_),
    .C(_8225_),
    .Y(_8247_)
);

NAND2X1 _18019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_21_bF$buf4),
    .Y(_7786_)
);

AOI21X1 _13994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3367_),
    .B(_3366_),
    .C(_3363_),
    .Y(_3376_)
);

NAND3X1 _13574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2894_),
    .B(_2899_),
    .C(_2870_),
    .Y(_2917_)
);

AOI21X1 _13154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2270_),
    .B(_2288_),
    .C(_2290_),
    .Y(_2457_)
);

NOR2X1 _23672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100__bF$buf3),
    .B(_6815__bF$buf3),
    .Y(_2068_)
);

OAI21X1 _23252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1610_),
    .B(_1608_),
    .C(_1607_),
    .Y(_1611_)
);

NAND3X1 _19800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9730_),
    .B(_9723_),
    .C(_9727_),
    .Y(_9739_)
);

FILL SFILL53880x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4234_),
    .B(_3955_),
    .C(_3980_),
    .Y(_4235_)
);

NOR2X1 _14359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3749_),
    .B(_3752_),
    .Y(_3774_)
);

FILL SFILL3720x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24037_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[27]),
    .CLK(clk_bF$buf6),
    .D(a[27])
);

FILL SFILL43960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5261_),
    .B(_5262_),
    .C(_5258_),
    .Y(_5266_)
);

OAI21X1 _15300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4805_),
    .B(_4801_),
    .C(_4769_),
    .Y(_4806_)
);

OR2X2 _18192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7966_),
    .B(_7970_),
    .Y(_7977_)
);

OAI21X1 _20797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf3),
    .B(_4551__bF$buf4),
    .C(_10831_),
    .Y(_10832_)
);

OAI21X1 _20377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9104__bF$buf0),
    .B(_6050__bF$buf2),
    .C(_10360_),
    .Y(_10371_)
);

NAND3X1 _16925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6585_),
    .B(_6586_),
    .C(_6584_),
    .Y(_6587_)
);

AOI21X1 _16505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6124_),
    .B(_6125_),
    .C(_6123_),
    .Y(_6126_)
);

AOI21X1 _19397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9292_),
    .B(_9296_),
    .C(_9284_),
    .Y(_9297_)
);

FILL SFILL69400x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_571_),
    .B(_604_),
    .C(_494_),
    .Y(_703_)
);

NAND3X1 _12425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7931_),
    .B(_7294_),
    .C(_7997_),
    .Y(_8008_)
);

AND2X2 _22943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1121_),
    .B(_1120_),
    .Y(_1274_)
);

INVX1 _12005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3394_),
    .Y(_3405_)
);

NAND3X1 _22523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_814_),
    .C(_813_),
    .Y(_815_)
);

NAND3X1 _22103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_354_),
    .B(_348_),
    .C(_353_),
    .Y(_355_)
);

NOR2X1 _23728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2092_),
    .B(_2083_),
    .Y(_2128_)
);

NAND2X1 _23308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1669_),
    .B(_1670_),
    .Y(_1671_)
);

FILL SFILL49080x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7633_),
    .B(_7637_),
    .Y(_7638_)
);

NAND3X1 _17463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7170_),
    .B(_7176_),
    .C(_6921_),
    .Y(_7177_)
);

NAND2X1 _17043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6691_),
    .B(_6688_),
    .Y(_6717_)
);

FILL SFILL33880x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8492_),
    .B(_8496_),
    .C(_8495_),
    .Y(_8497_)
);

NAND3X1 _18248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8019_),
    .B(_8024_),
    .C(_7780_),
    .Y(_8037_)
);

OAI21X1 _13383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2701_),
    .B(_2700_),
    .C(_2626_),
    .Y(_2708_)
);

NAND2X1 _23481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .B(_1859_),
    .Y(_1861_)
);

FILL SFILL23880x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1261_),
    .B(_1400_),
    .C(_1398_),
    .Y(_1402_)
);

FILL SFILL54280x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL63960x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4022_),
    .B(_4023_),
    .C(_4021_),
    .Y(_4027_)
);

NAND3X1 _14168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3560_),
    .B(_3565_),
    .C(_3538_),
    .Y(_3566_)
);

FILL SFILL8840x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL53880x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10151_),
    .B(_10150_),
    .C(_10147_),
    .Y(_10162_)
);

NAND3X1 _16734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6370_),
    .B(_6377_),
    .C(_6129_),
    .Y(_6378_)
);

NAND2X1 _16314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_23_bF$buf4),
    .Y(_5918_)
);

FILL SFILL53960x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7693_),
    .B(_7694_),
    .C(_7669_),
    .Y(_7698_)
);

AND2X2 _17519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_28_bF$buf0),
    .Y(_7237_)
);

NAND2X1 _12654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_7_bF$buf1),
    .Y(_10518_)
);

NOR2X1 _12234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5892_),
    .B(_5903_),
    .Y(_5914_)
);

AOI21X1 _22752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1029_),
    .B(_1030_),
    .C(_1028_),
    .Y(_1066_)
);

OAI21X1 _22332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_599_),
    .B(_600_),
    .C(_441_),
    .Y(_606_)
);

FILL SFILL29000x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3223_),
    .B(_3228_),
    .C(_2981_),
    .Y(_3229_)
);

NAND2X1 _13439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_16_bF$buf1),
    .Y(_2768_)
);

DFFPOSX1 _23957_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[11]),
    .CLK(clk_bF$buf2),
    .D(_0_[11])
);

FILL SFILL3720x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_2310_),
    .C(_2306_),
    .Y(_2314_)
);

INVX1 _23537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1915_),
    .Y(_1921_)
);

NAND2X1 _23117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1462_),
    .B(_1461_),
    .Y(_1463_)
);

FILL SFILL74360x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4256_),
    .B(_4255_),
    .C(_4254_),
    .Y(_4257_)
);

OAI21X1 _17692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7423_),
    .B(_7424_),
    .C(_7427_),
    .Y(_7428_)
);

OAI21X1 _17272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf1),
    .B(_2362__bF$buf2),
    .C(_6967_),
    .Y(_6968_)
);

FILL SFILL48920x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _18897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_7520__bF$buf0),
    .C(_4116__bF$buf1),
    .D(_7100__bF$buf2),
    .Y(_8749_)
);

OAI21X1 _18477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7905_),
    .B(_7889_),
    .C(_7896_),
    .Y(_8289_)
);

OAI21X1 _18057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf1),
    .B(_2560__bF$buf0),
    .C(_7823_),
    .Y(_7828_)
);

NOR3X1 _13192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2447_),
    .B(_2480_),
    .C(_2487_),
    .Y(_2499_)
);

FILL FILL74120x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1645_),
    .B(_1651_),
    .Y(_1652_)
);

NOR2X1 _11925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2519__bF$buf2),
    .Y(_2530_)
);

NAND2X1 _21603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11714_),
    .B(_11708_),
    .Y(_11715_)
);

NAND2X1 _14397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf4),
    .B(breg_16_bF$buf1),
    .Y(_3817_)
);

NOR2X1 _22808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1110_),
    .Y(_1126_)
);

OAI21X1 _16963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6627_),
    .B(_6628_),
    .C(_6623_),
    .Y(_6629_)
);

AND2X2 _16543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_16_bF$buf4),
    .Y(_6168_)
);

AOI21X1 _16123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5703_),
    .B(_5702_),
    .C(_5701_),
    .Y(_5708_)
);

FILL SFILL49000x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _17748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7488_),
    .Y(_7489_)
);

AND2X2 _17328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_21_bF$buf2),
    .Y(_7028_)
);

AOI21X1 _12883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1075_),
    .C(_1053_),
    .Y(_1118_)
);

NOR2X1 _12463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7065_),
    .B(_7087_),
    .Y(_8424_)
);

INVX1 _22981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .Y(_1315_)
);

FILL SFILL23880x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3612_),
    .B(_3701_),
    .Y(_3821_)
);

OR2X2 _22561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_851_),
    .Y(_857_)
);

FILL SFILL54280x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_386_),
    .C(_375_),
    .Y(_397_)
);

AOI21X1 _13668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2559_),
    .B(_2775_),
    .C(_2776_),
    .Y(_3019_)
);

OR2X2 _13248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2557_),
    .B(_2558_),
    .Y(_2559_)
);

NAND2X1 _23766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2127_),
    .B(_2150_),
    .Y(_2169_)
);

INVX1 _23346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .Y(_1713_)
);

FILL SFILL8840x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6594_),
    .B(_6589_),
    .C(_6596_),
    .Y(_6759_)
);

INVX4 _15814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_23_bF$buf2),
    .Y(_5369_)
);

NAND2X1 _18286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7750_),
    .B(_7760_),
    .Y(_8079_)
);

FILL SFILL29080x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .B(_52_),
    .C(_50_),
    .Y(_58_)
);

AOI21X1 _21412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11501_),
    .B(_11506_),
    .C(_11471_),
    .Y(_11507_)
);

FILL SFILL29000x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28760x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1696_),
    .B(_1707_),
    .C(_1718_),
    .Y(_1729_)
);

OAI21X1 _12519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7755_),
    .B(_7667_),
    .C(_7700_),
    .Y(_9038_)
);

INVX1 _22617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_915_),
    .Y(_918_)
);

NOR3X1 _16772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6409_),
    .B(_6410_),
    .C(_6405_),
    .Y(_6419_)
);

OAI21X1 _16352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5957_),
    .B(_5959_),
    .C(_5956_),
    .Y(_5960_)
);

BUFX2 BUFX2_insert360 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf3)
);

BUFX2 BUFX2_insert361 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf2)
);

BUFX2 BUFX2_insert362 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf1)
);

BUFX2 BUFX2_insert363 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(breg_0_bF$buf0)
);

AOI21X1 _17977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7729_),
    .B(_7724_),
    .C(_7710_),
    .Y(_7740_)
);

BUFX2 BUFX2_insert364 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[31]),
    .Y(areg_31_bF$buf4)
);

NOR2X1 _17557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6857_),
    .B(_7278_),
    .Y(_7279_)
);

BUFX2 BUFX2_insert365 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[31]),
    .Y(areg_31_bF$buf3)
);

BUFX2 BUFX2_insert366 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[31]),
    .Y(areg_31_bF$buf2)
);

AOI21X1 _17137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6429_),
    .B(_6431_),
    .C(_6818_),
    .Y(_6819_)
);

BUFX2 BUFX2_insert367 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[31]),
    .Y(areg_31_bF$buf1)
);

BUFX2 BUFX2_insert368 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[31]),
    .Y(areg_31_bF$buf0)
);

OAI21X1 _12692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10924_),
    .B(_10913_),
    .C(_10814_),
    .Y(_10935_)
);

BUFX2 BUFX2_insert369 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[28]),
    .Y(areg_28_bF$buf5)
);

NAND3X1 _12272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6297_),
    .B(_6319_),
    .C(_6308_),
    .Y(_6330_)
);

INVX1 _22790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1105_),
    .Y(_1106_)
);

NAND2X1 _22370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_646_),
    .B(_645_),
    .Y(_647_)
);

OAI21X1 _13897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf2),
    .B(_2586__bF$buf0),
    .C(_2796_),
    .Y(_3270_)
);

XNOR2X1 _13477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2809_),
    .B(_2806_),
    .Y(_2810_)
);

DFFPOSX1 _23995_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[49]),
    .CLK(clk_bF$buf6),
    .D(_0_[49])
);

AOI22X1 _23575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3497_),
    .B(_3511_),
    .C(_1961_),
    .D(_1960_),
    .Y(_1962_)
);

OAI21X1 _13057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2350_),
    .B(_2351_),
    .C(_2348_),
    .Y(_2352_)
);

AOI21X1 _23155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1492_),
    .B(_1493_),
    .C(_1491_),
    .Y(_1505_)
);

NAND3X1 _19703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9267_),
    .B(_9626_),
    .C(_9627_),
    .Y(_9633_)
);

FILL SFILL54040x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5154_),
    .B(_5159_),
    .C(_5158_),
    .Y(_5160_)
);

NOR2X1 _15203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4699_),
    .B(_4695_),
    .Y(_4700_)
);

OAI21X1 _18095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7438_),
    .B(_7480_),
    .C(_7472_),
    .Y(_7870_)
);

AOI21X1 _16828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6479_),
    .B(_6474_),
    .C(_6441_),
    .Y(_6480_)
);

OAI21X1 _16408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6018_),
    .B(_6019_),
    .C(_6017_),
    .Y(_6020_)
);

NOR2X1 _11963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2935_),
    .B(_2858_),
    .Y(_2946_)
);

NOR2X1 _21641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2763_),
    .B(_6686__bF$buf2),
    .Y(_11757_)
);

NAND3X1 _21221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11293_),
    .B(_11294_),
    .C(_11009_),
    .Y(_11298_)
);

AOI21X1 _12748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11516_),
    .B(_11505_),
    .C(_9641_),
    .Y(_11549_)
);

OAI21X1 _12328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6922_),
    .B(_6933_),
    .C(_6088_),
    .Y(_6944_)
);

NAND2X1 _22846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1152_),
    .Y(_1168_)
);

INVX1 _22426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .Y(_709_)
);

INVX2 _22006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_247_),
    .Y(_248_)
);

AOI21X1 _16581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5839_),
    .B(_5880_),
    .C(_5877_),
    .Y(_6210_)
);

NAND2X1 _16161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_21_bF$buf0),
    .Y(_5750_)
);

FILL SFILL8440x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_31_bF$buf1),
    .Y(_7531_)
);

NAND2X1 _17366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7069_),
    .B(_7070_),
    .Y(_7071_)
);

OAI21X1 _12081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3821_),
    .B(_3558_),
    .C(_3734_),
    .Y(_4237_)
);

FILL SFILL13800x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10607_),
    .Y(_10959_)
);

NAND2X1 _13286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(_2599_),
    .Y(_2600_)
);

OAI21X1 _23384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1750_),
    .B(_1749_),
    .C(_1612_),
    .Y(_1755_)
);

INVX2 _19932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9857_),
    .Y(_9885_)
);

NAND2X1 _19512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9418_),
    .B(_9423_),
    .Y(_9424_)
);

FILL SFILL64120x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_16_bF$buf2),
    .Y(_5411_)
);

OAI21X1 _15432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4941_),
    .B(_4942_),
    .C(_4656_),
    .Y(_4952_)
);

AND2X2 _15012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4183_),
    .B(_4175_),
    .Y(_4491_)
);

NAND3X1 _20089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10052_),
    .B(_10054_),
    .C(_10053_),
    .Y(_10055_)
);

NAND2X1 _16637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6269_),
    .B(_6270_),
    .Y(_6271_)
);

AOI21X1 _16217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5407_),
    .B(_5429_),
    .C(_5433_),
    .Y(_5811_)
);

AND2X2 _21870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_40_),
    .B(_97_),
    .Y(_99_)
);

OAI21X1 _21450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11543_),
    .B(_11542_),
    .C(_11540_),
    .Y(_11548_)
);

NAND3X1 _21030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11084_),
    .B(_11085_),
    .C(_11086_),
    .Y(_11087_)
);

FILL FILL74040x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_703_),
    .B(_691_),
    .C(_615_),
    .Y(_2142_)
);

NOR3X1 _12557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8939_),
    .B(_9290_),
    .C(_9356_),
    .Y(_9455_)
);

NOR3X1 _12137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3898_),
    .B(_3854_),
    .C(_3920_),
    .Y(_4851_)
);

NAND2X1 _22655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_28_bF$buf3),
    .Y(_959_)
);

INVX2 _22235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .Y(_499_)
);

FILL SFILL54040x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5982_),
    .B(_5987_),
    .C(_5835_),
    .Y(_6000_)
);

NAND2X1 _14703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4146_),
    .B(_4151_),
    .Y(_4152_)
);

FILL SFILL58760x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7314_),
    .B(_7320_),
    .C(_7270_),
    .Y(_7321_)
);

NOR2X1 _17175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6853_),
    .B(_6854_),
    .Y(_6861_)
);

OAI21X1 _15908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5119_),
    .B(_5110_),
    .C(_5115_),
    .Y(_5472_)
);

AND2X2 _20721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10745_),
    .B(_10746_),
    .Y(_10749_)
);

AOI21X1 _20301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10271_),
    .B(_10274_),
    .C(_10205_),
    .Y(_10289_)
);

FILL SFILL44040x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf2),
    .B(_8555_),
    .Y(_2392_)
);

NOR2X1 _23193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1540_),
    .B(_1258_),
    .Y(_1546_)
);

NAND3X1 _19741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9659_),
    .B(_9651_),
    .C(_9664_),
    .Y(_9675_)
);

AOI21X1 _19321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8831_),
    .B(_8828_),
    .C(_9213_),
    .Y(_9215_)
);

NOR2X1 _21926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_120_),
    .B(_125_),
    .Y(_161_)
);

INVX2 _21506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11608_),
    .Y(_11609_)
);

NAND3X1 _15661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5196_),
    .B(_5200_),
    .C(_5198_),
    .Y(_5202_)
);

NAND3X1 _15241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4732_),
    .B(_4718_),
    .C(_4722_),
    .Y(_4742_)
);

OAI21X1 _16866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf0),
    .B(_3253__bF$buf3),
    .C(_6521_),
    .Y(_6522_)
);

INVX1 _16446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6060_),
    .Y(_6061_)
);

NAND2X1 _16026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5600_),
    .B(_5601_),
    .Y(_5602_)
);

AOI21X1 _12786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11855_),
    .B(_11811_),
    .C(_11745_),
    .Y(_56_)
);

FILL SFILL13480x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6220_),
    .B(_7338_),
    .C(_7349_),
    .Y(_7360_)
);

OAI21X1 _22884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_9153_),
    .C(_1209_),
    .Y(_1210_)
);

NAND3X1 _22464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_744_),
    .C(_749_),
    .Y(_750_)
);

OAI21X1 _22044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_285_),
    .C(_284_),
    .Y(_290_)
);

FILL SFILL59160x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686__bF$buf1),
    .B(_7225__bF$buf2),
    .Y(_2064_)
);

XNOR2X1 _23249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1571_),
    .B(_1556_),
    .Y(_1607_)
);

NOR2X1 _14932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4394_),
    .B(_4395_),
    .Y(_4403_)
);

AOI21X1 _14512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .B(_3928_),
    .C(_3933_),
    .Y(_3944_)
);

OAI21X1 _15717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5261_),
    .B(_5262_),
    .C(_5258_),
    .Y(_5263_)
);

XNOR2X1 _20950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10688_),
    .B(_10999_),
    .Y(_0_[40])
);

NAND3X1 _20530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10537_),
    .B(_10538_),
    .C(_10536_),
    .Y(_10539_)
);

AND2X2 _20110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9711_),
    .B(_9704_),
    .Y(_10078_)
);

NOR3X1 _18189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7965_),
    .B(_7972_),
    .C(_7971_),
    .Y(_7973_)
);

INVX1 _19970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9567_),
    .Y(_9925_)
);

NAND3X1 _19550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9425_),
    .B(_9458_),
    .C(_9461_),
    .Y(_9465_)
);

OAI21X1 _19130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8692_),
    .B(_9003_),
    .C(_8829_),
    .Y(_9004_)
);

FILL SFILL54120x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11566_),
    .B(_11569_),
    .C(_11573_),
    .Y(_11860_)
);

NAND3X1 _21315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11393_),
    .B(_11398_),
    .C(_11399_),
    .Y(_11400_)
);

AOI21X1 _15890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .B(_5443_),
    .C(_5404_),
    .Y(_5452_)
);

OAI21X1 _15470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4987_),
    .B(_4990_),
    .C(_4971_),
    .Y(_4991_)
);

AOI22X1 _15050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_20_bF$buf3),
    .C(breg_4_bF$buf3),
    .D(areg_19_bF$buf0),
    .Y(_4532_)
);

FILL SFILL18680x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6311_),
    .B(_6312_),
    .Y(_6313_)
);

NAND3X1 _16255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5849_),
    .B(_5852_),
    .C(_5851_),
    .Y(_5853_)
);

FILL SFILL44040x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9839_),
    .B(_9850_),
    .C(_9861_),
    .Y(_9872_)
);

NOR2X1 _12175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5135_),
    .B(_5157_),
    .Y(_5267_)
);

INVX1 _22693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_860_),
    .Y(_1001_)
);

AOI21X1 _22273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .C(_326_),
    .Y(_541_)
);

AOI21X1 _18821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8663_),
    .B(_8664_),
    .C(_8662_),
    .Y(_8666_)
);

OAI21X1 _18401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf3),
    .B(_3529__bF$buf4),
    .C(_7802_),
    .Y(_8206_)
);

BUFX2 _23898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[16]),
    .Y(y[16])
);

NOR3X1 _23478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1851_),
    .B(_1852_),
    .C(_1853_),
    .Y(_1857_)
);

NAND3X1 _23058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1262_),
    .B(_1394_),
    .C(_1395_),
    .Y(_1398_)
);

NAND3X1 _19606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9525_),
    .B(_9526_),
    .C(_9524_),
    .Y(_9527_)
);

FILL SFILL69240x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4190_),
    .B(_4191_),
    .C(_4192_),
    .Y(_4194_)
);

AOI21X1 _14321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3730_),
    .B(_3733_),
    .C(_3729_),
    .Y(_3735_)
);

INVX1 _15946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5156_),
    .Y(_5514_)
);

OAI21X1 _15526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf2),
    .B(_2362__bF$buf5),
    .C(_5046_),
    .Y(_5053_)
);

AOI21X1 _15106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4200_),
    .B(_4286_),
    .C(_4593_),
    .Y(_4594_)
);

NAND3X1 _21964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_184_),
    .C(_171_),
    .Y(_203_)
);

FILL SFILL59240x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_26_bF$buf4),
    .Y(_11650_)
);

OAI21X1 _21124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11185_),
    .B(_11186_),
    .C(_11190_),
    .Y(_11191_)
);

FILL SFILL24120x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64280x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1061_),
    .B(_1060_),
    .Y(_1062_)
);

NAND3X1 _22329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_598_),
    .C(_601_),
    .Y(_602_)
);

NOR3X1 _16484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5708_),
    .B(_5709_),
    .C(_5710_),
    .Y(_6103_)
);

AOI21X1 _16064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5626_),
    .B(_5633_),
    .C(_5307_),
    .Y(_5644_)
);

FILL SFILL28760x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7413_),
    .B(_7407_),
    .C(_7378_),
    .Y(_7424_)
);

AND2X2 _17269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf2),
    .B(breg_15_bF$buf2),
    .Y(_6964_)
);

NOR2X1 _22082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_116_),
    .B(_331_),
    .Y(_332_)
);

AOI21X1 _18630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8454_),
    .B(_8455_),
    .C(_8071_),
    .Y(_8456_)
);

NAND3X1 _18210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7994_),
    .B(_7995_),
    .C(_7993_),
    .Y(_7996_)
);

FILL SFILL54120x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10498_),
    .B(_10851_),
    .C(_10506_),
    .Y(_10852_)
);

FILL SFILL33960x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .B(_2488_),
    .C(_2494_),
    .Y(_2495_)
);

AOI21X1 _23287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(_1638_),
    .C(_1551_),
    .Y(_1649_)
);

NAND3X1 _19835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9772_),
    .B(_9765_),
    .C(_9777_),
    .Y(_9778_)
);

AND2X2 _19415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9313_),
    .B(_9316_),
    .Y(_9317_)
);

NAND2X1 _14970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4439_),
    .B(_4443_),
    .Y(_4444_)
);

AOI21X1 _14550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3696_),
    .B(_3698_),
    .C(_3984_),
    .Y(_3985_)
);

NOR2X1 _14130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2990_),
    .B(_3251_),
    .Y(_3524_)
);

INVX1 _15755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4999_),
    .Y(_5304_)
);

NAND2X1 _15335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4841_),
    .B(_4844_),
    .Y(_4845_)
);

NAND2X1 _21773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11899_),
    .B(_11900_),
    .Y(_11901_)
);

NAND2X1 _21353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf0),
    .B(breg_22_bF$buf2),
    .Y(_11442_)
);

INVX2 _17901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7655_),
    .Y(_7657_)
);

XOR2X1 _22978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1310_),
    .B(_1299_),
    .Y(_1311_)
);

NAND2X1 _22558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_29_bF$buf1),
    .Y(_853_)
);

INVX1 _22138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_367_),
    .Y(_393_)
);

OAI21X1 _13821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3185_),
    .B(_3186_),
    .C(_3127_),
    .Y(_3188_)
);

OAI21X1 _13401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .B(_2726_),
    .C(_2724_),
    .Y(_2728_)
);

OAI21X1 _16293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf2),
    .B(_3961__bF$buf4),
    .C(_5887_),
    .Y(_5895_)
);

NAND3X1 _14606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3763_),
    .B(_3764_),
    .C(_3517_),
    .Y(_4046_)
);

FILL SFILL29000x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7212_),
    .B(_7209_),
    .Y(_7214_)
);

OAI21X1 _17078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6753_),
    .B(_6754_),
    .C(_6752_),
    .Y(_6755_)
);

FILL SFILL8920x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10304_),
    .B(_9996_),
    .C(_10642_),
    .Y(_10643_)
);

NAND3X1 _20204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10138_),
    .B(_10139_),
    .C(_10137_),
    .Y(_10182_)
);

NAND2X1 _23096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1438_),
    .B(_1439_),
    .Y(_1440_)
);

NOR2X1 _19644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9528_),
    .B(_9568_),
    .Y(_9569_)
);

FILL SFILL3800x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8717_),
    .B(_9107_),
    .Y(_9108_)
);

AOI21X1 _21829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11742_),
    .B(_11743_),
    .C(_11727_),
    .Y(_54_)
);

NAND3X1 _21409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11497_),
    .B(_11498_),
    .C(_11499_),
    .Y(_11503_)
);

FILL FILL74200x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf0),
    .B(areg_24_bF$buf0),
    .Y(_5556_)
);

NOR3X1 _15564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5093_),
    .B(_5092_),
    .C(_5094_),
    .Y(_5095_)
);

NAND3X1 _15144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4339_),
    .B(_4629_),
    .C(_4635_),
    .Y(_4636_)
);

FILL SFILL49240x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6415_),
    .B(_6412_),
    .Y(_6416_)
);

AOI21X1 _16349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5554_),
    .B(_5571_),
    .C(_5955_),
    .Y(_5956_)
);

AOI21X1 _21582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11370_),
    .B(_11404_),
    .C(_11408_),
    .Y(_11692_)
);

OAI21X1 _21162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10912_),
    .B(_11228_),
    .C(_11232_),
    .Y(_11233_)
);

AND2X2 _17710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_22_bF$buf4),
    .Y(_7447_)
);

NAND2X1 _12689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf6),
    .B(areg_12_bF$buf1),
    .Y(_10902_)
);

INVX1 _12269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6121_),
    .Y(_6297_)
);

INVX2 _22787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1102_),
    .Y(_1103_)
);

NAND2X1 _22367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_31_bF$buf2),
    .Y(_644_)
);

OAI21X1 _18915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8767_),
    .B(_8768_),
    .C(_8766_),
    .Y(_8769_)
);

OAI21X1 _13630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2975_),
    .C(_2976_),
    .Y(_2977_)
);

AOI21X1 _13210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .B(_2331_),
    .C(_2333_),
    .Y(_2518_)
);

AOI21X1 _14835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4007_),
    .B(_4010_),
    .C(_4296_),
    .Y(_4297_)
);

OAI21X1 _14415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3836_),
    .B(_3835_),
    .C(_3834_),
    .Y(_3837_)
);

FILL SFILL69000x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23960x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10890_),
    .B(_10892_),
    .C(_10893_),
    .Y(_10894_)
);

AOI21X1 _20433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10417_),
    .B(_10422_),
    .C(_10423_),
    .Y(_10433_)
);

OAI21X1 _20013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9961_),
    .B(_9964_),
    .C(_9966_),
    .Y(_9973_)
);

OAI21X1 _19873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9809_),
    .B(_9810_),
    .C(_9807_),
    .Y(_9820_)
);

OAI21X1 _19453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9357_),
    .B(_9358_),
    .C(_9355_),
    .Y(_9359_)
);

OAI21X1 _19033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8501_),
    .B(_8491_),
    .C(_8495_),
    .Y(_8898_)
);

OAI21X1 _21638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11752_),
    .B(_11475_),
    .C(_11498_),
    .Y(_11753_)
);

NAND3X1 _21218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11012_),
    .B(_11284_),
    .C(_11276_),
    .Y(_11294_)
);

AOI21X1 _12901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11603_),
    .B(_11614_),
    .C(_11592_),
    .Y(_1314_)
);

OAI21X1 _15793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5339_),
    .B(_5340_),
    .C(_5337_),
    .Y(_5346_)
);

OAI21X1 _15373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4842_),
    .B(_4843_),
    .C(_4817_),
    .Y(_4887_)
);

AOI21X1 _16998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6662_),
    .B(_6663_),
    .C(_6661_),
    .Y(_6667_)
);

AOI21X1 _16578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6200_),
    .B(_6204_),
    .C(_6205_),
    .Y(_6206_)
);

NAND2X1 _16158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5436_),
    .B(_5444_),
    .Y(_5746_)
);

OAI21X1 _21391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf3),
    .B(_6686__bF$buf2),
    .C(_11478_),
    .Y(_11484_)
);

OR2X2 _12498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7338_),
    .B(_8753_),
    .Y(_8808_)
);

NAND2X1 _12078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4149_),
    .B(_4182_),
    .Y(_4204_)
);

NAND3X1 _22596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_885_),
    .C(_894_),
    .Y(_895_)
);

AOI21X1 _22176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_161_),
    .C(_434_),
    .Y(_435_)
);

OAI21X1 _18724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8195_),
    .B(_8558_),
    .C(_8219_),
    .Y(_8559_)
);

AOI21X1 _18304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8093_),
    .B(_8098_),
    .C(_8086_),
    .Y(_8099_)
);

OAI21X1 _20909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10953_),
    .B(_10954_),
    .C(_10951_),
    .Y(_10955_)
);

FILL FILL74200x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9869_),
    .B(_9867_),
    .C(_9864_),
    .Y(_9881_)
);

NOR3X1 _19509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9414_),
    .B(_9416_),
    .C(_9415_),
    .Y(_9420_)
);

AOI21X1 _14644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4081_),
    .B(_4086_),
    .C(_4074_),
    .Y(_4087_)
);

NAND3X1 _14224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3621_),
    .B(_3623_),
    .C(_3622_),
    .Y(_3628_)
);

FILL SFILL49240x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5042_),
    .B(_5406_),
    .C(_5051_),
    .Y(_5407_)
);

NAND3X1 _15429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4651_),
    .B(_4944_),
    .C(_4947_),
    .Y(_4948_)
);

AOI21X1 _15009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4205_),
    .B(_4228_),
    .C(_4230_),
    .Y(_4487_)
);

AOI21X1 _20662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10674_),
    .B(_10672_),
    .C(_10683_),
    .Y(_10684_)
);

OAI21X1 _20242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf3),
    .B(_7520__bF$buf3),
    .C(_10222_),
    .Y(_10223_)
);

NOR3X1 _19682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9219_),
    .B(_9226_),
    .C(_9229_),
    .Y(_9611_)
);

OAI21X1 _19262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf1),
    .B(_7520__bF$buf0),
    .C(_9149_),
    .Y(_9150_)
);

INVX2 _21867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .Y(_96_)
);

NAND3X1 _21447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11258_),
    .B(_11541_),
    .C(_11544_),
    .Y(_11545_)
);

INVX1 _21027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11060_),
    .Y(_11084_)
);

OAI21X1 _12710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11121_),
    .B(_11055_),
    .C(_10693_),
    .Y(_11132_)
);

FILL SFILL23640x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4419_),
    .B(_4427_),
    .Y(_4677_)
);

OAI21X1 _13915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3288_),
    .B(_3289_),
    .C(_3287_),
    .Y(_3290_)
);

NOR3X1 _16387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5610_),
    .B(_5611_),
    .C(_5609_),
    .Y(_5997_)
);

FILL SFILL13640x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8779_),
    .B(_8374_),
    .C(_8781_),
    .Y(_8811_)
);

AOI21X1 _18533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8341_),
    .B(_8340_),
    .C(_8336_),
    .Y(_8351_)
);

AND2X2 _18113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf0),
    .B(areg_23_bF$buf2),
    .Y(_7890_)
);

NAND2X1 _20718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf1),
    .B(breg_25_bF$buf0),
    .Y(_10745_)
);

FILL SFILL74280x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _19738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9670_),
    .B(_9666_),
    .C(_9669_),
    .Y(_9671_)
);

AOI21X1 _19318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9209_),
    .B(_9210_),
    .C(_9208_),
    .Y(_9211_)
);

AOI21X1 _14873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4332_),
    .B(_4333_),
    .C(_4042_),
    .Y(_4339_)
);

AND2X2 _14453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf5),
    .B(areg_11_bF$buf0),
    .Y(_3879_)
);

NAND3X1 _14033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3418_),
    .B(_3411_),
    .C(_3395_),
    .Y(_3419_)
);

NAND2X1 _15658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4857_),
    .B(_5197_),
    .Y(_5198_)
);

OAI21X1 _15238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4736_),
    .B(_4737_),
    .C(_4735_),
    .Y(_4738_)
);

OAI21X1 _20891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10929_),
    .B(_10930_),
    .C(_10916_),
    .Y(_10936_)
);

OAI21X1 _20471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf1),
    .B(_3961__bF$buf1),
    .C(_10473_),
    .Y(_10475_)
);

NAND3X1 _20051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10008_),
    .B(_10012_),
    .C(_10011_),
    .Y(_10014_)
);

NAND2X1 _19491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf3),
    .B(breg_20_bF$buf1),
    .Y(_9401_)
);

NAND2X1 _19071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf3),
    .B(breg_24_bF$buf3),
    .Y(_8940_)
);

OAI21X1 _11998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3187_),
    .B(_3209_),
    .C(_3318_),
    .Y(_3329_)
);

OR2X2 _21676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11746_),
    .B(_11750_),
    .Y(_11795_)
);

INVX2 _21256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11334_),
    .Y(_11335_)
);

NAND3X1 _17804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7548_),
    .B(_7550_),
    .C(_7549_),
    .Y(_7551_)
);

NAND3X1 _13724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3059_),
    .B(_3069_),
    .C(_3067_),
    .Y(_3081_)
);

OAI21X1 _13304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2400_),
    .C(_2402_),
    .Y(_2621_)
);

NAND3X1 _23822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_29_bF$buf4),
    .B(breg[31]),
    .C(_2226_),
    .Y(_2230_)
);

OAI21X1 _23402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1773_),
    .C(_1770_),
    .Y(_1774_)
);

NAND2X1 _16196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5785_),
    .B(_5786_),
    .Y(_5787_)
);

NAND3X1 _14929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4393_),
    .B(_4398_),
    .C(_4396_),
    .Y(_4399_)
);

NAND3X1 _14509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3917_),
    .B(_3939_),
    .C(_3934_),
    .Y(_3940_)
);

OAI21X1 _18762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8279_),
    .B(_8600_),
    .C(_8419_),
    .Y(_8601_)
);

AOI21X1 _18342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8134_),
    .B(_8133_),
    .C(_8132_),
    .Y(_8141_)
);

FILL SFILL23720x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10995_),
    .B(_10996_),
    .C(_10994_),
    .Y(_10997_)
);

OR2X2 _20527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10490_),
    .B(_10494_),
    .Y(_10536_)
);

AOI21X1 _20107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9782_),
    .B(_9764_),
    .C(_9787_),
    .Y(_10075_)
);

AOI22X1 _19967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9920_),
    .B(_9921_),
    .C(_9919_),
    .D(_9918_),
    .Y(_9922_)
);

NAND3X1 _19547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9457_),
    .B(_9458_),
    .C(_9461_),
    .Y(_9462_)
);

NAND3X1 _19127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8999_),
    .B(_9000_),
    .C(_8998_),
    .Y(_9001_)
);

NAND3X1 _14682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4106_),
    .B(_4111_),
    .C(_4108_),
    .Y(_4129_)
);

NOR2X1 _14262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf1),
    .B(_2465__bF$buf0),
    .Y(_3670_)
);

FILL SFILL8680x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5137_),
    .B(_5143_),
    .C(_5145_),
    .Y(_5449_)
);

NAND2X1 _15467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4982_),
    .B(_4984_),
    .Y(_4988_)
);

NOR2X1 _15047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf1),
    .B(_3146__bF$buf0),
    .Y(_4529_)
);

INVX1 _20280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10264_),
    .Y(_10265_)
);

FILL SFILL8600x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11319_),
    .B(_11581_),
    .C(_11580_),
    .Y(_11587_)
);

AND2X2 _21065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10794_),
    .B(_10786_),
    .Y(_11126_)
);

NAND2X1 _17613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7335_),
    .B(_7340_),
    .Y(_7341_)
);

FILL SFILL74280x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8248_),
    .B(_8644_),
    .C(_8232_),
    .Y(_8662_)
);

NOR2X1 _13953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3062_),
    .B(_3331_),
    .Y(_3332_)
);

NAND2X1 _13533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_13_bF$buf1),
    .Y(_2872_)
);

AOI21X1 _13113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2397_),
    .B(_2401_),
    .C(_2386_),
    .Y(_2411_)
);

OAI21X1 _23631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(_2005_),
    .C(_2022_),
    .Y(_2024_)
);

OAI21X1 _23211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300__bF$buf3),
    .B(_5668__bF$buf1),
    .C(_1417_),
    .Y(_1566_)
);

FILL SFILL43800x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3880x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4185_),
    .B(_4186_),
    .C(_4184_),
    .Y(_4190_)
);

NOR3X1 _14318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3707_),
    .B(_3714_),
    .C(_3716_),
    .Y(_3731_)
);

NAND3X1 _18991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8849_),
    .B(_8850_),
    .C(_8848_),
    .Y(_8853_)
);

OAI21X1 _18571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8384_),
    .B(_8390_),
    .C(_8332_),
    .Y(_8392_)
);

NAND2X1 _18151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_24_bF$buf1),
    .Y(_7932_)
);

FILL SFILL64280x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10393_),
    .B(_10428_),
    .C(_10432_),
    .Y(_10787_)
);

AOI21X1 _20336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10311_),
    .B(_10316_),
    .C(_9993_),
    .Y(_10327_)
);

NAND3X1 _19776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9709_),
    .B(_9697_),
    .C(_9701_),
    .Y(_9713_)
);

NAND3X1 _19356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8883_),
    .B(_9243_),
    .C(_9238_),
    .Y(_9253_)
);

FILL SFILL64200x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf1),
    .B(areg_15_bF$buf1),
    .Y(_3921_)
);

NAND3X1 _14071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3305_),
    .B(_3250_),
    .C(_3306_),
    .Y(_3461_)
);

NAND2X1 _12804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf3),
    .B(areg_7_bF$buf0),
    .Y(_253_)
);

NOR3X1 _22902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1225_),
    .B(_1103_),
    .C(_1229_),
    .Y(_1230_)
);

FILL SFILL54200x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5231_),
    .B(_5232_),
    .C(_5150_),
    .Y(_5239_)
);

NAND2X1 _15276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4778_),
    .B(_4779_),
    .Y(_4780_)
);

AOI22X1 _21294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_25_bF$buf2),
    .C(areg_18_bF$buf2),
    .D(breg_24_bF$buf0),
    .Y(_11377_)
);

NAND2X1 _17842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7590_),
    .B(_7592_),
    .Y(_7593_)
);

NAND3X1 _17422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7118_),
    .B(_7121_),
    .C(_7115_),
    .Y(_7133_)
);

OAI21X1 _17002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6671_),
    .B(_6666_),
    .C(_6652_),
    .Y(_6672_)
);

NAND3X1 _22499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_787_),
    .C(_785_),
    .Y(_788_)
);

AOI21X1 _22079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_323_),
    .C(_321_),
    .Y(_328_)
);

AOI21X1 _18627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8448_),
    .B(_8452_),
    .C(_8072_),
    .Y(_8453_)
);

AOI21X1 _18207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7511_),
    .B(_7557_),
    .C(_7992_),
    .Y(_7993_)
);

OAI21X1 _13762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2638_),
    .B(_2849_),
    .C(_2848_),
    .Y(_3122_)
);

NOR2X1 _23860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8773_),
    .B(_7225__bF$buf1),
    .Y(_2269_)
);

NAND2X1 _13342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf2),
    .B(areg_14_bF$buf4),
    .Y(_2663_)
);

XOR2X1 _23440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1814_),
    .B(_1810_),
    .Y(_1815_)
);

XOR2X1 _23020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(_1350_),
    .Y(_1357_)
);

NAND3X1 _14967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4431_),
    .B(_4437_),
    .C(_4427_),
    .Y(_4441_)
);

AOI21X1 _14547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3981_),
    .B(_3980_),
    .C(_3979_),
    .Y(_3982_)
);

INVX2 _14127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3520_),
    .Y(_3521_)
);

OAI21X1 _18380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8176_),
    .B(_8175_),
    .C(_8173_),
    .Y(_8182_)
);

OAI21X1 _20985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf1),
    .B(_5668__bF$buf5),
    .C(_11025_),
    .Y(_11037_)
);

OAI21X1 _20565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10577_),
    .B(_10576_),
    .C(_10575_),
    .Y(_10578_)
);

OAI21X1 _20145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9776_),
    .B(_9766_),
    .C(_9770_),
    .Y(_10117_)
);

OAI21X1 _19585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf4),
    .B(_6686__bF$buf3),
    .C(_9493_),
    .Y(_9504_)
);

NAND2X1 _19165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf1),
    .B(areg_18_bF$buf5),
    .Y(_9043_)
);

FILL SFILL44120x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8566_),
    .B(_8610_),
    .C(_10057_),
    .Y(_10068_)
);

NAND3X1 _22711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1011_),
    .B(_1004_),
    .C(_1008_),
    .Y(_1021_)
);

NAND3X1 _15085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4499_),
    .B(_4515_),
    .C(_4520_),
    .Y(_4571_)
);

FILL SFILL43800x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3126_),
    .B(_3180_),
    .C(_3179_),
    .Y(_3184_)
);

BUFX2 _23916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[34]),
    .Y(y[34])
);

INVX1 _17651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7381_),
    .Y(_7383_)
);

NAND2X1 _17231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6577_),
    .B(_6583_),
    .Y(_6923_)
);

AND2X2 _18856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_25_bF$buf4),
    .Y(_8704_)
);

AND2X2 _18436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7838_),
    .B(_7884_),
    .Y(_8244_)
);

NAND2X1 _18016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7407_),
    .B(_7414_),
    .Y(_7783_)
);

OAI21X1 _13991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3135_),
    .B(_3137_),
    .C(_3132_),
    .Y(_3373_)
);

AOI21X1 _13571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2856_),
    .B(_2861_),
    .C(_2843_),
    .Y(_2914_)
);

AND2X2 _13151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .B(_2451_),
    .Y(_2454_)
);

OAI21X1 _14776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4230_),
    .B(_4231_),
    .C(_4205_),
    .Y(_4232_)
);

FILL SFILL13800x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3762_),
    .B(_3765_),
    .C(_3494_),
    .Y(_3771_)
);

DFFPOSX1 _24034_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[24]),
    .CLK(clk_bF$buf9),
    .D(a[24])
);

FILL SFILL58920x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _20794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10822_),
    .Y(_10829_)
);

OAI21X1 _20374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10367_),
    .B(_10366_),
    .C(_10357_),
    .Y(_10368_)
);

OR2X2 _16922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6539_),
    .B(_6544_),
    .Y(_6584_)
);

NAND2X1 _16502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5718_),
    .B(_5725_),
    .Y(_6123_)
);

NOR2X1 _19394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8907_),
    .B(_9293_),
    .Y(_9294_)
);

FILL SFILL44200x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_223_),
    .C(_11884_),
    .Y(_240_)
);

OAI21X1 _21579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11680_),
    .B(_11681_),
    .C(_11677_),
    .Y(_11688_)
);

INVX1 _21159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf2),
    .Y(_11229_)
);

NAND2X1 _17707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_20_bF$buf2),
    .Y(_7444_)
);

NAND3X1 _12842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_615_),
    .C(_659_),
    .Y(_680_)
);

NOR3X1 _12422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7898_),
    .B(_7909_),
    .C(_7887_),
    .Y(_7975_)
);

NAND2X1 _22940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1111_),
    .B(_1123_),
    .Y(_1270_)
);

NAND3X1 _12002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3361_),
    .B(_3033_),
    .C(_3000_),
    .Y(_3372_)
);

AND2X2 _22520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_567_),
    .B(_559_),
    .Y(_811_)
);

FILL SFILL69480x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_339_),
    .C(_344_),
    .Y(_351_)
);

FILL SFILL48920x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _13627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2751_),
    .B(_2974_),
    .Y(_0_[17])
);

NAND3X1 _13207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2501_),
    .B(_2505_),
    .C(_2509_),
    .Y(_2515_)
);

AOI21X1 _23725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2082_),
    .C(_2124_),
    .Y(_2125_)
);

OR2X2 _23305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1562_),
    .Y(_1668_)
);

NAND2X1 _16099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_25_bF$buf3),
    .Y(_5681_)
);

FILL SFILL13720x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6843_),
    .B(_7622_),
    .C(_7628_),
    .Y(_7634_)
);

OAI21X1 _17460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7167_),
    .B(_7168_),
    .C(_7015_),
    .Y(_7174_)
);

AOI21X1 _17040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6701_),
    .B(_6699_),
    .C(_6696_),
    .Y(_6713_)
);

AND2X2 _18665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg_27_bF$buf3),
    .Y(_8494_)
);

NOR3X1 _18245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7600_),
    .B(_7601_),
    .C(_7599_),
    .Y(_8034_)
);

NAND3X1 _13380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2619_),
    .C(_2612_),
    .Y(_2704_)
);

FILL SFILL38920x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4022_),
    .B(_4023_),
    .C(_4021_),
    .Y(_4024_)
);

NAND3X1 _14165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3551_),
    .B(_3549_),
    .C(_3545_),
    .Y(_3563_)
);

FILL SFILL3560x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9485_),
    .B(_10157_),
    .C(_10158_),
    .D(_9857_),
    .Y(_10159_)
);

FILL SFILL28920x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6367_),
    .B(_6368_),
    .C(_6219_),
    .Y(_6375_)
);

OAI21X1 _16311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5913_),
    .B(_5573_),
    .C(_5567_),
    .Y(_5915_)
);

NAND2X1 _21388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_26_bF$buf4),
    .Y(_11480_)
);

NAND3X1 _17936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7669_),
    .B(_7693_),
    .C(_7694_),
    .Y(_7695_)
);

OAI21X1 _17516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6826_),
    .B(_6820_),
    .C(_6829_),
    .Y(_7234_)
);

OAI21X1 _12651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8753_),
    .B(_10452_),
    .C(_10474_),
    .Y(_10485_)
);

NAND3X1 _12231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4051_),
    .B(_4862_),
    .C(_4873_),
    .Y(_5881_)
);

NAND3X1 _13856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2984_),
    .B(_3219_),
    .C(_3221_),
    .Y(_3226_)
);

NAND2X1 _13436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf1),
    .B(breg_15_bF$buf1),
    .Y(_2765_)
);

DFFPOSX1 _23954_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[8]),
    .CLK(clk_bF$buf2),
    .D(_0_[8])
);

NOR3X1 _13016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_2310_),
    .C(_2306_),
    .Y(_2311_)
);

NOR2X1 _23534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_1916_),
    .Y(_1918_)
);

NAND2X1 _23114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1455_),
    .Y(_1460_)
);

FILL SFILL18840x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _18894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8745_),
    .Y(_8746_)
);

NAND2X1 _18474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_21_bF$buf3),
    .Y(_8286_)
);

NAND2X1 _18054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_7825_)
);

NOR3X1 _20659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10649_),
    .B(_10653_),
    .C(_10656_),
    .Y(_10680_)
);

AND2X2 _20239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf3),
    .B(areg_29_bF$buf3),
    .Y(_10219_)
);

OAI21X1 _11922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_2453_),
    .C(_2486_),
    .Y(_2497_)
);

NAND3X1 _21600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11700_),
    .B(_11706_),
    .C(_11696_),
    .Y(_11711_)
);

OAI21X1 _19679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9591_),
    .B(_9597_),
    .C(_9601_),
    .Y(_9607_)
);

AND2X2 _19259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf5),
    .B(areg_29_bF$buf3),
    .Y(_9146_)
);

NAND2X1 _14394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3812_),
    .B(_3813_),
    .Y(_3814_)
);

DFFPOSX1 _24072_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[30]),
    .CLK(clk_bF$buf4),
    .D(b[30])
);

AOI21X1 _12707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11077_),
    .B(_11088_),
    .C(_11011_),
    .Y(_11099_)
);

XNOR2X1 _22805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1122_),
    .B(_1112_),
    .Y(_1123_)
);

NAND3X1 _15599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5122_),
    .B(_5117_),
    .C(_5120_),
    .Y(_5133_)
);

XNOR2X1 _15179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4672_),
    .B(_4671_),
    .Y(_4673_)
);

OAI21X1 _16960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_3958__bF$buf3),
    .C(_6229_),
    .Y(_6625_)
);

OAI21X1 _16540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5781_),
    .B(_6163_),
    .C(_5789_),
    .Y(_6164_)
);

NAND3X1 _16120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5703_),
    .B(_5701_),
    .C(_5702_),
    .Y(_5704_)
);

OAI21X1 _21197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10909_),
    .B(_10951_),
    .C(_11270_),
    .Y(_11271_)
);

AND2X2 _17745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_24_bF$buf3),
    .Y(_7486_)
);

NAND2X1 _17325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf0),
    .B(areg_19_bF$buf5),
    .Y(_7025_)
);

FILL SFILL59080x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1064_),
    .C(_1075_),
    .Y(_1086_)
);

NOR2X1 _12460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7109_),
    .B(_8359_),
    .Y(_8391_)
);

AOI21X1 _12040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2749_),
    .B(_3787_),
    .C(_2924_),
    .Y(_3788_)
);

FILL SFILL38920x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3003_),
    .B(_2999_),
    .C(_2995_),
    .Y(_3016_)
);

OAI21X1 _13245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2555_),
    .B(_2373_),
    .C(_2506_),
    .Y(_2556_)
);

INVX1 _23763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2134_),
    .Y(_2166_)
);

OAI21X1 _23343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1618_),
    .C(_1709_),
    .Y(_1710_)
);

FILL SFILL3560x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49080x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28920x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5360_),
    .B(_5364_),
    .Y(_5366_)
);

INVX2 _18283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8075_),
    .Y(_8076_)
);

NAND3X1 _20888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10927_),
    .B(_10931_),
    .C(_10915_),
    .Y(_10932_)
);

AND2X2 _20468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf4),
    .B(areg_21_bF$buf0),
    .Y(_10471_)
);

AND2X2 _20048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf1),
    .B(breg_27_bF$buf2),
    .Y(_10010_)
);

NOR2X1 _19488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9395_),
    .B(_9396_),
    .Y(_9397_)
);

OAI21X1 _19068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8535_),
    .B(_8530_),
    .C(_8538_),
    .Y(_8936_)
);

INVX1 _12936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1533_),
    .Y(_1696_)
);

AND2X2 _12516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7591_),
    .B(_8983_),
    .Y(_9005_)
);

NAND2X1 _22614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_914_),
    .Y(_915_)
);

XOR2X1 _23819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2222_),
    .B(_2225_),
    .Y(_2226_)
);

BUFX2 BUFX2_insert330 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf1)
);

BUFX2 BUFX2_insert331 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(breg_6_bF$buf0)
);

BUFX2 BUFX2_insert332 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .Y(_2287__bF$buf3)
);

BUFX2 BUFX2_insert333 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .Y(_2287__bF$buf2)
);

OAI21X1 _17974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7351_),
    .B(_7736_),
    .C(_7375_),
    .Y(_7737_)
);

BUFX2 BUFX2_insert334 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .Y(_2287__bF$buf1)
);

NAND2X1 _17554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_26_bF$buf1),
    .Y(_7276_)
);

BUFX2 BUFX2_insert335 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .Y(_2287__bF$buf0)
);

NOR2X1 _17134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf2),
    .B(_6815__bF$buf1),
    .Y(_6816_)
);

BUFX2 BUFX2_insert336 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf5)
);

BUFX2 BUFX2_insert337 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf4)
);

BUFX2 BUFX2_insert338 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf3)
);

BUFX2 BUFX2_insert339 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(breg_15_bF$buf2)
);

FILL SFILL74440x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8595_),
    .B(_8594_),
    .C(_8596_),
    .Y(_8597_)
);

AOI21X1 _18339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7784_),
    .B(_8136_),
    .C(_7787_),
    .Y(_8137_)
);

OAI21X1 _13894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf3),
    .B(_2362__bF$buf0),
    .C(_2996_),
    .Y(_3267_)
);

NAND2X1 _13474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf4),
    .B(breg_10_bF$buf3),
    .Y(_2807_)
);

DFFPOSX1 _23992_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[46]),
    .CLK(clk_bF$buf8),
    .D(_0_[46])
);

OAI21X1 _23572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2975_),
    .B(_2752_),
    .C(_1958_),
    .Y(_1959_)
);

OR2X2 _13054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .B(_2348_),
    .Y(_2349_)
);

NOR2X1 _23152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1353_),
    .Y(_1502_)
);

INVX2 _19700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9629_),
    .Y(_9630_)
);

OAI21X1 _14679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4124_),
    .B(_4123_),
    .C(_4122_),
    .Y(_4125_)
);

NAND2X1 _14259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3661_),
    .B(_3665_),
    .Y(_3666_)
);

FILL SFILL3720x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_19_bF$buf2),
    .Y(_5156_)
);

OAI21X1 _15200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf4),
    .B(_3526_),
    .C(_4695_),
    .Y(_4696_)
);

OAI21X1 _18092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7864_),
    .B(_7856_),
    .C(_7866_),
    .Y(_7867_)
);

AOI21X1 _20697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10720_),
    .B(_10721_),
    .C(_10706_),
    .Y(_10722_)
);

NAND2X1 _20277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10260_),
    .B(_10256_),
    .Y(_10262_)
);

AOI21X1 _16825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6152_),
    .B(_6153_),
    .C(_6137_),
    .Y(_6477_)
);

INVX2 _16405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5666_),
    .Y(_6017_)
);

XNOR2X1 _11960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2847_),
    .B(_2902_),
    .Y(_2913_)
);

AOI21X1 _19297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9185_),
    .B(_9187_),
    .C(_9141_),
    .Y(_9188_)
);

NAND3X1 _12745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11406_),
    .B(_11450_),
    .C(_11362_),
    .Y(_11516_)
);

NAND3X1 _12325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6099_),
    .B(_6900_),
    .C(_6834_),
    .Y(_6911_)
);

OAI21X1 _22843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1163_),
    .C(_1161_),
    .Y(_1165_)
);

NAND3X1 _22423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(_684_),
    .C(_696_),
    .Y(_706_)
);

AOI21X1 _22003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_212_),
    .C(_11888_),
    .Y(_245_)
);

AND2X2 _23628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2018_),
    .B(_2007_),
    .Y(_2020_)
);

NAND2X1 _23208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_23_bF$buf4),
    .B(breg_29_bF$buf1),
    .Y(_1562_)
);

FILL SFILL49080x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7108_),
    .B(_7113_),
    .C(_7112_),
    .Y(_7528_)
);

INVX1 _17363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7067_),
    .Y(_7068_)
);

FILL SFILL49000x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8432_),
    .B(_8434_),
    .C(_8847_),
    .Y(_8848_)
);

OAI21X1 _18568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7973_),
    .B(_7971_),
    .C(_8382_),
    .Y(_8388_)
);

OAI21X1 _18148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7562_),
    .B(_7927_),
    .C(_7552_),
    .Y(_7928_)
);

OAI21X1 _13283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf3),
    .B(_6044__bF$buf2),
    .C(_2393_),
    .Y(_2597_)
);

NOR3X1 _23381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1749_),
    .C(_1750_),
    .Y(_1752_)
);

FILL SFILL23880x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54280x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3640_),
    .B(_3916_),
    .C(_3648_),
    .Y(_3917_)
);

OAI21X1 _14068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3456_),
    .B(_3455_),
    .C(_3452_),
    .Y(_3457_)
);

FILL SFILL23800x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL73960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10045_),
    .Y(_10052_)
);

FILL SFILL13880x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_3958__bF$buf1),
    .Y(_6268_)
);

AOI21X1 _16214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5789_),
    .B(_5794_),
    .C(_5797_),
    .Y(_5808_)
);

NAND3X1 _17839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7583_),
    .B(_7434_),
    .C(_7588_),
    .Y(_7589_)
);

NAND3X1 _17419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7119_),
    .B(_7128_),
    .C(_7106_),
    .Y(_7129_)
);

OAI21X1 _12974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2034_),
    .B(_2045_),
    .C(_1990_),
    .Y(_2109_)
);

NAND3X1 _12554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9367_),
    .B(_9411_),
    .C(_8709_),
    .Y(_9422_)
);

AOI21X1 _12134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4642_),
    .B(_4686_),
    .C(_4072_),
    .Y(_4818_)
);

INVX1 _22652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .Y(_956_)
);

AOI21X1 _22232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_458_),
    .B(_457_),
    .C(_249_),
    .Y(_496_)
);

AOI21X1 _13759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2895_),
    .B(_3118_),
    .C(_3117_),
    .Y(_3119_)
);

XNOR2X1 _13339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2654_),
    .Y(_2659_)
);

NAND2X1 _23857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2250_),
    .B(_2248_),
    .Y(_2266_)
);

FILL SFILL3720x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf4),
    .B(areg_30_bF$buf4),
    .Y(_1812_)
);

AOI22X1 _23017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf0),
    .B(areg_31_bF$buf2),
    .C(breg_20_bF$buf4),
    .D(areg_30_bF$buf4),
    .Y(_1354_)
);

FILL SFILL43960x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4144_),
    .B(_4134_),
    .C(_4139_),
    .Y(_4148_)
);

AOI21X1 _17592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7312_),
    .B(_7311_),
    .C(_7310_),
    .Y(_7318_)
);

OAI21X1 _17172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf0),
    .B(_5318_),
    .C(_6857_),
    .Y(_6858_)
);

FILL SFILL49160x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf2),
    .B(_2287__bF$buf0),
    .C(_5419_),
    .Y(_5469_)
);

NAND2X1 _18797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf3),
    .B(breg_17_bF$buf0),
    .Y(_8639_)
);

NAND3X1 _18377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8079_),
    .B(_8174_),
    .C(_8178_),
    .Y(_8179_)
);

NOR2X1 _13092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11767_),
    .B(_2388_),
    .Y(_2389_)
);

NOR3X1 _23190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1404_),
    .B(_1526_),
    .C(_1530_),
    .Y(_1542_)
);

NAND3X1 _21923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_142_),
    .B(_149_),
    .C(_129_),
    .Y(_158_)
);

INVX1 _21503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11605_),
    .Y(_11606_)
);

NAND3X1 _14297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3660_),
    .B(_3654_),
    .C(_3662_),
    .Y(_3708_)
);

FILL SFILL33880x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1016_),
    .B(_1010_),
    .C(_979_),
    .Y(_1017_)
);

NOR2X1 _16863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf2),
    .B(_3526_),
    .Y(_6519_)
);

NAND2X1 _16443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5690_),
    .B(_5700_),
    .Y(_6058_)
);

NAND3X1 _16023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5592_),
    .B(_5511_),
    .C(_5598_),
    .Y(_5599_)
);

FILL SFILL18600x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6985_),
    .B(_6987_),
    .C(_6978_),
    .Y(_7379_)
);

NAND2X1 _17228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6914_),
    .B(_6918_),
    .Y(_6919_)
);

OAI21X1 _12783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_10650_),
    .C(_10573_),
    .Y(_23_)
);

NOR2X1 _12363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf3),
    .B(_5420__bF$buf2),
    .Y(_7327_)
);

OAI21X1 _22881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_8773_),
    .C(_1045_),
    .Y(_1207_)
);

FILL SFILL23880x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf2),
    .B(breg_27_bF$buf1),
    .Y(_747_)
);

NOR3X1 _22041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_256_),
    .C(_278_),
    .Y(_287_)
);

FILL SFILL39080x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf1),
    .B(_10869__bF$buf3),
    .C(_3365_),
    .Y(_3369_)
);

NAND3X1 _13568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2854_),
    .B(_2852_),
    .C(_2848_),
    .Y(_2910_)
);

FILL SFILL23800x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2449_),
    .Y(_2450_)
);

AOI21X1 _23666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1999_),
    .B(_1922_),
    .C(_2043_),
    .Y(_2061_)
);

OAI21X1 _23246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1468_),
    .B(_1465_),
    .C(_1460_),
    .Y(_1604_)
);

FILL SFILL8840x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5235_),
    .B(_5241_),
    .C(_5243_),
    .Y(_5260_)
);

NOR2X1 _18186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7969_),
    .B(_7968_),
    .Y(_7970_)
);

FILL SFILL13800x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6564_),
    .B(_6570_),
    .C(_6548_),
    .Y(_6580_)
);

OAI21X1 _21732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11845_),
    .B(_11848_),
    .C(_11850_),
    .Y(_11857_)
);

OAI21X1 _21312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11388_),
    .B(_11389_),
    .C(_11386_),
    .Y(_11397_)
);

FILL SFILL29000x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_593_),
    .Y(_637_)
);

NAND3X1 _12419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7503_),
    .B(_7404_),
    .C(_7481_),
    .Y(_7942_)
);

INVX2 _22937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1266_),
    .Y(_1267_)
);

AOI21X1 _22517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_639_),
    .C(_807_),
    .Y(_808_)
);

INVX2 _16672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6309_),
    .Y(_6310_)
);

AND2X2 _16252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_18_bF$buf0),
    .Y(_5850_)
);

NAND3X1 _17877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7617_),
    .B(_7621_),
    .C(_7625_),
    .Y(_7631_)
);

NAND3X1 _17457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6923_),
    .B(_7004_),
    .C(_7008_),
    .Y(_7171_)
);

NAND3X1 _17037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_29_bF$buf5),
    .C(_6704_),
    .Y(_6710_)
);

AOI21X1 _12592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8435_),
    .B(_8446_),
    .C(_7054_),
    .Y(_9839_)
);

NAND3X1 _12172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5233_),
    .B(_5124_),
    .C(_5168_),
    .Y(_5244_)
);

NAND2X1 _22690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_996_),
    .B(_995_),
    .Y(_997_)
);

NAND3X1 _22270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_529_),
    .C(_525_),
    .Y(_537_)
);

FILL SFILL64360x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3147_),
    .B(_3144_),
    .Y(_3161_)
);

NOR3X1 _13377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2651_),
    .B(_2685_),
    .C(_2691_),
    .Y(_2701_)
);

BUFX2 _23895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[13]),
    .Y(y[13])
);

OAI21X1 _23475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1853_),
    .B(_1852_),
    .C(_1851_),
    .Y(_1854_)
);

NAND3X1 _23055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1394_),
    .B(_1395_),
    .C(_1393_),
    .Y(_1396_)
);

AND2X2 _19603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9131_),
    .B(_9125_),
    .Y(_9524_)
);

FILL SFILL54040x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5510_),
    .B(_5505_),
    .Y(_5511_)
);

OAI21X1 _15523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf2),
    .B(_2362__bF$buf5),
    .C(_5042_),
    .Y(_5050_)
);

NAND3X1 _15103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4590_),
    .B(_4589_),
    .C(_4587_),
    .Y(_4591_)
);

NAND3X1 _16728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6130_),
    .B(_6215_),
    .C(_6214_),
    .Y(_6371_)
);

NAND3X1 _16308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5909_),
    .B(_5910_),
    .C(_5908_),
    .Y(_5911_)
);

AOI21X1 _21961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_90_),
    .C(_11889_),
    .Y(_200_)
);

OAI21X1 _21541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11409_),
    .B(_11407_),
    .C(_11400_),
    .Y(_11647_)
);

NOR2X1 _21121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10865_),
    .B(_10912_),
    .Y(_11188_)
);

NAND2X1 _12648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_7_bF$buf1),
    .Y(_10452_)
);

OAI21X1 _12228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5837_),
    .B(_5826_),
    .C(_5815_),
    .Y(_5848_)
);

NOR2X1 _22746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1058_),
    .Y(_1059_)
);

AOI21X1 _22326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .B(_596_),
    .C(_594_),
    .Y(_599_)
);

AOI21X1 _16481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6081_),
    .B(_6085_),
    .C(_6089_),
    .Y(_6100_)
);

OAI21X1 _16061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5638_),
    .B(_5639_),
    .C(_5635_),
    .Y(_5641_)
);

OAI21X1 _17686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7420_),
    .B(_7016_),
    .C(_7051_),
    .Y(_7421_)
);

NAND2X1 _17266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_17_bF$buf0),
    .Y(_6961_)
);

FILL SFILL13800x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10843_),
    .B(_10848_),
    .Y(_10849_)
);

OAI21X1 _13186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2484_),
    .B(_2485_),
    .C(_2481_),
    .Y(_2492_)
);

AOI21X1 _23284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1520_),
    .C(_1529_),
    .Y(_1646_)
);

NOR2X1 _19832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9408_),
    .B(_9774_),
    .Y(_9775_)
);

OAI21X1 _19412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9310_),
    .B(_9309_),
    .C(_9308_),
    .Y(_9314_)
);

NAND2X1 _11919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf3),
    .B(areg_1_bF$buf3),
    .Y(_2464_)
);

DFFPOSX1 _24069_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[27]),
    .CLK(clk_bF$buf4),
    .D(b[27])
);

FILL SFILL64120x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4961_),
    .B(_5296_),
    .Y(_5301_)
);

NOR3X1 _15332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4836_),
    .B(_4838_),
    .C(_4835_),
    .Y(_4842_)
);

NAND3X1 _16957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6610_),
    .B(_6617_),
    .C(_6621_),
    .Y(_6622_)
);

NOR2X1 _16537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6156_),
    .B(_6160_),
    .Y(_6161_)
);

INVX1 _16117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5675_),
    .Y(_5701_)
);

INVX2 _21770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11896_),
    .Y(_11897_)
);

NAND2X1 _21350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11433_),
    .B(_11437_),
    .Y(_11438_)
);

INVX1 _12877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11668_),
    .Y(_1053_)
);

NAND2X1 _12457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8348_),
    .B(_8304_),
    .Y(_8359_)
);

NAND2X1 _22975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1307_),
    .B(_1303_),
    .Y(_1308_)
);

AOI21X1 _12037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3734_),
    .B(_3745_),
    .C(_3547_),
    .Y(_3756_)
);

NOR2X1 _22555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_849_),
    .B(_625_),
    .Y(_850_)
);

OAI21X1 _22135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_6300__bF$buf3),
    .C(_381_),
    .Y(_390_)
);

FILL SFILL54040x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_20_bF$buf2),
    .Y(_5891_)
);

OAI21X1 _14603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4031_),
    .B(_4035_),
    .C(_4037_),
    .Y(_4043_)
);

NAND3X1 _17495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6793_),
    .B(_7211_),
    .C(_7210_),
    .Y(_7212_)
);

AOI21X1 _17075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6262_),
    .B(_6355_),
    .C(_6751_),
    .Y(_6752_)
);

NOR2X1 _15808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5357_),
    .B(_5358_),
    .Y(_5362_)
);

AOI21X1 _20621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10637_),
    .B(_10638_),
    .C(_10345_),
    .Y(_10640_)
);

AOI21X1 _20201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10160_),
    .B(_10166_),
    .C(_10144_),
    .Y(_10179_)
);

FILL SFILL44040x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1322_),
    .B(_1320_),
    .C(_1316_),
    .Y(_1437_)
);

OAI21X1 _19641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9549_),
    .B(_9553_),
    .C(_9173_),
    .Y(_9566_)
);

OAI21X1 _19221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8719_),
    .B(_8703_),
    .C(_8711_),
    .Y(_9105_)
);

NAND3X1 _21826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_35_),
    .C(_39_),
    .Y(_51_)
);

AOI21X1 _21406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11498_),
    .B(_11499_),
    .C(_11497_),
    .Y(_11500_)
);

OAI21X1 _15981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5551_),
    .B(_5550_),
    .C(_5543_),
    .Y(_5553_)
);

AOI21X1 _15561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5086_),
    .B(_5087_),
    .C(_5085_),
    .Y(_5092_)
);

AOI21X1 _15141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4627_),
    .B(_4626_),
    .C(_4349_),
    .Y(_4633_)
);

FILL SFILL23400x50 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6409_),
    .B(_6410_),
    .C(_6043_),
    .Y(_6413_)
);

FILL SFILL74120x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5950_),
    .B(_5952_),
    .C(_5951_),
    .Y(_5953_)
);

INVX8 _12686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf0),
    .Y(_10869_)
);

INVX1 _12266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6198_),
    .Y(_6264_)
);

INVX2 _22784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1099_),
    .Y(_1100_)
);

NOR2X1 _22364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_640_),
    .B(_634_),
    .Y(_641_)
);

OAI21X1 _18912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8333_),
    .B(_8765_),
    .C(_8342_),
    .Y(_8766_)
);

FILL SFILL59160x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23989_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[43]),
    .CLK(clk_bF$buf7),
    .D(_0_[43])
);

OAI21X1 _23569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1952_),
    .B(_1953_),
    .C(_1954_),
    .Y(_1955_)
);

FILL SFILL64120x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _23149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf2),
    .B(areg_30_bF$buf1),
    .C(breg_22_bF$buf4),
    .D(areg_29_bF$buf2),
    .Y(_1498_)
);

NAND3X1 _14832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4291_),
    .B(_4293_),
    .C(_4290_),
    .Y(_4294_)
);

INVX2 _14412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3809_),
    .Y(_3834_)
);

NAND2X1 _15617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_17_bF$buf5),
    .Y(_5153_)
);

OR2X2 _20850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10843_),
    .B(_10848_),
    .Y(_10890_)
);

NAND3X1 _20430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10393_),
    .B(_10428_),
    .C(_10424_),
    .Y(_10429_)
);

NAND3X1 _20010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9967_),
    .B(_9968_),
    .C(_9966_),
    .Y(_9969_)
);

OAI21X1 _18089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7842_),
    .B(_7847_),
    .C(_7849_),
    .Y(_7863_)
);

FILL SFILL49160x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _19870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9430_),
    .Y(_9816_)
);

INVX2 _19450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9320_),
    .Y(_9355_)
);

OAI21X1 _19030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8503_),
    .B(_8488_),
    .C(_8513_),
    .Y(_8894_)
);

FILL SFILL54120x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _11957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2749_),
    .B(_2869_),
    .Y(_2880_)
);

AOI21X1 _21635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11749_),
    .B(_11748_),
    .C(_11747_),
    .Y(_11750_)
);

NOR3X1 _21215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10964_),
    .B(_10971_),
    .C(_10974_),
    .Y(_11291_)
);

OAI21X1 _15790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5339_),
    .B(_5340_),
    .C(_5341_),
    .Y(_5342_)
);

OAI21X1 _15370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4882_),
    .B(_4881_),
    .C(_4880_),
    .Y(_4883_)
);

NAND3X1 _16995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6662_),
    .B(_6663_),
    .C(_6661_),
    .Y(_6664_)
);

NAND3X1 _16575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6193_),
    .B(_6186_),
    .C(_6191_),
    .Y(_6203_)
);

NAND2X1 _16155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5737_),
    .B(_5742_),
    .Y(_5743_)
);

FILL SFILL54200x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44040x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf4),
    .B(breg_6_bF$buf3),
    .C(areg_4_bF$buf1),
    .D(breg_7_bF$buf1),
    .Y(_8775_)
);

NAND3X1 _12075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg_5_bF$buf0),
    .C(_3536_),
    .Y(_4171_)
);

AOI21X1 _22593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_891_),
    .B(_887_),
    .C(_730_),
    .Y(_892_)
);

OAI21X1 _22173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_430_),
    .C(_428_),
    .Y(_432_)
);

OAI21X1 _18721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8547_),
    .B(_8546_),
    .C(_8543_),
    .Y(_8556_)
);

NOR2X1 _18301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7680_),
    .B(_8094_),
    .Y(_8096_)
);

NOR2X1 _20906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10951_),
    .B(_10909_),
    .Y(_10952_)
);

OAI21X1 _23798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2155_),
    .C(_2203_),
    .Y(_2204_)
);

NOR2X1 _23378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1623_),
    .B(_1624_),
    .Y(_1748_)
);

OAI21X1 _19926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf3),
    .B(_7100__bF$buf2),
    .C(_9866_),
    .Y(_9878_)
);

OAI21X1 _19506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9415_),
    .B(_9416_),
    .C(_9414_),
    .Y(_9417_)
);

FILL SFILL69240x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _14641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4078_),
    .B(_4079_),
    .Y(_4084_)
);

AOI21X1 _14221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3623_),
    .B(_3622_),
    .C(_3621_),
    .Y(_3625_)
);

FILL SFILL34040x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5403_),
    .B(_5399_),
    .Y(_5404_)
);

NOR3X1 _15426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4941_),
    .B(_4942_),
    .C(_4940_),
    .Y(_4945_)
);

AOI21X1 _15006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4475_),
    .B(_4482_),
    .C(_4483_),
    .Y(_4484_)
);

NAND2X1 _21864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_92_),
    .Y(_93_)
);

FILL SFILL59240x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11521_),
    .B(_11520_),
    .C(_11519_),
    .Y(_11542_)
);

AOI21X1 _21024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10817_),
    .B(_11080_),
    .C(_11079_),
    .Y(_11081_)
);

FILL SFILL23800x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf1),
    .B(_7225__bF$buf0),
    .Y(_952_)
);

OAI21X1 _22229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_491_),
    .B(_244_),
    .C(_474_),
    .Y(_492_)
);

INVX1 _13912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3259_),
    .Y(_3287_)
);

NAND3X1 _16384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5975_),
    .B(_5981_),
    .C(_5984_),
    .Y(_5994_)
);

FILL SFILL28760x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74120x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28680x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7309_),
    .B(_7313_),
    .C(_7273_),
    .Y(_7314_)
);

AND2X2 _17169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg_24_bF$buf4),
    .Y(_6854_)
);

FILL FILL74040x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8757_),
    .B(_8758_),
    .C(_8755_),
    .Y(_8807_)
);

OAI22X1 _18530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7518_),
    .B(_8346_),
    .C(_7962_),
    .D(_7958_),
    .Y(_8347_)
);

XNOR2X1 _18110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7885_),
    .B(_7883_),
    .Y(_7886_)
);

FILL SFILL54120x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10410_),
    .B(_10417_),
    .Y(_10742_)
);

NAND3X1 _13089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg_14_bF$buf2),
    .C(_2384_),
    .Y(_2385_)
);

AOI21X1 _23187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1255_),
    .B(_1094_),
    .C(_1538_),
    .Y(_1539_)
);

OAI21X1 _19735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf3),
    .B(_5668__bF$buf4),
    .C(_9655_),
    .Y(_9668_)
);

NAND2X1 _19315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9207_),
    .B(_9206_),
    .Y(_9208_)
);

NAND3X1 _14870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4047_),
    .B(_4334_),
    .C(_4331_),
    .Y(_4335_)
);

NAND2X1 _14450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_11_bF$buf3),
    .Y(_3875_)
);

AOI21X1 _14030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3413_),
    .B(_3414_),
    .C(_3397_),
    .Y(_3415_)
);

FILL SFILL59000x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33640x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39160x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf0),
    .B(areg_23_bF$buf3),
    .Y(_5195_)
);

INVX2 _15235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4711_),
    .Y(_4735_)
);

NOR2X1 _11995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3274_),
    .B(_3285_),
    .Y(_3296_)
);

FILL SFILL54120x50 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11779_),
    .B(_11770_),
    .C(_11755_),
    .Y(_11792_)
);

INVX2 _21253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11331_),
    .Y(_11332_)
);

NAND2X1 _17801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7526_),
    .B(_7522_),
    .Y(_7548_)
);

NOR2X1 _22878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3526_),
    .B(_9153_),
    .Y(_1203_)
);

OAI21X1 _22458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_512_),
    .B(_742_),
    .C(_741_),
    .Y(_743_)
);

AOI21X1 _22038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_279_),
    .C(_254_),
    .Y(_283_)
);

FILL SFILL69240x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3058_),
    .B(_3070_),
    .C(_3076_),
    .Y(_3078_)
);

AOI21X1 _13301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2425_),
    .B(_2440_),
    .C(_2615_),
    .Y(_2618_)
);

INVX1 _16193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5783_),
    .Y(_5784_)
);

NAND2X1 _14926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4394_),
    .B(_4395_),
    .Y(_4396_)
);

INVX1 _14506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3674_),
    .Y(_3937_)
);

AND2X2 _17398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7102_),
    .B(_7105_),
    .Y(_7106_)
);

FILL SFILL69160x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8520x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10340_),
    .B(_10652_),
    .C(_10689_),
    .Y(_10994_)
);

AOI21X1 _20524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10514_),
    .B(_10521_),
    .C(_10499_),
    .Y(_10533_)
);

NAND3X1 _20104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10065_),
    .B(_10070_),
    .C(_10071_),
    .Y(_10072_)
);

NAND3X1 _19964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9898_),
    .B(_9856_),
    .C(_9899_),
    .Y(_9919_)
);

NOR3X1 _19544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9445_),
    .B(_9441_),
    .C(_9443_),
    .Y(_9459_)
);

AND2X2 _19124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8581_),
    .B(_8572_),
    .Y(_8998_)
);

NAND3X1 _21729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11850_),
    .B(_11851_),
    .C(_11852_),
    .Y(_11853_)
);

NAND3X1 _21309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11371_),
    .B(_11387_),
    .C(_11392_),
    .Y(_11393_)
);

FILL FILL74200x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .B(_5441_),
    .C(_5405_),
    .Y(_5446_)
);

AND2X2 _15464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4984_),
    .B(_4982_),
    .Y(_4985_)
);

NAND2X1 _15044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4521_),
    .B(_4525_),
    .Y(_4526_)
);

FILL FILL74120x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6302_),
    .B(_6305_),
    .Y(_6306_)
);

OAI21X1 _16249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5483_),
    .B(_5473_),
    .C(_5477_),
    .Y(_5846_)
);

OAI21X1 _21482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11579_),
    .B(_11583_),
    .C(_11317_),
    .Y(_11584_)
);

AOI21X1 _21062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10815_),
    .B(_10903_),
    .C(_11122_),
    .Y(_11123_)
);

FILL SFILL18760x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL14040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7325_),
    .B(_7321_),
    .C(_7333_),
    .Y(_7337_)
);

FILL SFILL33960x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38520x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8238_),
    .B(_9729_),
    .C(_9740_),
    .Y(_9806_)
);

OAI21X1 _12169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_5190__bF$buf0),
    .C(_4423_),
    .Y(_5201_)
);

XNOR2X1 _22687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_993_),
    .B(_992_),
    .Y(_994_)
);

NOR3X1 _22267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .B(_532_),
    .C(_533_),
    .Y(_534_)
);

OAI22X1 _18815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7884_),
    .B(_8657_),
    .C(_8658_),
    .D(_8284_),
    .Y(_8659_)
);

OAI21X1 _13950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf5),
    .B(_7711__bF$buf1),
    .C(_3071_),
    .Y(_3328_)
);

NAND2X1 _13530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2862_),
    .B(_2867_),
    .Y(_2868_)
);

OAI21X1 _13110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2407_),
    .B(_2088_),
    .C(_2001_),
    .Y(_2408_)
);

FILL SFILL39160x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4185_),
    .B(_4186_),
    .C(_4184_),
    .Y(_4187_)
);

NOR3X1 _14315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3720_),
    .B(_3727_),
    .C(_3592_),
    .Y(_3728_)
);

FILL SFILL23960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10766_),
    .B(_10771_),
    .C(_10773_),
    .Y(_10784_)
);

AOI21X1 _20333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9967_),
    .B(_9968_),
    .C(_9639_),
    .Y(_10324_)
);

OAI21X1 _19773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9706_),
    .B(_9705_),
    .C(_9709_),
    .Y(_9710_)
);

NOR3X1 _19353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8854_),
    .B(_8857_),
    .C(_8860_),
    .Y(_9250_)
);

AOI21X1 _21958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_194_),
    .C(_193_),
    .Y(_196_)
);

NAND3X1 _21538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11607_),
    .B(_11635_),
    .C(_11632_),
    .Y(_11644_)
);

NAND3X1 _21118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11177_),
    .B(_11180_),
    .C(_11183_),
    .Y(_11184_)
);

NAND2X1 _12801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_9_bF$buf1),
    .Y(_221_)
);

NAND3X1 _15693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5104_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5236_)
);

INVX2 _15273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4776_),
    .Y(_4777_)
);

OAI21X1 _16898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf0),
    .B(_2560__bF$buf1),
    .C(_6553_),
    .Y(_6557_)
);

NAND3X1 _16478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6058_),
    .B(_6095_),
    .C(_6090_),
    .Y(_6096_)
);

NAND3X1 _16058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5620_),
    .C(_5622_),
    .Y(_5637_)
);

NAND2X1 _21291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf0),
    .B(breg_25_bF$buf2),
    .Y(_11374_)
);

CLKBUF1 CLKBUF1_insert90 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert91 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert92 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert93 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert94 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

FILL SFILL43640x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _12398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .Y(_7711_)
);

NAND3X1 _22496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_782_),
    .C(_784_),
    .Y(_785_)
);

AOI21X1 _22076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_117_),
    .B(_118_),
    .C(_103_),
    .Y(_325_)
);

NAND3X1 _18624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8075_),
    .B(_8444_),
    .C(_8445_),
    .Y(_8450_)
);

AOI21X1 _18204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7988_),
    .B(_7989_),
    .C(_7987_),
    .Y(_7990_)
);

NAND3X1 _20809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10837_),
    .B(_10821_),
    .C(_10841_),
    .Y(_10845_)
);

FILL FILL74200x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf0),
    .B(_3402__bF$buf1),
    .C(_9408_),
    .Y(_9771_)
);

NOR3X1 _19409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9297_),
    .B(_9283_),
    .C(_9302_),
    .Y(_9310_)
);

OAI21X1 _14964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4436_),
    .B(_4435_),
    .C(_4437_),
    .Y(_4438_)
);

XOR2X1 _14544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3954_),
    .B(_3949_),
    .Y(_3979_)
);

AOI21X1 _14124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3458_),
    .B(_3465_),
    .C(_3248_),
    .Y(_3518_)
);

NAND2X1 _15749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4957_),
    .B(_5292_),
    .Y(_5297_)
);

AOI22X1 _15329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4530_),
    .B(_4531_),
    .C(_4837_),
    .D(_4529_),
    .Y(_4838_)
);

AOI21X1 _20982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11029_),
    .B(_11033_),
    .C(_11021_),
    .Y(_11034_)
);

AOI21X1 _20562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10217_),
    .B(_10223_),
    .C(_10226_),
    .Y(_10575_)
);

NAND2X1 _20142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf2),
    .B(breg_21_bF$buf4),
    .Y(_10114_)
);

OAI21X1 _19582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9500_),
    .B(_9498_),
    .C(_9490_),
    .Y(_9501_)
);

OAI21X1 _19162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8671_),
    .B(_8638_),
    .C(_8663_),
    .Y(_9040_)
);

FILL SFILL33960x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _21767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11893_),
    .Y(_11894_)
);

NAND3X1 _21347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11423_),
    .B(_11419_),
    .C(_11431_),
    .Y(_11435_)
);

NAND2X1 _12610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_12_bF$buf3),
    .Y(_10035_)
);

AOI21X1 _15082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4557_),
    .B(_4549_),
    .C(_4535_),
    .Y(_4568_)
);

AOI21X1 _13815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3180_),
    .B(_3179_),
    .C(_3126_),
    .Y(_3181_)
);

BUFX2 _23913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[31]),
    .Y(y[31])
);

OAI21X1 _16287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5514_),
    .B(_5887_),
    .C(_5522_),
    .Y(_5888_)
);

XNOR2X1 _18853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8700_),
    .B(_8697_),
    .Y(_8701_)
);

AOI21X1 _18433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8233_),
    .B(_8234_),
    .C(_8226_),
    .Y(_8241_)
);

NAND2X1 _18013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7774_),
    .B(_7779_),
    .Y(_7780_)
);

AOI21X1 _20618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10630_),
    .B(_10635_),
    .C(_10346_),
    .Y(_10636_)
);

OAI21X1 _19638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9555_),
    .B(_9561_),
    .C(_9183_),
    .Y(_9562_)
);

NAND2X1 _19218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf1),
    .B(areg_23_bF$buf1),
    .Y(_9100_)
);

NAND3X1 _14773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4222_),
    .B(_4228_),
    .C(_4206_),
    .Y(_4229_)
);

OAI21X1 _14353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3768_),
    .B(_3767_),
    .C(_3494_),
    .Y(_3769_)
);

FILL SFILL13960x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24031_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[21]),
    .CLK(clk_bF$buf4),
    .D(a[21])
);

NAND3X1 _15978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .B(_5548_),
    .C(_5547_),
    .Y(_5549_)
);

NAND3X1 _15558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5086_),
    .B(_5087_),
    .C(_5085_),
    .Y(_5088_)
);

NAND3X1 _15138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4625_),
    .B(_4628_),
    .C(_4348_),
    .Y(_4629_)
);

AND2X2 _20791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf2),
    .B(areg_21_bF$buf0),
    .Y(_10826_)
);

NAND2X1 _20371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_10365_)
);

OAI21X1 _19391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf1),
    .B(_5668__bF$buf4),
    .C(_8907_),
    .Y(_9291_)
);

OR2X2 _21996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_236_),
    .B(_230_),
    .Y(_237_)
);

NAND3X1 _21576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11648_),
    .B(_11678_),
    .C(_11684_),
    .Y(_11685_)
);

NAND2X1 _21156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf0),
    .B(areg_27_bF$buf0),
    .Y(_11226_)
);

XOR2X1 _17704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7392_),
    .B(_7440_),
    .Y(_7441_)
);

OAI21X1 _18909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8757_),
    .B(_8758_),
    .C(_8761_),
    .Y(_8762_)
);

AOI22X1 _13624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .B(_2971_),
    .C(_2963_),
    .D(_2958_),
    .Y(_2972_)
);

OAI21X1 _13204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2511_),
    .C(_2509_),
    .Y(_2512_)
);

AOI21X1 _23722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2058_),
    .B(_2098_),
    .C(_2121_),
    .Y(_2122_)
);

NOR2X1 _23302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf2),
    .B(_7225__bF$buf2),
    .Y(_1665_)
);

AND2X2 _16096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf0),
    .B(breg_25_bF$buf3),
    .Y(_5678_)
);

NAND2X1 _14829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4288_),
    .B(_4289_),
    .Y(_4290_)
);

AOI21X1 _14409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3815_),
    .B(_3814_),
    .C(_3811_),
    .Y(_3830_)
);

NAND2X1 _18662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_29_bF$buf3),
    .Y(_8491_)
);

OAI21X1 _18242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8012_),
    .B(_8018_),
    .C(_8021_),
    .Y(_8031_)
);

AOI21X1 _20847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10868_),
    .B(_10875_),
    .C(_10852_),
    .Y(_10887_)
);

AOI21X1 _20427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10410_),
    .B(_10416_),
    .C(_10394_),
    .Y(_10426_)
);

AOI21X1 _20007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9273_),
    .B(_9607_),
    .C(_9614_),
    .Y(_9966_)
);

OAI22X1 _19867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9100_),
    .B(_9811_),
    .C(_9812_),
    .D(_9484_),
    .Y(_9813_)
);

AOI21X1 _19447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9032_),
    .B(_9013_),
    .C(_9035_),
    .Y(_9352_)
);

NAND2X1 _19027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8572_),
    .B(_8581_),
    .Y(_8891_)
);

NAND2X1 _14582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4020_),
    .B(_4018_),
    .Y(_4021_)
);

NAND3X1 _14162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3539_),
    .B(_3553_),
    .C(_3559_),
    .Y(_3560_)
);

FILL SFILL8680x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5334_),
    .B(_5335_),
    .C(_5333_),
    .Y(_5339_)
);

AOI21X1 _15367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4535_),
    .B(_4557_),
    .C(_4879_),
    .Y(_4880_)
);

NAND3X1 _20180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10146_),
    .B(_10153_),
    .C(_10154_),
    .Y(_10155_)
);

FILL SFILL8600x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11476_),
    .Y(_11477_)
);

OAI21X1 _17933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7691_),
    .B(_7684_),
    .C(_7670_),
    .Y(_7692_)
);

OAI21X1 _17513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6837_),
    .B(_6817_),
    .C(_7230_),
    .Y(_7231_)
);

FILL SFILL74280x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8529_),
    .B(_8545_),
    .C(_8551_),
    .Y(_8552_)
);

OAI21X1 _13853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3218_),
    .B(_3222_),
    .C(_2983_),
    .Y(_3223_)
);

OAI21X1 _13433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2580_),
    .C(_2612_),
    .Y(_2762_)
);

DFFPOSX1 _23951_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[5]),
    .CLK(clk_bF$buf7),
    .D(_0_[5])
);

NAND3X1 _13013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .B(_2292_),
    .C(_2289_),
    .Y(_2308_)
);

AOI21X1 _23531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .B(_1893_),
    .C(_1912_),
    .Y(_1915_)
);

NAND2X1 _23111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1355_),
    .B(_1351_),
    .Y(_1457_)
);

FILL SFILL74200x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4078_),
    .B(_4079_),
    .Y(_4080_)
);

XNOR2X1 _14218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3597_),
    .B(_3620_),
    .Y(_3621_)
);

AND2X2 _18891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_27_bF$buf2),
    .Y(_8743_)
);

NAND2X1 _18471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7911_),
    .B(_7916_),
    .Y(_8283_)
);

INVX1 _18051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7820_),
    .Y(_7822_)
);

FILL SFILL64280x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _20656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10649_),
    .B(_10339_),
    .C(_10653_),
    .Y(_10677_)
);

NAND2X1 _20236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_11_bF$buf1),
    .B(areg_27_bF$buf3),
    .Y(_10216_)
);

NAND3X1 _19676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9602_),
    .B(_9603_),
    .C(_9601_),
    .Y(_9604_)
);

AOI21X1 _19256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8339_),
    .B(_9142_),
    .C(_8757_),
    .Y(_9143_)
);

FILL SFILL64200x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf0),
    .B(_2763_),
    .Y(_3811_)
);

FILL SFILL33720x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9225_),
    .B(_9027_),
    .C(_9257_),
    .Y(_11066_)
);

OR2X2 _22802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_959_),
    .B(_1119_),
    .Y(_1120_)
);

INVX2 _15596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5105_),
    .Y(_5130_)
);

INVX1 _15176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4669_),
    .Y(_4670_)
);

AOI21X1 _13909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3269_),
    .B(_3265_),
    .C(_3272_),
    .Y(_3283_)
);

NAND3X1 _21194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11015_),
    .B(_11128_),
    .C(_11127_),
    .Y(_11268_)
);

NAND2X1 _17742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7477_),
    .B(_7482_),
    .Y(_7483_)
);

NOR2X1 _17322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7019_),
    .B(_7021_),
    .Y(_7022_)
);

FILL SFILL74120x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _22399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_677_),
    .B(_676_),
    .Y(_678_)
);

AOI21X1 _18947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8406_),
    .B(_8404_),
    .C(_8803_),
    .Y(_8804_)
);

OAI21X1 _18527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_7100__bF$buf3),
    .C(_8338_),
    .Y(_8344_)
);

INVX2 _18107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7882_),
    .Y(_7883_)
);

INVX1 _13662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2764_),
    .Y(_3013_)
);

NAND2X1 _13242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2370_),
    .B(_2372_),
    .Y(_2553_)
);

NOR2X1 _23760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2151_),
    .Y(_2162_)
);

OR2X2 _23340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .B(_1704_),
    .Y(_1706_)
);

NAND3X1 _14867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4057_),
    .B(_4326_),
    .C(_4321_),
    .Y(_4332_)
);

XOR2X1 _14447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3870_),
    .B(_3871_),
    .Y(_3872_)
);

AOI21X1 _14027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3150_),
    .B(_3153_),
    .C(_3160_),
    .Y(_3412_)
);

FILL SFILL8600x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8071_),
    .Y(_8072_)
);

FILL SFILL13640x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10923_),
    .B(_10925_),
    .C(_10917_),
    .Y(_10929_)
);

XNOR2X1 _20465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10467_),
    .B(_10465_),
    .Y(_10468_)
);

NAND2X1 _20045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf4),
    .B(breg_29_bF$buf0),
    .Y(_10007_)
);

NAND2X1 _19485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf0),
    .B(breg_21_bF$buf4),
    .Y(_9394_)
);

AND2X2 _19065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8929_),
    .B(_8932_),
    .Y(_8933_)
);

XNOR2X1 _12933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(_1653_),
    .Y(_1663_)
);

INVX2 _12513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8961_),
    .Y(_8972_)
);

NAND3X1 _22611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_905_),
    .C(_906_),
    .Y(_912_)
);

FILL SFILL38840x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3068_),
    .B(_3073_),
    .Y(_3074_)
);

NOR2X1 _23816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8759_),
    .B(_6815__bF$buf1),
    .Y(_2223_)
);

BUFX2 BUFX2_insert300 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .Y(_2825__bF$buf4)
);

BUFX2 BUFX2_insert301 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .Y(_2825__bF$buf3)
);

BUFX2 BUFX2_insert302 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .Y(_2825__bF$buf2)
);

BUFX2 BUFX2_insert303 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .Y(_2825__bF$buf1)
);

BUFX2 BUFX2_insert304 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825_),
    .Y(_2825__bF$buf0)
);

OAI21X1 _17971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7726_),
    .B(_7725_),
    .C(_7723_),
    .Y(_7734_)
);

BUFX2 BUFX2_insert305 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf5)
);

OAI21X1 _17551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6890_),
    .B(_7271_),
    .C(_6882_),
    .Y(_7273_)
);

BUFX2 BUFX2_insert306 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf4)
);

OAI21X1 _17131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6774_),
    .B(_6776_),
    .C(_6764_),
    .Y(_6813_)
);

BUFX2 BUFX2_insert307 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf3)
);

BUFX2 BUFX2_insert308 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf2)
);

BUFX2 BUFX2_insert309 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[18]),
    .Y(breg_18_bF$buf1)
);

AND2X2 _18756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8167_),
    .B(_8162_),
    .Y(_8594_)
);

OAI21X1 _18336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf1),
    .B(_5315__bF$buf3),
    .C(_8126_),
    .Y(_8134_)
);

XOR2X1 _13891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2996_),
    .B(_3262_),
    .Y(_3264_)
);

AOI21X1 _13471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .B(_2597_),
    .C(_2802_),
    .Y(_2804_)
);

NAND3X1 _13051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1096_),
    .B(_1140_),
    .C(_1162_),
    .Y(_2346_)
);

FILL SFILL54200x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4099_),
    .Y(_4122_)
);

FILL SFILL13800x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _14256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3656_),
    .B(_3659_),
    .C(_3655_),
    .Y(_3663_)
);

FILL SFILL13720x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10358_),
    .B(_10362_),
    .C(_10366_),
    .Y(_10719_)
);

AOI22X1 _20274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf4),
    .B(areg_31_bF$buf3),
    .C(breg[8]),
    .D(areg_30_bF$buf2),
    .Y(_10259_)
);

NAND3X1 _16822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6466_),
    .B(_6470_),
    .C(_6473_),
    .Y(_6474_)
);

AOI21X1 _16402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5996_),
    .B(_6002_),
    .C(_5743_),
    .Y(_6014_)
);

OAI21X1 _19294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8816_),
    .B(_8783_),
    .C(_9184_),
    .Y(_9185_)
);

NAND2X1 _21899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf0),
    .B(areg_29_bF$buf1),
    .Y(_131_)
);

NAND3X1 _21479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11322_),
    .B(_11574_),
    .C(_11577_),
    .Y(_11580_)
);

AOI21X1 _21059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11113_),
    .B(_11114_),
    .C(_11112_),
    .Y(_11119_)
);

OAI21X1 _17607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7331_),
    .B(_7330_),
    .C(_7333_),
    .Y(_7334_)
);

OAI21X1 _12742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11472_),
    .B(_11461_),
    .C(_11450_),
    .Y(_11483_)
);

AOI21X1 _12322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6856_),
    .B(_6867_),
    .C(_6791_),
    .Y(_6878_)
);

INVX2 _22840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .Y(_1161_)
);

NOR3X1 _22420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_464_),
    .C(_468_),
    .Y(_702_)
);

FILL SFILL69480x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_11882_),
    .C(_226_),
    .Y(_241_)
);

AND2X2 _13947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf1),
    .B(breg_10_bF$buf5),
    .Y(_3325_)
);

NOR3X1 _13527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2859_),
    .B(_2854_),
    .C(_2860_),
    .Y(_2865_)
);

NAND2X1 _13107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2396_),
    .Y(_2405_)
);

XNOR2X1 _23625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2016_),
    .B(_2011_),
    .Y(_2017_)
);

NAND2X1 _23205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1558_),
    .Y(_1559_)
);

AND2X2 _17780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7517_),
    .B(_7518_),
    .Y(_7524_)
);

OAI21X1 _17360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6731_),
    .B(_7063_),
    .C(_6721_),
    .Y(_7064_)
);

AOI21X1 _18985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8843_),
    .B(_8844_),
    .C(_8842_),
    .Y(_8845_)
);

NAND3X1 _18565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8355_),
    .B(_8349_),
    .C(_8353_),
    .Y(_8385_)
);

OAI21X1 _18145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7924_),
    .B(_7923_),
    .C(_7922_),
    .Y(_7925_)
);

INVX2 _13280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .Y(_2594_)
);

FILL SFILL38920x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL38840x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3705_),
    .B(_3704_),
    .C(_3669_),
    .Y(_3914_)
);

NAND3X1 _14065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3430_),
    .B(_3436_),
    .C(_3434_),
    .Y(_3454_)
);

FILL SFILL3560x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3480x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10047_),
    .B(_10048_),
    .Y(_10049_)
);

OAI21X1 _16631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5964_),
    .B(_6263_),
    .C(_5954_),
    .Y(_6265_)
);

NAND3X1 _16211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5782_),
    .B(_5798_),
    .C(_5803_),
    .Y(_5805_)
);

FILL SFILL28840x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11075_),
    .B(_11083_),
    .Y(_11370_)
);

AOI21X1 _17836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7581_),
    .B(_7579_),
    .C(_7578_),
    .Y(_7586_)
);

AOI21X1 _17416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7123_),
    .B(_7125_),
    .C(_7108_),
    .Y(_7126_)
);

NAND3X1 _12971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2066_),
    .B(_1914_),
    .C(_2001_),
    .Y(_2077_)
);

OAI21X1 _12551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9334_),
    .B(_9345_),
    .C(_9301_),
    .Y(_9389_)
);

OAI21X1 _12131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4774_),
    .B(_4763_),
    .C(_4730_),
    .Y(_4785_)
);

AOI21X1 _13756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3105_),
    .B(_3104_),
    .C(_3101_),
    .Y(_3116_)
);

NOR2X1 _13336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .B(_2655_),
    .Y(_2656_)
);

NAND2X1 _23854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2252_),
    .B(_2245_),
    .Y(_2263_)
);

NOR2X1 _23434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1733_),
    .Y(_1809_)
);

OAI21X1 _23014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1204_),
    .C(_1208_),
    .Y(_1351_)
);

FILL SFILL18840x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf3),
    .B(breg_14_bF$buf0),
    .Y(_5466_)
);

OAI21X1 _18794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8258_),
    .B(_8225_),
    .C(_8251_),
    .Y(_8636_)
);

AOI21X1 _18374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8162_),
    .B(_8166_),
    .C(_8121_),
    .Y(_8176_)
);

NOR2X1 _20979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10713_),
    .B(_11030_),
    .Y(_11031_)
);

NOR2X1 _20559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10222_),
    .B(_10570_),
    .Y(_10571_)
);

NAND2X1 _20139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9836_),
    .B(_9843_),
    .Y(_10110_)
);

OAI21X1 _21920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_150_),
    .C(_127_),
    .Y(_154_)
);

OAI21X1 _21500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11438_),
    .B(_11563_),
    .C(_11555_),
    .Y(_11602_)
);

NAND3X1 _19999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9952_),
    .B(_9951_),
    .C(_9950_),
    .Y(_9957_)
);

NAND2X1 _19579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf5),
    .B(areg_27_bF$buf2),
    .Y(_9497_)
);

AOI21X1 _19159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9022_),
    .B(_9026_),
    .C(_9014_),
    .Y(_9036_)
);

NAND3X1 _14294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3694_),
    .B(_3689_),
    .C(_3676_),
    .Y(_3705_)
);

FILL SFILL69080x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8687_),
    .B(_9991_),
    .Y(_10002_)
);

AOI21X1 _22705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1013_),
    .B(_1012_),
    .C(_1005_),
    .Y(_1014_)
);

AND2X2 _15499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4694_),
    .B(_5021_),
    .Y(_5023_)
);

NOR3X1 _15079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4255_),
    .B(_4254_),
    .C(_4256_),
    .Y(_4564_)
);

XOR2X1 _16860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6455_),
    .B(_6514_),
    .Y(_6515_)
);

INVX1 _16440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6053_),
    .Y(_6054_)
);

AOI21X1 _16020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5590_),
    .B(_5589_),
    .C(_5588_),
    .Y(_5595_)
);

INVX2 _21097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11134_),
    .Y(_11161_)
);

OAI21X1 _17645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7361_),
    .B(_7365_),
    .C(_7367_),
    .Y(_7376_)
);

NAND3X1 _17225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6902_),
    .B(_6912_),
    .C(_6906_),
    .Y(_6916_)
);

NAND2X1 _12780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11822_),
    .B(_11800_),
    .Y(_11898_)
);

OAI21X1 _12360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6812_),
    .B(_6791_),
    .C(_6703_),
    .Y(_7294_)
);

FILL SFILL38920x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3364_),
    .B(_3365_),
    .Y(_3366_)
);

AOI21X1 _13565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2893_),
    .B(_2890_),
    .C(_2875_),
    .Y(_2907_)
);

NAND2X1 _13145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2441_),
    .B(_2446_),
    .Y(_2447_)
);

NAND2X1 _23663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .B(_2057_),
    .Y(_2058_)
);

OAI21X1 _23243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1600_),
    .B(_1599_),
    .C(_1597_),
    .Y(_1601_)
);

DFFPOSX1 _24028_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[18]),
    .CLK(clk_bF$buf5),
    .D(a[18])
);

FILL SFILL28920x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5249_),
    .B(_5008_),
    .C(_5255_),
    .Y(_5257_)
);

NAND2X1 _18183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_2_bF$buf4),
    .B(areg_31_bF$buf1),
    .Y(_7967_)
);

NAND2X1 _20788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf1),
    .B(breg_20_bF$buf2),
    .Y(_10822_)
);

NAND2X1 _20368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10359_),
    .B(_10360_),
    .Y(_10361_)
);

NAND3X1 _16916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6572_),
    .B(_6546_),
    .C(_6576_),
    .Y(_6577_)
);

AND2X2 _19388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_8_bF$buf2),
    .B(breg_28_bF$buf2),
    .Y(_9287_)
);

FILL SFILL18520x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_9104__bF$buf1),
    .C(_593_),
    .Y(_604_)
);

AOI21X1 _12416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7810_),
    .B(_7777_),
    .C(_7635_),
    .Y(_7909_)
);

INVX1 _22934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .Y(_1264_)
);

AOI21X1 _22514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_803_),
    .B(_804_),
    .C(_796_),
    .Y(_805_)
);

NAND2X1 _23719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .B(_2105_),
    .Y(_2118_)
);

OAI21X1 _17874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7626_),
    .B(_7627_),
    .C(_7625_),
    .Y(_7628_)
);

AOI21X1 _17454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7149_),
    .B(_7155_),
    .C(_7062_),
    .Y(_7168_)
);

OAI21X1 _17034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6706_),
    .B(_6700_),
    .C(_6695_),
    .Y(_6707_)
);

FILL SFILL53960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf3),
    .B(_6815__bF$buf1),
    .Y(_8487_)
);

NAND3X1 _18239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7664_),
    .B(_7776_),
    .C(_7778_),
    .Y(_8027_)
);

NAND3X1 _13794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3150_),
    .B(_3153_),
    .C(_3151_),
    .Y(_3158_)
);

NAND3X1 _13374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2626_),
    .B(_2692_),
    .C(_2697_),
    .Y(_2698_)
);

BUFX2 _23892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[10]),
    .Y(y[10])
);

AOI21X1 _23472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1623_),
    .B(_1742_),
    .C(_1750_),
    .Y(_1851_)
);

AOI21X1 _23052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1099_),
    .B(_1242_),
    .C(_1248_),
    .Y(_1393_)
);

AOI21X1 _19600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9168_),
    .B(_9171_),
    .C(_9178_),
    .Y(_9520_)
);

NAND3X1 _14999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4468_),
    .B(_4474_),
    .C(_4453_),
    .Y(_4475_)
);

AOI21X1 _14579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4012_),
    .B(_4016_),
    .C(_3866_),
    .Y(_4017_)
);

NOR2X1 _14159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3540_),
    .B(_3555_),
    .Y(_3556_)
);

OAI21X1 _15940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .B(_5501_),
    .C(_5503_),
    .Y(_5507_)
);

AND2X2 _15520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf0),
    .B(breg_16_bF$buf2),
    .Y(_5046_)
);

NAND2X1 _15100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4585_),
    .B(_4586_),
    .Y(_4587_)
);

AOI21X1 _20597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10543_),
    .B(_10548_),
    .C(_10462_),
    .Y(_10613_)
);

NAND3X1 _20177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10147_),
    .B(_10151_),
    .C(_10150_),
    .Y(_10152_)
);

AOI21X1 _16725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6349_),
    .B(_6355_),
    .C(_6262_),
    .Y(_6368_)
);

INVX2 _16305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .Y(_5908_)
);

FILL SFILL59080x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9070_),
    .B(_9077_),
    .C(_9039_),
    .Y(_9078_)
);

FILL SFILL69400x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43880x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10408_),
    .B(_10375_),
    .Y(_10419_)
);

AOI21X1 _12225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3460_),
    .B(_4785_),
    .C(_4807_),
    .Y(_5815_)
);

NAND2X1 _22743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1055_),
    .B(_872_),
    .Y(_1056_)
);

NAND3X1 _22323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_579_),
    .B(_584_),
    .C(_588_),
    .Y(_596_)
);

FILL SFILL33880x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _23948_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[2]),
    .CLK(clk_bF$buf2),
    .D(_0_[2])
);

XNOR2X1 _23528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1909_),
    .B(_1901_),
    .Y(_1910_)
);

OAI21X1 _23108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1192_),
    .B(_1348_),
    .C(_1452_),
    .Y(_1453_)
);

NAND3X1 _17683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7401_),
    .B(_7406_),
    .C(_7408_),
    .Y(_7418_)
);

AOI21X1 _17263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6556_),
    .B(_6559_),
    .C(_6563_),
    .Y(_6958_)
);

FILL SFILL49000x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8738_),
    .B(_8737_),
    .C(_8736_),
    .Y(_8739_)
);

NAND2X1 _18468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8274_),
    .B(_8278_),
    .Y(_8279_)
);

AND2X2 _18048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_16_bF$buf1),
    .B(breg_16_bF$buf3),
    .Y(_7818_)
);

AOI21X1 _13183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2445_),
    .B(_2444_),
    .C(_2443_),
    .Y(_2489_)
);

OAI21X1 _23281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1630_),
    .B(_1634_),
    .C(_1636_),
    .Y(_1643_)
);

FILL SFILL23880x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _11916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2420_),
    .Y(_2431_)
);

AOI21X1 _14388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3549_),
    .B(_3545_),
    .C(_3552_),
    .Y(_3807_)
);

DFFPOSX1 _24066_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[24]),
    .CLK(clk_bF$buf4),
    .D(b[24])
);

FILL SFILL53880x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _16954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6234_),
    .B(_6618_),
    .Y(_6619_)
);

NAND3X1 _16534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6152_),
    .B(_6137_),
    .C(_6153_),
    .Y(_6158_)
);

AOI21X1 _16114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5370_),
    .B(_5697_),
    .C(_5374_),
    .Y(_5698_)
);

FILL SFILL8760x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _17739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7474_),
    .B(_7475_),
    .C(_7473_),
    .Y(_7479_)
);

NAND2X1 _17319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_18_bF$buf0),
    .Y(_7018_)
);

AOI21X1 _12874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_856_),
    .B(_900_),
    .C(_133_),
    .Y(_1020_)
);

AOI21X1 _12454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8260_),
    .B(_8271_),
    .C(_6955_),
    .Y(_8326_)
);

NAND2X1 _22972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf5),
    .B(areg_26_bF$buf0),
    .Y(_1305_)
);

AOI21X1 _12034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3712_),
    .B(_3690_),
    .C(_3558_),
    .Y(_3723_)
);

NAND2X1 _22552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_844_),
    .Y(_847_)
);

NOR3X1 _22132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_386_),
    .C(_382_),
    .Y(_387_)
);

OAI21X1 _13659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3008_),
    .B(_3007_),
    .C(_3003_),
    .Y(_3009_)
);

AOI21X1 _13239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2528_),
    .B(_2529_),
    .C(_2336_),
    .Y(_2549_)
);

AND2X2 _23757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2119_),
    .B(_2159_),
    .Y(_2160_)
);

FILL SFILL3720x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf4),
    .B(areg_29_bF$buf5),
    .Y(_1703_)
);

FILL SFILL43960x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4038_),
    .B(_4039_),
    .C(_4037_),
    .Y(_4040_)
);

NAND3X1 _17492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7208_),
    .B(_6809_),
    .C(_7202_),
    .Y(_7209_)
);

NAND3X1 _17072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6748_),
    .B(_6745_),
    .C(_6746_),
    .Y(_6749_)
);

FILL SFILL48920x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5357_),
    .B(_5358_),
    .Y(_5359_)
);

OAI21X1 _18697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8130_),
    .B(_8125_),
    .C(_8133_),
    .Y(_8529_)
);

AOI21X1 _18277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8067_),
    .B(_7652_),
    .C(_8068_),
    .Y(_8069_)
);

NAND2X1 _23090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .B(_1426_),
    .Y(_1433_)
);

FILL SFILL64360x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_44_),
    .C(_47_),
    .Y(_48_)
);

OAI21X1 _21403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10861_),
    .B(_11480_),
    .C(_11177_),
    .Y(_11497_)
);

XNOR2X1 _14197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3597_),
    .B(_3594_),
    .Y(_3598_)
);

OAI21X1 _22608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_904_),
    .C(_725_),
    .Y(_908_)
);

FILL SFILL49080x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6392_),
    .B(_6398_),
    .C(_6045_),
    .Y(_6410_)
);

NAND2X1 _16343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5927_),
    .B(_5923_),
    .Y(_5950_)
);

FILL SFILL49000x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert270 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217_),
    .Y(_7217__bF$buf3)
);

BUFX2 BUFX2_insert271 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217_),
    .Y(_7217__bF$buf2)
);

BUFX2 BUFX2_insert272 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217_),
    .Y(_7217__bF$buf1)
);

BUFX2 BUFX2_insert273 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217_),
    .Y(_7217__bF$buf0)
);

NAND3X1 _17968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7710_),
    .B(_7729_),
    .C(_7724_),
    .Y(_7730_)
);

BUFX2 BUFX2_insert274 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6050_),
    .Y(_6050__bF$buf3)
);

NAND3X1 _17548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7226_),
    .B(_7267_),
    .C(_7268_),
    .Y(_7269_)
);

BUFX2 BUFX2_insert275 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6050_),
    .Y(_6050__bF$buf2)
);

BUFX2 BUFX2_insert276 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6050_),
    .Y(_6050__bF$buf1)
);

INVX1 _17128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6793_),
    .Y(_6809_)
);

BUFX2 BUFX2_insert277 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6050_),
    .Y(_6050__bF$buf0)
);

BUFX2 BUFX2_insert278 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf4)
);

BUFX2 BUFX2_insert279 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[11]),
    .Y(areg_11_bF$buf3)
);

AND2X2 _12683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf0),
    .B(areg_11_bF$buf1),
    .Y(_10836_)
);

XOR2X1 _12263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5442_),
    .B(_6220_),
    .Y(_6231_)
);

AOI21X1 _22781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(_1081_),
    .C(_947_),
    .Y(_1097_)
);

FILL SFILL23880x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_632_),
    .B(_619_),
    .C(_631_),
    .Y(_638_)
);

FILL SFILL39080x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2765_),
    .B(_2996_),
    .C(_2995_),
    .Y(_3260_)
);

XNOR2X1 _13468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2799_),
    .B(_2795_),
    .Y(_2800_)
);

DFFPOSX1 _23986_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[40]),
    .CLK(clk_bF$buf7),
    .D(_0_[40])
);

NAND3X1 _13048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .B(_2335_),
    .C(_2337_),
    .Y(_2343_)
);

INVX1 _23566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6804_),
    .Y(_1952_)
);

NAND2X1 _23146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_23_bF$buf2),
    .B(areg_28_bF$buf2),
    .Y(_1495_)
);

FILL SFILL39000x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4888_),
    .B(_5149_),
    .C(_4878_),
    .Y(_5150_)
);

AOI21X1 _18086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7809_),
    .B(_7806_),
    .C(_7791_),
    .Y(_7860_)
);

FILL SFILL13800x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6467_),
    .B(_6468_),
    .C(_6469_),
    .Y(_6470_)
);

OAI21X1 _11954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2759_),
    .B(_2814_),
    .C(_2836_),
    .Y(_2847_)
);

XNOR2X1 _21632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11725_),
    .B(_11719_),
    .Y(_11747_)
);

OAI21X1 _21212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11266_),
    .B(_11274_),
    .C(_11279_),
    .Y(_11288_)
);

FILL SFILL29000x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74440x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8522_),
    .B(_9587_),
    .C(_11439_),
    .Y(_11450_)
);

AOI21X1 _12319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5661_),
    .B(_5683_),
    .C(_5409_),
    .Y(_6845_)
);

AOI21X1 _22837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_1050_),
    .C(_1157_),
    .Y(_1158_)
);

OAI21X1 _22417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_679_),
    .C(_686_),
    .Y(_699_)
);

FILL SFILL74360x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6653_),
    .Y(_6661_)
);

NAND3X1 _16572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6199_),
    .B(_6161_),
    .C(_6192_),
    .Y(_6200_)
);

NAND3X1 _16152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5725_),
    .B(_5730_),
    .C(_5735_),
    .Y(_5740_)
);

OAI21X1 _17777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_7520__bF$buf0),
    .C(_7517_),
    .Y(_7521_)
);

NAND3X1 _17357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7058_),
    .B(_7059_),
    .C(_7060_),
    .Y(_7061_)
);

NAND2X1 _12492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf1),
    .B(breg[8]),
    .Y(_8742_)
);

OAI21X1 _12072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf0),
    .B(_4116__bF$buf4),
    .C(_4127_),
    .Y(_4138_)
);

NAND2X1 _22590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_607_),
    .Y(_888_)
);

OR2X2 _22170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_398_),
    .Y(_428_)
);

NAND3X1 _20903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10947_),
    .B(_10945_),
    .C(_10948_),
    .Y(_10949_)
);

NOR2X1 _13697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562__bF$buf3),
    .B(_2379_),
    .Y(_3051_)
);

NAND2X1 _13277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg_9_bF$buf2),
    .Y(_2591_)
);

NAND2X1 _23795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2165_),
    .Y(_2201_)
);

NAND3X1 _23375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1736_),
    .B(_1727_),
    .C(_1732_),
    .Y(_1745_)
);

OAI21X1 _19923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9874_),
    .B(_9873_),
    .C(_9863_),
    .Y(_9875_)
);

AOI21X1 _19503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9017_),
    .B(_9021_),
    .C(_9024_),
    .Y(_9414_)
);

NOR3X1 _15843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5394_),
    .B(_5396_),
    .C(_5395_),
    .Y(_5401_)
);

AOI21X1 _15423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4931_),
    .B(_4923_),
    .C(_4673_),
    .Y(_4942_)
);

NAND3X1 _15003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4462_),
    .B(_4467_),
    .C(_4469_),
    .Y(_4481_)
);

NAND3X1 _16628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6258_),
    .B(_6259_),
    .C(_6260_),
    .Y(_6261_)
);

NOR2X1 _16208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5419_),
    .B(_5795_),
    .Y(_5801_)
);

NAND3X1 _21861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_80_),
    .C(_85_),
    .Y(_90_)
);

NAND2X1 _21441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11536_),
    .B(_11537_),
    .Y(_11539_)
);

NOR3X1 _21021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11061_),
    .B(_11064_),
    .C(_11065_),
    .Y(_11078_)
);

NOR2X1 _12968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1925_),
    .B(_2023_),
    .Y(_2045_)
);

FILL SFILL23800x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _12548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9334_),
    .B(_9301_),
    .C(_9345_),
    .Y(_9356_)
);

NAND3X1 _12128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4533_),
    .B(_4577_),
    .C(_4599_),
    .Y(_4752_)
);

NAND2X1 _22646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_882_),
    .Y(_949_)
);

AOI22X1 _22226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_477_),
    .B(_482_),
    .C(_229_),
    .D(_234_),
    .Y(_489_)
);

FILL SFILL8840x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5829_),
    .B(_5824_),
    .C(_5831_),
    .Y(_5991_)
);

FILL SFILL13880x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7295_),
    .B(_7299_),
    .C(_7307_),
    .Y(_7311_)
);

NAND2X1 _17166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg_26_bF$buf2),
    .Y(_6851_)
);

FILL SFILL74120x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10699_),
    .B(_10738_),
    .C(_10736_),
    .Y(_10739_)
);

NOR2X1 _13086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1511_),
    .B(_2381_),
    .Y(_2382_)
);

NAND2X1 _23184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1531_),
    .B(_1536_),
    .Y(_1537_)
);

AOI21X1 _19732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9659_),
    .B(_9664_),
    .C(_9651_),
    .Y(_9665_)
);

AOI21X1 _19312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9204_),
    .B(_9197_),
    .C(_9095_),
    .Y(_9205_)
);

NAND3X1 _21917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_139_),
    .C(_148_),
    .Y(_151_)
);

OAI21X1 _15652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5191_),
    .B(_5189_),
    .C(_5188_),
    .Y(_5192_)
);

AOI21X1 _15232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4476_),
    .B(_4731_),
    .C(_4729_),
    .Y(_4732_)
);

FILL SFILL64040x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6192_),
    .B(_6200_),
    .Y(_6512_)
);

NAND2X1 _16437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg_27_bF$buf5),
    .Y(_6051_)
);

NAND3X1 _16017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5513_),
    .B(_5584_),
    .C(_5591_),
    .Y(_5592_)
);

FILL SFILL64440x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _11992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3088_),
    .B(_3154_),
    .Y(_3263_)
);

NAND3X1 _21670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11763_),
    .B(_11777_),
    .C(_11766_),
    .Y(_11788_)
);

INVX1 _21250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11327_),
    .Y(_11328_)
);

NAND3X1 _12777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11745_),
    .B(_11855_),
    .C(_11811_),
    .Y(_11866_)
);

NAND2X1 _12357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6209_),
    .B(_6286_),
    .Y(_7261_)
);

INVX1 _22875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1044_),
    .Y(_1200_)
);

OAI21X1 _22455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(_509_),
    .C(_517_),
    .Y(_740_)
);

OAI21X1 _22035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_277_),
    .C(_272_),
    .Y(_280_)
);

NAND2X1 _16190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf2),
    .B(breg_16_bF$buf4),
    .Y(_5781_)
);

INVX1 _14923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4392_),
    .Y(_4393_)
);

NAND3X1 _14503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3924_),
    .B(_3928_),
    .C(_3933_),
    .Y(_3934_)
);

NOR2X1 _17395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7096_),
    .B(_7097_),
    .Y(_7103_)
);

NOR3X1 _15708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5246_),
    .B(_5247_),
    .C(_5243_),
    .Y(_5253_)
);

OAI21X1 _20941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10982_),
    .B(_10978_),
    .C(_10984_),
    .Y(_10991_)
);

NAND3X1 _20521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10520_),
    .B(_10506_),
    .C(_10510_),
    .Y(_10530_)
);

OAI21X1 _20101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10061_),
    .B(_10060_),
    .C(_10058_),
    .Y(_10069_)
);

FILL SFILL44040x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9914_),
    .B(_9555_),
    .Y(_9916_)
);

OAI21X1 _19541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9450_),
    .B(_9454_),
    .C(_9425_),
    .Y(_9456_)
);

AOI21X1 _19121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8602_),
    .B(_8681_),
    .C(_8690_),
    .Y(_8995_)
);

AOI21X1 _21726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11323_),
    .B(_11568_),
    .C(_11575_),
    .Y(_11850_)
);

NOR2X1 _21306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11072_),
    .B(_11383_),
    .Y(_11390_)
);

OAI21X1 _15881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5440_),
    .B(_5441_),
    .C(_5437_),
    .Y(_5443_)
);

NOR2X1 _15461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4978_),
    .B(_4980_),
    .Y(_4982_)
);

NOR3X1 _15041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4517_),
    .B(_4519_),
    .C(_4516_),
    .Y(_4523_)
);

NOR2X1 _16666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6296_),
    .B(_6298_),
    .Y(_6303_)
);

OAI21X1 _16246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf1),
    .B(_2465__bF$buf1),
    .C(_5468_),
    .Y(_5843_)
);

NAND3X1 _12586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6955_),
    .B(_8183_),
    .C(_8227_),
    .Y(_9773_)
);

NAND2X1 _12166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5135_),
    .B(_5157_),
    .Y(_5168_)
);

NAND3X1 _22684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_988_),
    .B(_983_),
    .C(_990_),
    .Y(_991_)
);

AOI21X1 _22264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_255_),
    .B(_280_),
    .C(_278_),
    .Y(_531_)
);

AOI21X1 _18812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8645_),
    .B(_8642_),
    .C(_8640_),
    .Y(_8656_)
);

BUFX2 _23889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[7]),
    .Y(y[7])
);

NAND3X1 _23469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1840_),
    .C(_1741_),
    .Y(_1847_)
);

FILL SFILL64120x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(_1378_),
    .C(_1381_),
    .Y(_1389_)
);

XNOR2X1 _14732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4161_),
    .B(_4156_),
    .Y(_4184_)
);

NAND3X1 _14312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3639_),
    .B(_3717_),
    .C(_3718_),
    .Y(_3725_)
);

NOR3X1 _15937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5500_),
    .B(_5501_),
    .C(_5503_),
    .Y(_5504_)
);

OAI21X1 _15517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4400_),
    .B(_5042_),
    .C(_4718_),
    .Y(_5043_)
);

NAND3X1 _20750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10742_),
    .B(_10779_),
    .C(_10774_),
    .Y(_10780_)
);

NAND3X1 _20330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10305_),
    .B(_10309_),
    .C(_10313_),
    .Y(_10320_)
);

FILL SFILL28680x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL FILL74040x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _19770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9691_),
    .B(_9694_),
    .C(_9695_),
    .Y(_9706_)
);

OAI21X1 _19350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9233_),
    .B(_9237_),
    .C(_9240_),
    .Y(_9246_)
);

FILL SFILL54120x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_192_),
    .Y(_193_)
);

NOR3X1 _21535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11638_),
    .B(_11639_),
    .C(_11640_),
    .Y(_11641_)
);

NAND2X1 _21115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf2),
    .B(areg_28_bF$buf0),
    .Y(_11181_)
);

AOI21X1 _15690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5217_),
    .B(_5222_),
    .C(_5178_),
    .Y(_5232_)
);

XNOR2X1 _15270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4772_),
    .B(_4770_),
    .Y(_4773_)
);

FILL SFILL18680x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6552_),
    .B(_6553_),
    .Y(_6554_)
);

NOR3X1 _16475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5764_),
    .B(_5766_),
    .C(_5759_),
    .Y(_6093_)
);

NAND3X1 _16055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5626_),
    .B(_5633_),
    .C(_5307_),
    .Y(_5634_)
);

FILL SFILL44040x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL54120x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7667_),
    .Y(_7678_)
);

INVX1 _22493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_776_),
    .Y(_782_)
);

NAND3X1 _22073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_317_),
    .B(_305_),
    .C(_310_),
    .Y(_322_)
);

AOI21X1 _18621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8444_),
    .B(_8445_),
    .C(_8075_),
    .Y(_8447_)
);

AND2X2 _18201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7949_),
    .B(_7954_),
    .Y(_7987_)
);

NAND3X1 _20806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10835_),
    .B(_10837_),
    .C(_10841_),
    .Y(_10842_)
);

XNOR2X1 _23698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2095_),
    .B(_2063_),
    .Y(_2096_)
);

NAND3X1 _23278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1637_),
    .B(_1638_),
    .C(_1636_),
    .Y(_1639_)
);

AND2X2 _19826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf5),
    .B(breg_19_bF$buf3),
    .Y(_9768_)
);

AOI21X1 _19406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9306_),
    .B(_9303_),
    .C(_9281_),
    .Y(_9307_)
);

AOI21X1 _14961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4430_),
    .B(_4429_),
    .C(_4428_),
    .Y(_4435_)
);

FILL SFILL69240x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3974_),
    .B(_3973_),
    .C(_3957_),
    .Y(_3976_)
);

NOR2X1 _14121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3510_),
    .B(_2979_),
    .Y(_3515_)
);

FILL SFILL69160x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5293_),
    .B(_4948_),
    .C(_5294_),
    .Y(_5295_)
);

AOI21X1 _15326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4826_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4835_)
);

FILL SFILL38760x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _21764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11890_),
    .Y(_11891_)
);

OAI21X1 _21344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11429_),
    .B(_11427_),
    .C(_11431_),
    .Y(_11432_)
);

FILL SFILL38680x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64360x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64280x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1144_),
    .B(_1301_),
    .C(_1300_),
    .Y(_1302_)
);

FILL SFILL64120x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _22549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_26_bF$buf0),
    .C(breg_22_bF$buf4),
    .D(areg_25_bF$buf1),
    .Y(_843_)
);

NAND2X1 _22129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_18_bF$buf3),
    .B(areg_27_bF$buf0),
    .Y(_383_)
);

AOI21X1 _13812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3177_),
    .B(_3170_),
    .C(_3127_),
    .Y(_3178_)
);

BUFX2 _23910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[28]),
    .Y(y[28])
);

AOI21X1 _16284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5577_),
    .B(_5572_),
    .C(_5542_),
    .Y(_5885_)
);

FILL FILL74120x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _17489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7197_),
    .Y(_7205_)
);

NAND2X1 _17069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6743_),
    .B(_6744_),
    .Y(_6745_)
);

FILL SFILL18760x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL14040x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _18850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8696_),
    .Y(_8697_)
);

OAI21X1 _18430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf4),
    .B(_3958__bF$buf3),
    .C(_7838_),
    .Y(_8237_)
);

NAND3X1 _18010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7760_),
    .B(_7764_),
    .C(_7772_),
    .Y(_7776_)
);

FILL SFILL54120x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10627_),
    .B(_10626_),
    .C(_10625_),
    .Y(_10633_)
);

NOR2X1 _23087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1428_),
    .B(_1429_),
    .Y(_1430_)
);

AOI21X1 _19635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9544_),
    .B(_9539_),
    .C(_9530_),
    .Y(_9559_)
);

NAND2X1 _19215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8725_),
    .B(_8730_),
    .Y(_9097_)
);

INVX1 _14770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3952_),
    .Y(_4225_)
);

OAI21X1 _14350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3762_),
    .B(_3765_),
    .C(_3487_),
    .Y(_3766_)
);

FILL SFILL59320x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf1),
    .B(areg_23_bF$buf1),
    .Y(_5546_)
);

NAND2X1 _15555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5081_),
    .B(_5084_),
    .Y(_5085_)
);

OAI21X1 _15135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4622_),
    .B(_4623_),
    .C(_4352_),
    .Y(_4626_)
);

NAND2X1 _21993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_229_),
    .Y(_235_)
);

NOR3X1 _21573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11460_),
    .B(_11458_),
    .C(_11454_),
    .Y(_11682_)
);

OAI21X1 _21153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11214_),
    .B(_11215_),
    .C(_11212_),
    .Y(_11223_)
);

AND2X2 _17701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7044_),
    .B(_7038_),
    .Y(_7438_)
);

XNOR2X1 _22778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_1093_),
    .Y(_0_[48])
);

AOI21X1 _22358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_630_),
    .C(_616_),
    .Y(_634_)
);

INVX4 _18906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_30_bF$buf5),
    .Y(_8759_)
);

FILL SFILL69240x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2752_),
    .B(_2967_),
    .C(_2964_),
    .Y(_2969_)
);

AOI21X1 _13201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1881_),
    .B(_2321_),
    .C(_2507_),
    .Y(_2509_)
);

OAI21X1 _16093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4973_),
    .B(_5674_),
    .C(_5317_),
    .Y(_5675_)
);

NAND3X1 _14826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4280_),
    .B(_4286_),
    .C(_4200_),
    .Y(_4287_)
);

OAI21X1 _14406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf1),
    .B(_2560__bF$buf4),
    .C(_3813_),
    .Y(_3827_)
);

FILL SFILL29000x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6995_),
    .B(_6994_),
    .C(_6991_),
    .Y(_6996_)
);

FILL SFILL69160x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8520x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10860_),
    .B(_10874_),
    .C(_10864_),
    .Y(_10884_)
);

OAI21X1 _20424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10116_),
    .B(_10184_),
    .C(_10138_),
    .Y(_10423_)
);

OAI21X1 _20004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9946_),
    .B(_9953_),
    .C(_9956_),
    .Y(_9963_)
);

AOI21X1 _19864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9799_),
    .B(_9798_),
    .C(_9796_),
    .Y(_9810_)
);

NAND3X1 _19444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9342_),
    .B(_9347_),
    .C(_9348_),
    .Y(_9349_)
);

INVX2 _19024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8887_),
    .Y(_8888_)
);

FILL SFILL24040x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11733_),
    .B(_11730_),
    .C(_11728_),
    .Y(_11743_)
);

NAND3X1 _21209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11280_),
    .B(_11283_),
    .C(_11279_),
    .Y(_11284_)
);

NAND3X1 _15784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5333_),
    .B(_5334_),
    .C(_5335_),
    .Y(_5336_)
);

NAND3X1 _15364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4874_),
    .B(_4876_),
    .C(_4875_),
    .Y(_4877_)
);

NAND2X1 _16989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6654_),
    .B(_6655_),
    .Y(_6656_)
);

AOI21X1 _16569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6194_),
    .B(_6195_),
    .C(_6188_),
    .Y(_6196_)
);

OAI21X1 _16149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5733_),
    .B(_5734_),
    .C(_5735_),
    .Y(_5736_)
);

AND2X2 _21382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf0),
    .B(areg_26_bF$buf4),
    .Y(_11474_)
);

FILL SFILL18760x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33560x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7686_),
    .B(_7687_),
    .C(_7672_),
    .Y(_7688_)
);

INVX1 _17510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7226_),
    .Y(_7227_)
);

FILL SFILL33960x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7964_),
    .B(_7986_),
    .C(_7876_),
    .Y(_8709_)
);

INVX2 _12069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4094_),
    .Y(_4105_)
);

NAND3X1 _22587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_882_),
    .C(_883_),
    .Y(_885_)
);

NAND3X1 _22167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_402_),
    .B(_415_),
    .C(_412_),
    .Y(_425_)
);

OAI21X1 _18715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10869__bF$buf1),
    .B(_3781__bF$buf2),
    .C(_8191_),
    .Y(_8549_)
);

NAND3X1 _13850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3215_),
    .B(_3216_),
    .C(_2987_),
    .Y(_3219_)
);

AOI21X1 _13430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2710_),
    .C(_2579_),
    .Y(_2758_)
);

AOI21X1 _13010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2299_),
    .B(_2304_),
    .C(_2142_),
    .Y(_2305_)
);

NOR2X1 _14635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3790_),
    .B(_4076_),
    .Y(_4077_)
);

NAND3X1 _14215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3599_),
    .B(_3614_),
    .C(_3617_),
    .Y(_3618_)
);

FILL SFILL23960x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9987_),
    .B(_10673_),
    .Y(_10674_)
);

XOR2X1 _20233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10157_),
    .B(_10212_),
    .Y(_10213_)
);

AOI21X1 _19673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9224_),
    .B(_9222_),
    .C(_9600_),
    .Y(_9601_)
);

OAI21X1 _19253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9139_),
    .B(_9138_),
    .C(_9136_),
    .Y(_9140_)
);

OAI21X1 _21858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_84_),
    .B(_83_),
    .C(_85_),
    .Y(_86_)
);

NAND2X1 _21438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11532_),
    .B(_11534_),
    .Y(_11535_)
);

OAI22X1 _21018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10466_),
    .B(_11072_),
    .C(_11073_),
    .D(_10816_),
    .Y(_11074_)
);

AOI21X1 _12701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10891_),
    .B(_10935_),
    .C(_10803_),
    .Y(_11043_)
);

AOI21X1 _15593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5116_),
    .B(_5115_),
    .C(_5111_),
    .Y(_5127_)
);

OAI21X1 _15173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4353_),
    .B(_4095_),
    .C(_4666_),
    .Y(_4667_)
);

NOR2X1 _13906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2768_),
    .B(_2993_),
    .Y(_3280_)
);

AND2X2 _16798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_24_bF$buf5),
    .Y(_6447_)
);

OAI21X1 _16378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5985_),
    .B(_5986_),
    .C(_5984_),
    .Y(_5987_)
);

NAND2X1 _21191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11262_),
    .B(_11263_),
    .Y(_11265_)
);

FILL SFILL59240x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6516_),
    .B(_6604_),
    .Y(_6615_)
);

INVX1 _22396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_448_),
    .Y(_675_)
);

AOI21X1 _18944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8799_),
    .B(_8800_),
    .C(_8798_),
    .Y(_8801_)
);

OAI21X1 _18524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_7100__bF$buf3),
    .C(_8333_),
    .Y(_8341_)
);

OAI21X1 _18104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7578_),
    .B(_7879_),
    .C(_7566_),
    .Y(_7880_)
);

OAI21X1 _20709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10734_),
    .B(_10730_),
    .C(_10700_),
    .Y(_10735_)
);

FILL FILL74200x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _19729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9293_),
    .B(_9660_),
    .Y(_9661_)
);

AOI21X1 _19309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9176_),
    .B(_9183_),
    .C(_9193_),
    .Y(_9201_)
);

NAND3X1 _14864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4316_),
    .B(_4320_),
    .C(_4322_),
    .Y(_4329_)
);

NOR2X1 _14444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf0),
    .B(_2379_),
    .Y(_3869_)
);

NOR2X1 _14024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3399_),
    .B(_3400_),
    .Y(_3409_)
);

FILL SFILL33640x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _15649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5182_),
    .Y(_5188_)
);

AOI21X1 _15229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4717_),
    .B(_4716_),
    .C(_4713_),
    .Y(_4728_)
);

NAND3X1 _20882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10917_),
    .B(_10923_),
    .C(_10925_),
    .Y(_10926_)
);

INVX2 _20462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10464_),
    .Y(_10465_)
);

NOR2X1 _20042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5190__bF$buf1),
    .B(_6815__bF$buf2),
    .Y(_10004_)
);

NAND2X1 _19482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9080_),
    .B(_9085_),
    .Y(_9391_)
);

OAI21X1 _19062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8926_),
    .B(_8925_),
    .C(_8924_),
    .Y(_8930_)
);

FILL SFILL33960x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _11989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_2376__bF$buf0),
    .Y(_3231_)
);

NAND3X1 _21667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11753_),
    .B(_11780_),
    .C(_11784_),
    .Y(_11785_)
);

OAI21X1 _21247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11130_),
    .B(_11282_),
    .C(_11272_),
    .Y(_11325_)
);

XNOR2X1 _12930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1620_),
    .B(_1586_),
    .Y(_1631_)
);

NAND2X1 _12510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8928_),
    .B(_8895_),
    .Y(_8939_)
);

NAND2X1 _13715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf4),
    .B(breg_10_bF$buf3),
    .Y(_3071_)
);

NAND2X1 _23813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2180_),
    .B(_2178_),
    .Y(_2220_)
);

AOI21X1 _16187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5777_),
    .B(_5776_),
    .C(_5775_),
    .Y(_5778_)
);

FILL SFILL69400x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8188_),
    .B(_8268_),
    .C(_8277_),
    .Y(_8591_)
);

OAI21X1 _18333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8130_),
    .B(_8129_),
    .C(_8125_),
    .Y(_8131_)
);

FILL SFILL69320x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10986_),
    .B(_10985_),
    .C(_10984_),
    .Y(_10987_)
);

OAI21X1 _20518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10524_),
    .B(_10525_),
    .C(_10523_),
    .Y(_10526_)
);

XNOR2X1 _19958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9911_),
    .B(_9902_),
    .Y(_9912_)
);

NAND3X1 _19538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9435_),
    .B(_9438_),
    .C(_9448_),
    .Y(_9452_)
);

NAND3X1 _19118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8989_),
    .B(_8990_),
    .C(_8985_),
    .Y(_8991_)
);

AOI21X1 _14673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4104_),
    .B(_4103_),
    .C(_4100_),
    .Y(_4119_)
);

OAI21X1 _14253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3655_),
    .B(_3656_),
    .C(_3659_),
    .Y(_3660_)
);

OAI21X1 _15878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5424_),
    .B(_5425_),
    .C(_5422_),
    .Y(_5439_)
);

NOR2X1 _15458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4977_),
    .B(_4976_),
    .Y(_4978_)
);

AOI22X1 _15038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4238_),
    .C(_4518_),
    .D(_4261_),
    .Y(_4519_)
);

FILL SFILL59320x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10708_),
    .B(_10709_),
    .Y(_10716_)
);

OAI21X1 _20271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9901_),
    .B(_9905_),
    .C(_9908_),
    .Y(_10256_)
);

INVX1 _19291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9175_),
    .Y(_9182_)
);

OAI21X1 _21896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11765_),
    .B(_11771_),
    .C(_11760_),
    .Y(_128_)
);

OAI21X1 _21476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11575_),
    .B(_11576_),
    .C(_11324_),
    .Y(_11577_)
);

AOI21X1 _21056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10889_),
    .B(_10894_),
    .C(_10896_),
    .Y(_11116_)
);

AOI21X1 _17604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7314_),
    .B(_7320_),
    .C(_7270_),
    .Y(_7331_)
);

AOI21X1 _18809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8285_),
    .B(_8651_),
    .C(_8650_),
    .Y(_8652_)
);

INVX1 _13944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3321_),
    .Y(_3322_)
);

NAND3X1 _13524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2843_),
    .B(_2856_),
    .C(_2861_),
    .Y(_2862_)
);

NAND3X1 _13104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2397_),
    .C(_2401_),
    .Y(_2402_)
);

NOR2X1 _23622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1886_),
    .B(_2013_),
    .Y(_2014_)
);

NOR2X1 _23202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf4),
    .B(_7225__bF$buf2),
    .Y(_1556_)
);

AOI21X1 _14729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4169_),
    .B(_4168_),
    .C(_4165_),
    .Y(_4180_)
);

OAI21X1 _14309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3636_),
    .B(_3634_),
    .C(_3593_),
    .Y(_3721_)
);

NAND2X1 _18982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8841_),
    .B(_8840_),
    .Y(_8842_)
);

AND2X2 _18562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8374_),
    .B(_8378_),
    .Y(_8382_)
);

AND2X2 _18142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7464_),
    .B(_7456_),
    .Y(_7922_)
);

NOR3X1 _20747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10480_),
    .B(_10482_),
    .C(_10476_),
    .Y(_10777_)
);

NAND3X1 _20327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9993_),
    .B(_10311_),
    .C(_10316_),
    .Y(_10317_)
);

OAI22X1 _19767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9009_),
    .B(_9702_),
    .C(_9393_),
    .D(_9396_),
    .Y(_9703_)
);

NAND3X1 _19347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9241_),
    .B(_9242_),
    .C(_9240_),
    .Y(_9243_)
);

NOR3X1 _14482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3894_),
    .B(_3900_),
    .C(_3901_),
    .Y(_3911_)
);

NAND3X1 _14062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3443_),
    .B(_3450_),
    .C(_3310_),
    .Y(_3451_)
);

FILL SFILL8680x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _15687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4882_),
    .B(_4881_),
    .C(_4880_),
    .Y(_5229_)
);

NAND2X1 _15267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf1),
    .B(breg_14_bF$buf2),
    .Y(_4770_)
);

FILL SFILL69000x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_12_bF$buf4),
    .B(breg_26_bF$buf3),
    .Y(_10045_)
);

FILL SFILL8600x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11327_),
    .B(_11366_),
    .C(_11365_),
    .Y(_11367_)
);

NAND3X1 _17833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7582_),
    .B(_7436_),
    .C(_7573_),
    .Y(_7583_)
);

NAND3X1 _17413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_30_bF$buf5),
    .C(_7122_),
    .Y(_7123_)
);

FILL SFILL74280x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8437_),
    .B(_8442_),
    .C(_8076_),
    .Y(_8443_)
);

OAI22X1 _13753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_3111_),
    .C(_3112_),
    .D(_2871_),
    .Y(_3113_)
);

NOR2X1 _13333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf0),
    .B(_9104__bF$buf1),
    .Y(_2653_)
);

INVX1 _23851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .Y(_2260_)
);

OAI21X1 _23431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1714_),
    .B(_1713_),
    .C(_1804_),
    .Y(_1806_)
);

NAND2X1 _23011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_21_bF$buf3),
    .B(areg_29_bF$buf1),
    .Y(_1348_)
);

FILL SFILL74200x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4430_),
    .B(_4429_),
    .C(_4428_),
    .Y(_4431_)
);

NAND2X1 _14538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_21_bF$buf1),
    .Y(_3972_)
);

NAND2X1 _14118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3491_),
    .B(_3239_),
    .Y(_3511_)
);

FILL SFILL69480x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8616_),
    .B(_8619_),
    .C(_8622_),
    .Y(_8633_)
);

OAI21X1 _18371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7874_),
    .B(_7873_),
    .C(_7871_),
    .Y(_8173_)
);

FILL SFILL64280x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI22X1 _20976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf1),
    .B(_6050__bF$buf3),
    .C(_2287__bF$buf1),
    .D(_5668__bF$buf5),
    .Y(_11028_)
);

INVX2 _20556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10567_),
    .Y(_10568_)
);

NAND3X1 _20136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10104_),
    .B(_10105_),
    .C(_10106_),
    .Y(_10107_)
);

OAI21X1 _19996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9946_),
    .B(_9953_),
    .C(_9644_),
    .Y(_9954_)
);

NAND2X1 _19576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9492_),
    .B(_9493_),
    .Y(_9494_)
);

NAND3X1 _19156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9028_),
    .B(_9032_),
    .C(_9013_),
    .Y(_9033_)
);

NOR3X1 _14291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3417_),
    .B(_3412_),
    .C(_3415_),
    .Y(_3702_)
);

FILL SFILL33720x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9477_),
    .B(_9521_),
    .C(_8544_),
    .Y(_9970_)
);

INVX1 _22702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_980_),
    .Y(_1011_)
);

NAND2X1 _15496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_20_bF$buf2),
    .Y(_5020_)
);

NAND3X1 _15076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4550_),
    .B(_4543_),
    .C(_4548_),
    .Y(_4561_)
);

AOI21X1 _13809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3158_),
    .B(_3162_),
    .C(_3140_),
    .Y(_3174_)
);

BUFX2 _23907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[25]),
    .Y(y[25])
);

OAI21X1 _21094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11157_),
    .B(_11156_),
    .C(_11140_),
    .Y(_11158_)
);

INVX2 _17642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7345_),
    .Y(_7373_)
);

OAI21X1 _17222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6909_),
    .B(_6910_),
    .C(_6912_),
    .Y(_6913_)
);

FILL SFILL74040x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_557_),
    .C(_555_),
    .Y(_569_)
);

OAI21X1 _18847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8330_),
    .B(_8693_),
    .C(_8405_),
    .Y(_8694_)
);

OAI21X1 _18427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_3146__bF$buf1),
    .C(_8224_),
    .Y(_8234_)
);

OAI21X1 _18007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7769_),
    .B(_7770_),
    .C(_7772_),
    .Y(_7773_)
);

INVX1 _13982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3362_),
    .Y(_3363_)
);

OAI21X1 _13562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2892_),
    .C(_2877_),
    .Y(_2904_)
);

NAND2X1 _13142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2439_),
    .B(_2430_),
    .Y(_2444_)
);

AND2X2 _23660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_1998_),
    .Y(_2054_)
);

INVX1 _23240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .Y(_1597_)
);

NAND3X1 _14767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4213_),
    .B(_4217_),
    .C(_4221_),
    .Y(_4222_)
);

NAND3X1 _14347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3757_),
    .B(_3519_),
    .C(_3760_),
    .Y(_3763_)
);

DFFPOSX1 _24025_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[15]),
    .CLK(clk_bF$buf5),
    .D(a[15])
);

FILL SFILL8600x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7960_),
    .B(_7961_),
    .C(_7962_),
    .Y(_7963_)
);

XOR2X1 _20785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10755_),
    .B(_10818_),
    .Y(_10819_)
);

INVX2 _20365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10357_),
    .Y(_10358_)
);

NAND3X1 _16913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6569_),
    .B(_6556_),
    .C(_6559_),
    .Y(_6574_)
);

OAI21X1 _19385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8909_),
    .B(_8899_),
    .C(_8903_),
    .Y(_9284_)
);

FILL SFILL44040x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(_560_),
    .C(_538_),
    .Y(_571_)
);

NAND3X1 _12413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7821_),
    .B(_7865_),
    .C(_7558_),
    .Y(_7876_)
);

AOI21X1 _22931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1259_),
    .B(_942_),
    .C(_1257_),
    .Y(_1261_)
);

NAND3X1 _22511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_800_),
    .C(_798_),
    .Y(_802_)
);

OAI21X1 _13618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2961_),
    .B(_2962_),
    .C(_2755_),
    .Y(_2965_)
);

AOI21X1 _23716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .B(_942_),
    .C(_2114_),
    .Y(_2115_)
);

AOI21X1 _17871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6811_),
    .B(_7195_),
    .C(_7199_),
    .Y(_7625_)
);

NOR3X1 _17451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6739_),
    .B(_6740_),
    .C(_6738_),
    .Y(_7165_)
);

NAND2X1 _17031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf5),
    .B(areg_28_bF$buf3),
    .Y(_6704_)
);

FILL SFILL28840x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _18656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2792_),
    .B(_7225__bF$buf3),
    .Y(_8484_)
);

NAND3X1 _18236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8022_),
    .B(_8023_),
    .C(_8021_),
    .Y(_8024_)
);

AOI21X1 _13791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3153_),
    .B(_3151_),
    .C(_3150_),
    .Y(_3155_)
);

OAI21X1 _13371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_2690_),
    .C(_2686_),
    .Y(_2695_)
);

AOI21X1 _14996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4470_),
    .B(_4471_),
    .C(_4455_),
    .Y(_4472_)
);

NAND3X1 _14576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4009_),
    .B(_4010_),
    .C(_4007_),
    .Y(_4014_)
);

FILL SFILL13800x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3549_),
    .B(_3545_),
    .C(_3552_),
    .Y(_3553_)
);

FILL SFILL13720x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10535_),
    .B(_10539_),
    .C(_10547_),
    .Y(_10610_)
);

AND2X2 _20174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf5),
    .B(areg_23_bF$buf1),
    .Y(_10149_)
);

NOR3X1 _16722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5972_),
    .B(_5973_),
    .C(_5971_),
    .Y(_6365_)
);

AOI21X1 _16302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5544_),
    .B(_5548_),
    .C(_5550_),
    .Y(_5905_)
);

AOI21X1 _19194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9048_),
    .B(_9052_),
    .C(_9062_),
    .Y(_9075_)
);

FILL SFILL23720x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11892_),
    .B(_13_),
    .C(_9_),
    .Y(_21_)
);

AOI21X1 _21379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11468_),
    .B(_11469_),
    .C(_11467_),
    .Y(_11470_)
);

AOI21X1 _17927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7236_),
    .B(_7241_),
    .C(_7244_),
    .Y(_7685_)
);

AND2X2 _17507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6902_),
    .B(_6894_),
    .Y(_7224_)
);

OAI21X1 _12642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10342_),
    .B(_10332_),
    .C(_10353_),
    .Y(_10386_)
);

NAND3X1 _12222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5694_),
    .B(_5651_),
    .C(_4992_),
    .Y(_5792_)
);

XNOR2X1 _22740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1051_),
    .B(_1040_),
    .Y(_1052_)
);

NAND3X1 _22320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_591_),
    .C(_540_),
    .Y(_592_)
);

FILL SFILL48920x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3195_),
    .B(_3203_),
    .C(_3047_),
    .Y(_3216_)
);

BUFX2 _23945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[63]),
    .Y(y[63])
);

OAI21X1 _13427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2754_),
    .B(_2553_),
    .C(_2722_),
    .Y(_2755_)
);

NOR2X1 _13007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2238_),
    .B(_2301_),
    .Y(_2302_)
);

AOI21X1 _23525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_24_bF$buf4),
    .B(areg_31_bF$buf4),
    .C(_1906_),
    .Y(_1907_)
);

NAND3X1 _23105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1447_),
    .B(_1442_),
    .C(_1449_),
    .Y(_1450_)
);

FILL SFILL13720x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7413_),
    .B(_7378_),
    .C(_7407_),
    .Y(_7414_)
);

OAI21X1 _17260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6940_),
    .B(_6945_),
    .C(_6947_),
    .Y(_6954_)
);

AND2X2 _18885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8319_),
    .B(_8312_),
    .Y(_8736_)
);

AOI21X1 _18465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8269_),
    .B(_8270_),
    .C(_8272_),
    .Y(_8276_)
);

OAI21X1 _18045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7813_),
    .B(_7814_),
    .C(_7812_),
    .Y(_7815_)
);

AOI21X1 _13180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .B(_2473_),
    .C(_2456_),
    .Y(_2485_)
);

INVX1 _11913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2387_),
    .Y(_2398_)
);

FILL SFILL38840x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3793_),
    .B(_3797_),
    .C(_3786_),
    .Y(_3804_)
);

DFFPOSX1 _24063_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[21]),
    .CLK(clk_bF$buf1),
    .D(b[21])
);

OAI22X1 _16951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6044__bF$buf0),
    .B(_3958__bF$buf1),
    .C(_7217__bF$buf1),
    .D(_3402__bF$buf3),
    .Y(_6616_)
);

NAND3X1 _16531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6151_),
    .B(_6152_),
    .C(_6153_),
    .Y(_6155_)
);

AOI21X1 _16111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5692_),
    .B(_5693_),
    .C(_5691_),
    .Y(_5695_)
);

FILL SFILL28840x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10953_),
    .B(_10954_),
    .Y(_11261_)
);

OAI21X1 _17736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7473_),
    .B(_7474_),
    .C(_7475_),
    .Y(_7476_)
);

OAI21X1 _17316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6745_),
    .B(_7014_),
    .C(_6735_),
    .Y(_7015_)
);

OAI21X1 _12871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_889_),
    .B(_878_),
    .C(_144_),
    .Y(_987_)
);

AOI21X1 _12451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7043_),
    .B(_6012_),
    .C(_7065_),
    .Y(_8293_)
);

NAND2X1 _12031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3612_),
    .B(_3679_),
    .Y(_3690_)
);

INVX1 _13656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2992_),
    .Y(_3006_)
);

NAND3X1 _13236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2523_),
    .C(_2526_),
    .Y(_2546_)
);

NAND2X1 _23754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2122_),
    .B(_2154_),
    .Y(_2157_)
);

INVX1 _23334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .Y(_1700_)
);

FILL SFILL18840x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5355_),
    .B(_5353_),
    .Y(_5356_)
);

AOI21X1 _18694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8148_),
    .B(_8144_),
    .C(_8149_),
    .Y(_8526_)
);

NAND2X1 _18274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8058_),
    .B(_8066_),
    .Y(_8067_)
);

NAND3X1 _20879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10918_),
    .B(_10921_),
    .C(_10920_),
    .Y(_10922_)
);

OAI21X1 _20459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10279_),
    .B(_10281_),
    .C(_10271_),
    .Y(_10461_)
);

NOR2X1 _20039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf3),
    .B(_7225__bF$buf3),
    .Y(_10000_)
);

NOR3X1 _21820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_29_),
    .B(_33_),
    .C(_32_),
    .Y(_44_)
);

OAI22X1 _21400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10912_),
    .B(_11228_),
    .C(_11492_),
    .D(_11226_),
    .Y(_11493_)
);

NAND3X1 _19899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9757_),
    .B(_9847_),
    .C(_9842_),
    .Y(_9848_)
);

NAND2X1 _19479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9382_),
    .B(_9386_),
    .Y(_9387_)
);

NOR3X1 _19059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8911_),
    .B(_8897_),
    .C(_8918_),
    .Y(_8926_)
);

NAND2X1 _14194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf1),
    .B(breg_13_bF$buf3),
    .Y(_3595_)
);

FILL SFILL69080x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48920x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf0),
    .B(breg_10_bF$buf3),
    .Y(_1598_)
);

NAND2X1 _12507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8874_),
    .B(_8863_),
    .Y(_8906_)
);

NAND3X1 _22605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_902_),
    .C(_728_),
    .Y(_905_)
);

NAND3X1 _15399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4914_),
    .B(_4907_),
    .C(_4766_),
    .Y(_4915_)
);

OAI21X1 _16760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6397_),
    .B(_6395_),
    .C(_6047_),
    .Y(_6406_)
);

AOI21X1 _16340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5935_),
    .B(_5933_),
    .C(_5931_),
    .Y(_5946_)
);

FILL SFILL34200x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert240 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf2)
);

BUFX2 BUFX2_insert241 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf1)
);

BUFX2 BUFX2_insert242 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[17]),
    .Y(areg_17_bF$buf0)
);

BUFX2 BUFX2_insert243 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf5)
);

OAI21X1 _17965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf0),
    .B(_3781__bF$buf2),
    .C(_7286_),
    .Y(_7727_)
);

BUFX2 BUFX2_insert244 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf4)
);

BUFX2 BUFX2_insert245 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf3)
);

OAI21X1 _17545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7259_),
    .B(_7265_),
    .C(_7227_),
    .Y(_7266_)
);

BUFX2 BUFX2_insert246 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf2)
);

INVX1 _17125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6805_),
    .Y(_6806_)
);

BUFX2 BUFX2_insert247 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf1)
);

BUFX2 BUFX2_insert248 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[27]),
    .Y(breg_27_bF$buf0)
);

FILL SFILL59080x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9159_),
    .B(_9049_),
    .C(_9103_),
    .Y(_10803_)
);

BUFX2 BUFX2_insert249 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[14]),
    .Y(areg_14_bF$buf4)
);

OAI22X1 _12260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4281_),
    .B(_6187_),
    .C(_5025_),
    .D(_5069_),
    .Y(_6198_)
);

FILL SFILL38920x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _13885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3256_),
    .Y(_3257_)
);

DFFPOSX1 _23983_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[37]),
    .CLK(clk_bF$buf3),
    .D(_0_[37])
);

NAND2X1 _13465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_13_bF$buf0),
    .Y(_2797_)
);

OAI21X1 _13045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2338_),
    .B(_2339_),
    .C(_2337_),
    .Y(_2340_)
);

INVX1 _23563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .Y(_1950_)
);

NAND3X1 _23143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1482_),
    .C(_1477_),
    .Y(_1492_)
);

FILL SFILL3560x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28920x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5143_),
    .B(_5144_),
    .C(_5145_),
    .Y(_5147_)
);

OAI21X1 _18083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7807_),
    .B(_7808_),
    .C(_7793_),
    .Y(_7857_)
);

NAND3X1 _20688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10707_),
    .B(_10711_),
    .C(_10710_),
    .Y(_10712_)
);

NAND3X1 _20268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10246_),
    .B(_10238_),
    .C(_10243_),
    .Y(_10252_)
);

AOI21X1 _16816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5679_),
    .B(_6446_),
    .C(_6074_),
    .Y(_6467_)
);

NAND2X1 _11951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf1),
    .B(breg_1_bF$buf3),
    .Y(_2814_)
);

NOR3X1 _19288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9162_),
    .B(_9158_),
    .C(_9161_),
    .Y(_9178_)
);

NAND3X1 _12736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9981_),
    .B(_11406_),
    .C(_11362_),
    .Y(_11417_)
);

AOI21X1 _12316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6658_),
    .B(_6692_),
    .C(_6352_),
    .Y(_6812_)
);

NAND2X1 _22834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1154_),
    .Y(_1155_)
);

NAND3X1 _22414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_686_),
    .C(_695_),
    .Y(_696_)
);

FILL SFILL18840x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _23619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_2009_),
    .Y(_2010_)
);

NAND2X1 _17774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_28_bF$buf5),
    .Y(_7518_)
);

NAND2X1 _17354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6622_),
    .B(_6630_),
    .Y(_7058_)
);

FILL SFILL74360x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10579_),
    .B(_10574_),
    .Y(_10945_)
);

AOI21X1 _18979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8838_),
    .B(_8833_),
    .C(_8598_),
    .Y(_8839_)
);

NAND2X1 _18559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8374_),
    .B(_8378_),
    .Y(_8379_)
);

OAI21X1 _18139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7509_),
    .B(_7487_),
    .C(_7500_),
    .Y(_7918_)
);

AOI21X1 _13694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2918_),
    .B(_2909_),
    .C(_2841_),
    .Y(_3048_)
);

XOR2X1 _23792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2197_),
    .B(_2168_),
    .Y(_2198_)
);

INVX1 _13274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2587_),
    .Y(_2588_)
);

OAI21X1 _23372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1741_),
    .B(_1737_),
    .C(_1622_),
    .Y(_1742_)
);

NAND2X1 _19920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_28_bF$buf1),
    .Y(_9871_)
);

NOR2X1 _19500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9403_),
    .B(_9404_),
    .Y(_9410_)
);

XNOR2X1 _14899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4365_),
    .B(_4363_),
    .Y(_4366_)
);

NAND3X1 _14479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3868_),
    .B(_3902_),
    .C(_3906_),
    .Y(_3907_)
);

NOR3X1 _14059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3440_),
    .B(_3441_),
    .C(_3436_),
    .Y(_3447_)
);

FILL SFILL3720x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5395_),
    .B(_5396_),
    .C(_5394_),
    .Y(_5397_)
);

NOR3X1 _15420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4609_),
    .B(_4611_),
    .C(_4608_),
    .Y(_4938_)
);

INVX2 _15000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4449_),
    .Y(_4476_)
);

FILL SFILL3640x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf4),
    .B(areg_24_bF$buf2),
    .Y(_10503_)
);

OAI21X1 _20077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9726_),
    .B(_9724_),
    .C(_9717_),
    .Y(_10042_)
);

AND2X2 _16625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5866_),
    .B(_5858_),
    .Y(_6258_)
);

NAND3X1 _16205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5789_),
    .B(_5794_),
    .C(_5797_),
    .Y(_5798_)
);

FILL SFILL59080x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8962_),
    .B(_8963_),
    .C(_8960_),
    .Y(_8968_)
);

FILL SFILL69400x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf3),
    .B(areg_8_bF$buf4),
    .Y(_2012_)
);

NAND3X1 _12545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9192_),
    .B(_9126_),
    .C(_9170_),
    .Y(_9323_)
);

OAI21X1 _12125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3723_),
    .B(_3756_),
    .C(_3788_),
    .Y(_4719_)
);

OAI21X1 _22643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .B(_734_),
    .C(_766_),
    .Y(_946_)
);

NOR3X1 _22223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_476_),
    .C(_479_),
    .Y(_486_)
);

XNOR2X1 _23848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2256_),
    .Y(_0_[61])
);

XOR2X1 _23428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1801_),
    .B(_1782_),
    .Y(_1802_)
);

NAND3X1 _23008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1343_),
    .C(_1341_),
    .Y(_1344_)
);

FILL SFILL49080x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7303_),
    .B(_7304_),
    .C(_7307_),
    .Y(_7308_)
);

NAND2X1 _17163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6458_),
    .B(_6466_),
    .Y(_6848_)
);

FILL SFILL18600x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49000x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8628_),
    .B(_8620_),
    .C(_8607_),
    .Y(_8629_)
);

OAI21X1 _18368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8164_),
    .B(_8165_),
    .C(_8122_),
    .Y(_8169_)
);

INVX4 _13083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf3),
    .Y(_2379_)
);

OAI21X1 _23181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_1528_),
    .C(_1527_),
    .Y(_1534_)
);

FILL SFILL23880x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_11815_),
    .C(_147_),
    .Y(_148_)
);

OAI21X1 _14288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3688_),
    .B(_3683_),
    .C(_3691_),
    .Y(_3698_)
);

FILL SFILL53880x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6508_),
    .B(_6503_),
    .Y(_6509_)
);

AND2X2 _16434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5725_),
    .B(_5718_),
    .Y(_6048_)
);

OAI21X1 _16014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5581_),
    .B(_5582_),
    .C(_5542_),
    .Y(_5589_)
);

OAI21X1 _17639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7359_),
    .B(_7356_),
    .C(_7353_),
    .Y(_7369_)
);

AOI21X1 _17219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6904_),
    .B(_6905_),
    .C(_6903_),
    .Y(_6909_)
);

INVX1 _12774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11756_),
    .Y(_11833_)
);

NAND2X1 _12354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg_9_bF$buf2),
    .Y(_7228_)
);

OR2X2 _22872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1191_),
    .Y(_1197_)
);

INVX1 _22452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_736_),
    .Y(_737_)
);

AOI21X1 _22032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .B(_262_),
    .C(_259_),
    .Y(_277_)
);

NAND2X1 _13979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf5),
    .B(areg_12_bF$buf0),
    .Y(_3359_)
);

OAI21X1 _13559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2898_),
    .B(_2897_),
    .C(_2896_),
    .Y(_2899_)
);

OAI21X1 _13139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2437_),
    .B(_2438_),
    .C(_2439_),
    .Y(_2440_)
);

NOR2X1 _23657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2051_),
    .B(_2050_),
    .Y(_0_[56])
);

FILL SFILL3720x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _23237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1589_),
    .B(_1577_),
    .Y(_1594_)
);

FILL SFILL43960x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4124_),
    .B(_4122_),
    .C(_4113_),
    .Y(_4389_)
);

AND2X2 _14500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_17_bF$buf1),
    .Y(_3930_)
);

INVX8 _17392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_27_bF$buf4),
    .Y(_7100_)
);

FILL SFILL43880x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48840x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5009_),
    .B(_5099_),
    .C(_5098_),
    .Y(_5250_)
);

OAI21X1 _18597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8400_),
    .B(_8407_),
    .C(_8410_),
    .Y(_8420_)
);

AND2X2 _18177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf5),
    .B(areg_28_bF$buf5),
    .Y(_7960_)
);

FILL FILL74040x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11831_),
    .B(_11838_),
    .C(_11840_),
    .Y(_11847_)
);

NAND3X1 _21303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11378_),
    .B(_11382_),
    .C(_11386_),
    .Y(_11387_)
);

NAND3X1 _14097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3475_),
    .B(_3479_),
    .C(_3483_),
    .Y(_3489_)
);

FILL SFILL33880x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(_1256_),
    .C(_1254_),
    .Y(_1257_)
);

NAND2X1 _22508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_797_),
    .Y(_798_)
);

FILL SFILL49080x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _16663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_25_bF$buf0),
    .Y(_6300_)
);

NAND2X1 _16243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_14_bF$buf3),
    .Y(_5840_)
);

FILL SFILL49000x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7604_),
    .B(_7610_),
    .C(_7613_),
    .Y(_7620_)
);

NAND3X1 _17448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7141_),
    .B(_7148_),
    .C(_7151_),
    .Y(_7161_)
);

AOI22X1 _17028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf0),
    .B(areg_29_bF$buf5),
    .C(breg_1_bF$buf4),
    .D(areg_28_bF$buf3),
    .Y(_6700_)
);

NAND3X1 _12583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9598_),
    .B(_9631_),
    .C(_9663_),
    .Y(_9740_)
);

NOR2X1 _12163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_3646__bF$buf1),
    .Y(_5135_)
);

NOR2X1 _22681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf3),
    .B(_5676_),
    .Y(_988_)
);

FILL SFILL23880x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _22261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_514_),
    .B(_519_),
    .C(_508_),
    .Y(_528_)
);

NAND2X1 _13788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3147_),
    .B(_3144_),
    .Y(_3151_)
);

NOR3X1 _13368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_2690_),
    .C(_2686_),
    .Y(_2691_)
);

BUFX2 _23886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[4]),
    .Y(y[4])
);

NOR3X1 _23466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1843_),
    .B(_1745_),
    .C(_1842_),
    .Y(_1844_)
);

NAND3X1 _23046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1381_),
    .B(_1382_),
    .C(_1385_),
    .Y(_1386_)
);

FILL SFILL8840x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .B(_5490_),
    .C(_5471_),
    .Y(_5501_)
);

NOR2X1 _15514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5034_),
    .B(_5039_),
    .Y(_5040_)
);

NAND3X1 _16719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6342_),
    .B(_6348_),
    .C(_6351_),
    .Y(_6361_)
);

AOI21X1 _21952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_189_),
    .B(_187_),
    .C(_93_),
    .Y(_190_)
);

AOI21X1 _21532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11331_),
    .B(_11354_),
    .C(_11352_),
    .Y(_11638_)
);

OAI21X1 _21112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf3),
    .B(_6300__bF$buf3),
    .C(_11173_),
    .Y(_11178_)
);

AOI21X1 _12639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8720_),
    .B(_8906_),
    .C(_8884_),
    .Y(_10353_)
);

NOR3X1 _12219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5716_),
    .B(_5727_),
    .C(_5738_),
    .Y(_5749_)
);

OR2X2 _22737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1043_),
    .B(_1048_),
    .Y(_1049_)
);

AOI21X1 _22317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_583_),
    .B(_581_),
    .C(_580_),
    .Y(_589_)
);

FILL SFILL43960x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6550_),
    .Y(_6551_)
);

NAND3X1 _16472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6081_),
    .B(_6085_),
    .C(_6089_),
    .Y(_6090_)
);

NOR3X1 _16052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5623_),
    .B(_5624_),
    .C(_5622_),
    .Y(_5631_)
);

FILL SFILL64040x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL19000x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7409_),
    .B(_7410_),
    .C(_7402_),
    .Y(_7411_)
);

AOI21X1 _17257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6946_),
    .B(_6950_),
    .C(_6931_),
    .Y(_6951_)
);

AOI21X1 _12392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6472_),
    .B(_6593_),
    .C(_6527_),
    .Y(_7645_)
);

NOR2X1 _22490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_777_),
    .Y(_778_)
);

OAI21X1 _22070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_314_),
    .C(_317_),
    .Y(_318_)
);

NOR2X1 _20803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10831_),
    .B(_10838_),
    .Y(_10839_)
);

NAND2X1 _13597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .B(_2789_),
    .Y(_2942_)
);

OAI21X1 _13177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2472_),
    .B(_2471_),
    .C(_2458_),
    .Y(_2482_)
);

OR2X2 _23695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2083_),
    .B(_2092_),
    .Y(_2093_)
);

AOI21X1 _23275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .B(_1509_),
    .C(_1518_),
    .Y(_1636_)
);

OAI21X1 _19823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9410_),
    .B(_9401_),
    .C(_9405_),
    .Y(_9765_)
);

OAI21X1 _19403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9299_),
    .B(_9300_),
    .C(_9298_),
    .Y(_9304_)
);

NAND3X1 _15743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5284_),
    .B(_5291_),
    .C(_4964_),
    .Y(_5292_)
);

NAND2X1 _15323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4238_),
    .B(_4831_),
    .Y(_4832_)
);

INVX2 _16948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6611_),
    .Y(_6612_)
);

AOI21X1 _16528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5761_),
    .B(_5763_),
    .C(_5769_),
    .Y(_6151_)
);

INVX1 _16108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5677_),
    .Y(_5691_)
);

OAI21X1 _21761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11715_),
    .B(_11827_),
    .C(_11837_),
    .Y(_11888_)
);

AOI21X1 _21341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11411_),
    .B(_11418_),
    .C(_11368_),
    .Y(_11429_)
);

FILL SFILL8920x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(_943_),
    .C(_921_),
    .Y(_954_)
);

FILL SFILL23800x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8194_),
    .B(_8172_),
    .C(_8128_),
    .Y(_8260_)
);

OAI21X1 _22966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_989_),
    .B(_1139_),
    .C(_1146_),
    .Y(_1299_)
);

OAI21X1 _12028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf2),
    .B(_3646__bF$buf1),
    .C(_2814_),
    .Y(_3657_)
);

NOR2X1 _22546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5369_),
    .B(_5921__bF$buf3),
    .Y(_840_)
);

OAI21X1 _22126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_7100__bF$buf0),
    .C(_379_),
    .Y(_380_)
);

FILL SFILL8840x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5866_),
    .B(_5871_),
    .C(_5872_),
    .Y(_5882_)
);

FILL SFILL13880x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7197_),
    .B(_7201_),
    .C(_6810_),
    .Y(_7202_)
);

NAND3X1 _17066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6735_),
    .B(_6741_),
    .C(_6648_),
    .Y(_6742_)
);

FILL SFILL74120x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13800x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10622_),
    .B(_10629_),
    .C(_10348_),
    .Y(_10630_)
);

NOR2X1 _23084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .B(_1426_),
    .Y(_1427_)
);

INVX1 _19632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9173_),
    .Y(_9556_)
);

OAI21X1 _19212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9093_),
    .B(_9091_),
    .C(_9090_),
    .Y(_9094_)
);

OAI22X1 _21817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11661_),
    .B(_40_),
    .C(_11724_),
    .D(_11719_),
    .Y(_41_)
);

NAND2X1 _15972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf2),
    .B(areg_21_bF$buf2),
    .Y(_5543_)
);

NOR3X1 _15552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5018_),
    .B(_5024_),
    .C(_5029_),
    .Y(_5082_)
);

AOI21X1 _15132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4606_),
    .B(_4612_),
    .C(_4359_),
    .Y(_4623_)
);

OAI21X1 _16757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6401_),
    .B(_6402_),
    .C(_6400_),
    .Y(_6403_)
);

NAND2X1 _16337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5564_),
    .B(_5932_),
    .Y(_5943_)
);

NAND3X1 _21990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11881_),
    .B(_226_),
    .C(_227_),
    .Y(_231_)
);

NAND3X1 _21570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11671_),
    .B(_11675_),
    .C(_11677_),
    .Y(_11678_)
);

AOI21X1 _21150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11213_),
    .B(_11218_),
    .C(_11133_),
    .Y(_11219_)
);

AND2X2 _12677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10737_),
    .B(_10748_),
    .Y(_10770_)
);

OAI21X1 _12257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5530_),
    .B(_6143_),
    .C(_6154_),
    .Y(_6165_)
);

OR2X2 _22775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1087_),
    .B(_1085_),
    .Y(_1091_)
);

NAND2X1 _22355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_628_),
    .Y(_631_)
);

NAND3X1 _18903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8750_),
    .B(_8754_),
    .C(_8755_),
    .Y(_8756_)
);

OAI21X1 _16090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5670_),
    .B(_4979_),
    .C(_5345_),
    .Y(_5671_)
);

AOI21X1 _14823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4278_),
    .B(_4277_),
    .C(_4276_),
    .Y(_4284_)
);

INVX2 _14403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3823_),
    .Y(_3824_)
);

OAI21X1 _17295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6979_),
    .B(_6980_),
    .C(_6976_),
    .Y(_6993_)
);

AND2X2 _15608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4793_),
    .B(_4788_),
    .Y(_5143_)
);

OAI21X1 _20841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10878_),
    .B(_10879_),
    .C(_10877_),
    .Y(_10881_)
);

NAND3X1 _20421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10415_),
    .B(_10401_),
    .C(_10405_),
    .Y(_10420_)
);

NAND3X1 _20001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9957_),
    .B(_9958_),
    .C(_9956_),
    .Y(_9960_)
);

FILL SFILL44040x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9511_),
    .B(_9805_),
    .C(_9804_),
    .Y(_9807_)
);

OAI21X1 _19441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9338_),
    .B(_9337_),
    .C(_9335_),
    .Y(_9346_)
);

AOI21X1 _19021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8849_),
    .B(_8850_),
    .C(_8482_),
    .Y(_8885_)
);

FILL SFILL8920x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _11948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2584_),
    .C(_2770_),
    .Y(_2781_)
);

OAI21X1 _21626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11735_),
    .B(_11739_),
    .C(_11727_),
    .Y(_11740_)
);

NOR2X1 _21206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11259_),
    .B(_11262_),
    .Y(_11281_)
);

INVX1 _15781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4974_),
    .Y(_5333_)
);

XNOR2X1 _15361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4852_),
    .B(_4872_),
    .Y(_4874_)
);

NOR2X1 _16986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf3),
    .B(_3961__bF$buf2),
    .Y(_6653_)
);

AOI21X1 _16566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5782_),
    .B(_5803_),
    .C(_5807_),
    .Y(_6193_)
);

AOI21X1 _16146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5728_),
    .B(_5729_),
    .C(_5726_),
    .Y(_5733_)
);

NAND2X1 _12486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8643_),
    .B(_8665_),
    .Y(_8676_)
);

OAI21X1 _12066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3876_),
    .B(_3471_),
    .C(_4061_),
    .Y(_4072_)
);

NAND3X1 _22584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_835_),
    .C(_837_),
    .Y(_882_)
);

OAI21X1 _22164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_416_),
    .C(_401_),
    .Y(_422_)
);

AOI21X1 _18712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8539_),
    .B(_8538_),
    .C(_8537_),
    .Y(_8546_)
);

FILL SFILL59160x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2169_),
    .B(_2193_),
    .Y(_2194_)
);

AOI21X1 _23369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1731_),
    .B(_1730_),
    .C(_1728_),
    .Y(_1738_)
);

FILL SFILL64120x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_27_bF$buf3),
    .Y(_9868_)
);

INVX1 _14632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4073_),
    .Y(_4074_)
);

AND2X2 _14212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3604_),
    .B(_3602_),
    .Y(_3615_)
);

AOI21X1 _15837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5026_),
    .B(_5028_),
    .C(_5022_),
    .Y(_5394_)
);

NAND3X1 _15417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4925_),
    .B(_4915_),
    .C(_4922_),
    .Y(_4935_)
);

AOI21X1 _20650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9260_),
    .B(_8878_),
    .C(_10669_),
    .Y(_10670_)
);

NAND3X1 _20230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9908_),
    .B(_9910_),
    .C(_9902_),
    .Y(_10210_)
);

AOI21X1 _19670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9595_),
    .B(_9596_),
    .C(_9594_),
    .Y(_9597_)
);

AND2X2 _19250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8730_),
    .B(_8725_),
    .Y(_9136_)
);

FILL SFILL54120x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_77_),
    .C(_76_),
    .Y(_83_)
);

OAI21X1 _21435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10565_),
    .B(_11237_),
    .C(_11531_),
    .Y(_11532_)
);

NAND3X1 _21015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11068_),
    .B(_11070_),
    .C(_11069_),
    .Y(_11071_)
);

FILL SFILL54040x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf2),
    .B(_2465__bF$buf4),
    .C(_5114_),
    .Y(_5123_)
);

NOR2X1 _15170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4659_),
    .B(_4661_),
    .Y(_4663_)
);

NOR2X1 _13903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3261_),
    .B(_3264_),
    .Y(_3277_)
);

NAND2X1 _16795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf2),
    .B(breg_26_bF$buf0),
    .Y(_6444_)
);

AOI21X1 _16375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5511_),
    .B(_5598_),
    .C(_5983_),
    .Y(_5984_)
);

FILL SFILL44040x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _12295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf4),
    .Y(_6582_)
);

FILL SFILL54040x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _22393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_439_),
    .B(_667_),
    .Y(_672_)
);

NAND2X1 _18941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8796_),
    .B(_8795_),
    .Y(_8798_)
);

AND2X2 _18521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf3),
    .B(areg_26_bF$buf3),
    .Y(_8338_)
);

OAI21X1 _18101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7875_),
    .B(_7874_),
    .C(_7873_),
    .Y(_7877_)
);

AOI21X1 _20706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10727_),
    .B(_10728_),
    .C(_10702_),
    .Y(_10732_)
);

INVX1 _23598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .Y(_1987_)
);

NOR3X1 _23178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1528_),
    .C(_1529_),
    .Y(_1530_)
);

OAI22X1 _19726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6582__bF$buf1),
    .B(_6050__bF$buf1),
    .C(_7711__bF$buf3),
    .D(_5668__bF$buf4),
    .Y(_9658_)
);

AOI21X1 _19306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8800_),
    .B(_8798_),
    .C(_8821_),
    .Y(_9198_)
);

OAI21X1 _14861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4323_),
    .B(_4324_),
    .C(_4322_),
    .Y(_4326_)
);

FILL SFILL69240x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3860_),
    .B(_3864_),
    .Y(_3866_)
);

NAND3X1 _14021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3398_),
    .B(_3404_),
    .C(_3401_),
    .Y(_3406_)
);

FILL SFILL69160x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _15646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5183_),
    .B(_5184_),
    .Y(_5185_)
);

OAI22X1 _15226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4159_),
    .B(_4723_),
    .C(_4724_),
    .D(_4449_),
    .Y(_4725_)
);

XNOR2X1 _11986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2497_),
    .B(_2616_),
    .Y(_3198_)
);

NOR3X1 _21664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11775_),
    .B(_11777_),
    .C(_11774_),
    .Y(_11782_)
);

OAI21X1 _21244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11321_),
    .B(_11012_),
    .C(_11287_),
    .Y(_11322_)
);

FILL SFILL28760x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3720x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1038_),
    .B(_1192_),
    .Y(_1193_)
);

FILL SFILL3640x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _22449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf3),
    .B(_7225__bF$buf0),
    .Y(_733_)
);

OAI21X1 _22029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2884__bF$buf2),
    .B(_6050__bF$buf3),
    .C(_261_),
    .Y(_273_)
);

INVX1 _13712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3061_),
    .Y(_3068_)
);

INVX1 _23810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .Y(_2216_)
);

XNOR2X1 _16184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5751_),
    .B(_5747_),
    .Y(_5775_)
);

FILL FILL74120x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4385_),
    .B(_4367_),
    .Y(_4386_)
);

FILL SFILL28680x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_26_bF$buf1),
    .Y(_7096_)
);

FILL SFILL49160x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8586_),
    .B(_8585_),
    .C(_8581_),
    .Y(_8587_)
);

NAND2X1 _18330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf2),
    .B(breg_24_bF$buf3),
    .Y(_8127_)
);

FILL SFILL54120x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10638_),
    .B(_10345_),
    .C(_10645_),
    .Y(_10984_)
);

AOI21X1 _20515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9797_),
    .B(_10502_),
    .C(_10161_),
    .Y(_10523_)
);

XNOR2X1 _19955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9901_),
    .B(_9905_),
    .Y(_9909_)
);

OAI21X1 _19535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9443_),
    .B(_9445_),
    .C(_9448_),
    .Y(_9449_)
);

NAND3X1 _19115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8974_),
    .B(_8978_),
    .C(_8980_),
    .Y(_8988_)
);

OAI21X1 _14670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3646__bF$buf3),
    .B(_2560__bF$buf4),
    .C(_4102_),
    .Y(_4115_)
);

AOI21X1 _14250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3647_),
    .B(_3645_),
    .C(_3642_),
    .Y(_3656_)
);

FILL SFILL59320x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33640x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5405_),
    .B(_5430_),
    .C(_5435_),
    .Y(_5436_)
);

FILL SFILL39160x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _15455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg_24_bF$buf1),
    .C(areg[0]),
    .D(breg_25_bF$buf0),
    .Y(_4975_)
);

AOI21X1 _15035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4509_),
    .B(_4510_),
    .C(_4508_),
    .Y(_4516_)
);

AOI21X1 _21893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_124_),
    .C(_121_),
    .Y(_125_)
);

NAND3X1 _21473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11323_),
    .B(_11567_),
    .C(_11568_),
    .Y(_11574_)
);

OAI21X1 _21053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11107_),
    .B(_11108_),
    .C(_11058_),
    .Y(_11113_)
);

OAI21X1 _17601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7326_),
    .B(_6924_),
    .C(_7004_),
    .Y(_7328_)
);

NAND2X1 _22678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf0),
    .B(breg_25_bF$buf1),
    .Y(_984_)
);

NOR3X1 _22258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_521_),
    .C(_523_),
    .Y(_524_)
);

NAND3X1 _18806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8639_),
    .B(_8647_),
    .C(_8648_),
    .Y(_8649_)
);

FILL SFILL69240x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _13941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3316_),
    .B(_3317_),
    .Y(_3319_)
);

NOR2X1 _13521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2857_),
    .B(_2851_),
    .Y(_2859_)
);

INVX1 _13101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .Y(_2399_)
);

OAI21X1 _14726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7217__bF$buf2),
    .B(_10869__bF$buf2),
    .C(_4167_),
    .Y(_4177_)
);

NAND3X1 _14306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3706_),
    .B(_3666_),
    .C(_3700_),
    .Y(_3718_)
);

AOI21X1 _17198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6543_),
    .B(_6541_),
    .C(_6885_),
    .Y(_6886_)
);

FILL SFILL69160x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69080x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8520x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10766_),
    .B(_10771_),
    .C(_10773_),
    .Y(_10774_)
);

AOI21X1 _20324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10307_),
    .B(_10308_),
    .C(_10306_),
    .Y(_10314_)
);

OAI21X1 _19764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549__bF$buf2),
    .B(_5315__bF$buf4),
    .C(_9692_),
    .Y(_9700_)
);

AOI21X1 _19344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8479_),
    .B(_8856_),
    .C(_9239_),
    .Y(_9240_)
);

FILL SFILL28760x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_181_),
    .B(_185_),
    .Y(_186_)
);

NAND3X1 _21529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11619_),
    .B(_11610_),
    .C(_11623_),
    .Y(_11634_)
);

NAND2X1 _21109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11172_),
    .B(_11173_),
    .Y(_11174_)
);

FILL SFILL3800x50 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5211_),
    .B(_5216_),
    .C(_5219_),
    .Y(_5226_)
);

AOI21X1 _15264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4570_),
    .B(_4576_),
    .C(_4497_),
    .Y(_4767_)
);

FILL FILL74120x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _16889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf3),
    .B(breg_16_bF$buf4),
    .Y(_6547_)
);

NAND3X1 _16469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6083_),
    .B(_6084_),
    .C(_6082_),
    .Y(_6085_)
);

NAND3X1 _16049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5361_),
    .B(_5359_),
    .C(_5356_),
    .Y(_5627_)
);

OAI21X1 _21282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11363_),
    .B(_11357_),
    .C(_11328_),
    .Y(_11364_)
);

FILL SFILL18760x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7570_),
    .B(_7571_),
    .C(_7485_),
    .Y(_7579_)
);

NAND3X1 _17410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7107_),
    .B(_7118_),
    .C(_7115_),
    .Y(_7119_)
);

FILL SFILL33960x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf0),
    .B(areg_7_bF$buf1),
    .C(breg_4_bF$buf5),
    .D(areg_6_bF$buf4),
    .Y(_7623_)
);

NAND2X1 _22487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_21_bF$buf4),
    .B(breg_26_bF$buf0),
    .Y(_775_)
);

NOR3X1 _22067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_301_),
    .C(_304_),
    .Y(_315_)
);

NAND3X1 _18615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8433_),
    .B(_8434_),
    .C(_8432_),
    .Y(_8440_)
);

NAND3X1 _13750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3100_),
    .B(_3107_),
    .C(_3108_),
    .Y(_3109_)
);

NAND3X1 _13330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2646_),
    .B(_2648_),
    .C(_2647_),
    .Y(_2649_)
);

FILL SFILL39160x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4387_),
    .B(_4386_),
    .Y(_4428_)
);

OAI21X1 _14535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3963_),
    .B(_3968_),
    .C(_3956_),
    .Y(_3969_)
);

NAND3X1 _14115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3507_),
    .B(_2537_),
    .C(_1271_),
    .Y(_3508_)
);

FILL SFILL23960x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf2),
    .B(breg_28_bF$buf4),
    .Y(_11025_)
);

AND2X2 _20553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf2),
    .B(areg_30_bF$buf2),
    .Y(_10565_)
);

NAND2X1 _20133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9728_),
    .B(_9736_),
    .Y(_10104_)
);

NAND3X1 _19993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9941_),
    .B(_9944_),
    .C(_9756_),
    .Y(_9951_)
);

INVX2 _19573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9490_),
    .Y(_9491_)
);

NOR3X1 _19153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9015_),
    .B(_9024_),
    .C(_9025_),
    .Y(_9030_)
);

FILL SFILL69320x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11883_),
    .B(_11601_),
    .C(_11846_),
    .Y(_11884_)
);

OAI21X1 _21338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11424_),
    .B(_11133_),
    .C(_11222_),
    .Y(_11425_)
);

AOI22X1 _12601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9883_),
    .B(_8402_),
    .C(_9904_),
    .D(_9926_),
    .Y(_9937_)
);

XNOR2X1 _15493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5016_),
    .B(_5011_),
    .Y(_5017_)
);

NAND3X1 _15073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4535_),
    .B(_4557_),
    .C(_4549_),
    .Y(_4558_)
);

AOI21X1 _13806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2893_),
    .B(_2875_),
    .C(_2897_),
    .Y(_3171_)
);

BUFX2 _23904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[22]),
    .Y(y[22])
);

AOI21X1 _16698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6333_),
    .B(_6332_),
    .C(_6331_),
    .Y(_6338_)
);

OAI21X1 _16278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5877_),
    .B(_5873_),
    .C(_5839_),
    .Y(_5878_)
);

NAND2X1 _21091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_19_bF$buf4),
    .B(areg_23_bF$buf3),
    .Y(_11155_)
);

FILL SFILL59240x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376__bF$buf3),
    .B(_5420__bF$buf1),
    .C(_5475_),
    .Y(_5519_)
);

OAI21X1 _22296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_564_),
    .B(_565_),
    .C(_557_),
    .Y(_566_)
);

OAI21X1 _18844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8690_),
    .B(_8689_),
    .C(_8688_),
    .Y(_8691_)
);

OAI22X1 _18424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362__bF$buf2),
    .B(_3146__bF$buf1),
    .C(_2560__bF$buf0),
    .D(_2884__bF$buf3),
    .Y(_8231_)
);

AOI21X1 _18004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7759_),
    .B(_7750_),
    .C(_7706_),
    .Y(_7770_)
);

NAND3X1 _20609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10619_),
    .B(_10620_),
    .C(_10461_),
    .Y(_10626_)
);

FILL FILL74200x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9547_),
    .B(_9546_),
    .C(_9531_),
    .Y(_9552_)
);

INVX2 _19209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9006_),
    .Y(_9090_)
);

AND2X2 _14764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf3),
    .B(areg_18_bF$buf4),
    .Y(_4219_)
);

OAI21X1 _14344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3758_),
    .B(_3759_),
    .C(_3521_),
    .Y(_3760_)
);

DFFPOSX1 _24022_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[12]),
    .CLK(clk_bF$buf1),
    .D(a[12])
);

FILL SFILL49240x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5538_),
    .B(_5534_),
    .Y(_5539_)
);

OAI21X1 _15549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5076_),
    .B(_5077_),
    .C(_5073_),
    .Y(_5078_)
);

NOR3X1 _15129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4312_),
    .B(_4313_),
    .C(_4311_),
    .Y(_4619_)
);

NAND2X1 _20782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf5),
    .B(breg_23_bF$buf3),
    .Y(_10816_)
);

INVX2 _20362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10354_),
    .Y(_10355_)
);

OAI21X1 _16910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6565_),
    .B(_6566_),
    .C(_6569_),
    .Y(_6570_)
);

OAI21X1 _19382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8911_),
    .B(_8897_),
    .C(_8921_),
    .Y(_9281_)
);

FILL SFILL33960x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_226_),
    .B(_227_),
    .C(_11881_),
    .Y(_228_)
);

NAND3X1 _21567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11672_),
    .B(_11673_),
    .C(_11674_),
    .Y(_11675_)
);

AOI21X1 _21147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10932_),
    .B(_10938_),
    .C(_10258_),
    .Y(_11216_)
);

OR2X2 _12830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_527_),
    .Y(_538_)
);

NOR3X1 _12410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7799_),
    .B(_7645_),
    .C(_7788_),
    .Y(_7843_)
);

AOI21X1 _13615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2947_),
    .B(_2952_),
    .C(_2757_),
    .Y(_2962_)
);

NAND2X1 _23713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1948_),
    .B(_1989_),
    .Y(_2112_)
);

INVX8 _16087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_27_bF$buf0),
    .Y(_5668_)
);

FILL SFILL23960x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8426_),
    .B(_8427_),
    .C(_8187_),
    .Y(_8481_)
);

AOI21X1 _18233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7434_),
    .B(_7588_),
    .C(_8020_),
    .Y(_8021_)
);

FILL SFILL69320x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10149_),
    .B(_10855_),
    .C(_10515_),
    .Y(_10877_)
);

OAI21X1 _20418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10412_),
    .B(_10411_),
    .C(_10415_),
    .Y(_10416_)
);

NAND3X1 _19858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9794_),
    .B(_9801_),
    .C(_9802_),
    .Y(_9803_)
);

NAND3X1 _19438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9321_),
    .B(_9341_),
    .C(_9336_),
    .Y(_9342_)
);

OAI21X1 _19018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8880_),
    .B(_8475_),
    .C(_8866_),
    .Y(_8881_)
);

AOI21X1 _14993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4165_),
    .B(_4169_),
    .C(_4172_),
    .Y(_4469_)
);

AOI21X1 _14573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4009_),
    .B(_4010_),
    .C(_4007_),
    .Y(_4011_)
);

OAI21X1 _14153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf2),
    .B(_2586__bF$buf0),
    .C(_3314_),
    .Y(_3550_)
);

AOI21X1 _15778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5011_),
    .B(_5328_),
    .C(_5013_),
    .Y(_5329_)
);

OAI21X1 _15358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4869_),
    .B(_4868_),
    .C(_4867_),
    .Y(_4870_)
);

NAND3X1 _20591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10604_),
    .B(_10605_),
    .C(_10603_),
    .Y(_10607_)
);

NAND2X1 _20171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf1),
    .B(areg_21_bF$buf3),
    .Y(_10146_)
);

AOI21X1 _19191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8662_),
    .B(_8664_),
    .C(_8670_),
    .Y(_9072_)
);

NOR3X1 _21796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_15_),
    .B(_16_),
    .C(_17_),
    .Y(_18_)
);

XNOR2X1 _21376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11444_),
    .B(_11466_),
    .Y(_11467_)
);

NOR2X1 _17924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7674_),
    .B(_7675_),
    .Y(_7682_)
);

NAND2X1 _17504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6908_),
    .B(_7184_),
    .Y(_7221_)
);

AND2X2 _18709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8191_),
    .B(_8192_),
    .Y(_8542_)
);

NOR3X1 _13844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2938_),
    .B(_2939_),
    .C(_2937_),
    .Y(_3213_)
);

AOI21X1 _13424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2741_),
    .B(_2742_),
    .C(_2527_),
    .Y(_2752_)
);

BUFX2 _23942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[60]),
    .Y(y[60])
);

NAND3X1 _13004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2293_),
    .C(_2298_),
    .Y(_2299_)
);

NAND2X1 _23522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_25_bF$buf4),
    .B(areg_31_bF$buf4),
    .Y(_1904_)
);

NOR2X1 _23102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6300__bF$buf2),
    .B(_5676_),
    .Y(_1447_)
);

OAI22X1 _14629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_3781__bF$buf0),
    .C(_2376__bF$buf2),
    .D(_4069_),
    .Y(_4070_)
);

AOI21X1 _14209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3609_),
    .B(_3608_),
    .C(_3607_),
    .Y(_3610_)
);

OAI21X1 _18882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8357_),
    .B(_8355_),
    .C(_8349_),
    .Y(_8733_)
);

NAND3X1 _18462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8269_),
    .B(_8270_),
    .C(_8272_),
    .Y(_8273_)
);

XNOR2X1 _18042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7790_),
    .B(_7784_),
    .Y(_7812_)
);

NOR3X1 _20647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9244_),
    .B(_8881_),
    .C(_9248_),
    .Y(_10667_)
);

NAND2X1 _20227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9921_),
    .B(_9920_),
    .Y(_10207_)
);

INVX8 _11910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_3_bF$buf4),
    .Y(_2365_)
);

NAND2X1 _19667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9593_),
    .B(_9592_),
    .Y(_9594_)
);

OAI21X1 _19247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8768_),
    .B(_8744_),
    .C(_8756_),
    .Y(_9133_)
);

FILL SFILL23640x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _14382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3785_),
    .B(_3800_),
    .Y(_3801_)
);

DFFPOSX1 _24060_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[18]),
    .CLK(clk_bF$buf5),
    .D(b[18])
);

FILL SFILL8680x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5118_),
    .B(_5119_),
    .C(_5110_),
    .Y(_5120_)
);

NAND3X1 _15167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_23_bF$buf3),
    .C(_4365_),
    .Y(_4660_)
);

FILL SFILL8600x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13640x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11257_),
    .B(_11255_),
    .C(_11256_),
    .Y(_11258_)
);

AOI21X1 _17733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7467_),
    .B(_7468_),
    .C(_7466_),
    .Y(_7473_)
);

NAND3X1 _17313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6923_),
    .B(_7010_),
    .C(_7011_),
    .Y(_7012_)
);

FILL SFILL74280x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8790_),
    .B(_8793_),
    .C(_8740_),
    .Y(_8794_)
);

OAI21X1 _18518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7929_),
    .B(_8333_),
    .C(_7938_),
    .Y(_8334_)
);

AOI21X1 _13653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2795_),
    .B(_2798_),
    .C(_3002_),
    .Y(_3003_)
);

OAI21X1 _13233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2542_),
    .B(_2541_),
    .C(_2355_),
    .Y(_2543_)
);

XNOR2X1 _23751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2152_),
    .B(_2125_),
    .Y(_2154_)
);

NAND2X1 _23331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1577_),
    .B(_1589_),
    .Y(_1697_)
);

FILL SFILL74200x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4032_),
    .B(_4034_),
    .C(_4025_),
    .Y(_4322_)
);

NAND3X1 _14438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3852_),
    .B(_3858_),
    .C(_3848_),
    .Y(_3862_)
);

INVX8 _14018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_19_bF$buf2),
    .Y(_3402_)
);

FILL SFILL64200x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8486_),
    .B(_8514_),
    .C(_8510_),
    .Y(_8523_)
);

AOI21X1 _18271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8048_),
    .B(_8051_),
    .C(_7659_),
    .Y(_8064_)
);

FILL SFILL64280x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _20876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf1),
    .B(areg_31_bF$buf3),
    .Y(_10919_)
);

OAI21X1 _20456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10451_),
    .B(_10450_),
    .C(_10448_),
    .Y(_10458_)
);

AOI21X1 _20036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9941_),
    .B(_9944_),
    .C(_9756_),
    .Y(_9997_)
);

AOI21X1 _19896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9509_),
    .B(_9515_),
    .C(_9516_),
    .Y(_9845_)
);

NAND3X1 _19476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9374_),
    .B(_9380_),
    .C(_9370_),
    .Y(_9384_)
);

AOI21X1 _19056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8922_),
    .B(_8919_),
    .C(_8894_),
    .Y(_8923_)
);

AOI21X1 _14191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3357_),
    .B(_3442_),
    .C(_3447_),
    .Y(_3592_)
);

INVX2 _12924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .Y(_1565_)
);

AOI21X1 _12504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7569_),
    .B(_7624_),
    .C(_7602_),
    .Y(_8874_)
);

NAND3X1 _22602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_891_),
    .C(_887_),
    .Y(_902_)
);

FILL SFILL54200x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4910_),
    .B(_4911_),
    .C(_4902_),
    .Y(_4912_)
);

AND2X2 _13709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2807_),
    .B(_3062_),
    .Y(_3064_)
);

OAI21X1 _23807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2115_),
    .B(_2209_),
    .C(_2212_),
    .Y(_2213_)
);

BUFX2 BUFX2_insert210 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[26]),
    .Y(areg_26_bF$buf2)
);

BUFX2 BUFX2_insert211 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[26]),
    .Y(areg_26_bF$buf1)
);

BUFX2 BUFX2_insert212 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[26]),
    .Y(areg_26_bF$buf0)
);

BUFX2 BUFX2_insert213 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf4)
);

BUFX2 BUFX2_insert214 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf3)
);

NAND3X1 _17962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7716_),
    .B(_7720_),
    .C(_7723_),
    .Y(_7724_)
);

AOI21X1 _17542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7256_),
    .B(_7257_),
    .C(_7232_),
    .Y(_7263_)
);

BUFX2 BUFX2_insert215 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf2)
);

BUFX2 BUFX2_insert216 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf1)
);

XNOR2X1 _17122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6418_),
    .B(_6803_),
    .Y(_0_[29])
);

BUFX2 BUFX2_insert217 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf0)
);

BUFX2 BUFX2_insert218 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[23]),
    .Y(areg_23_bF$buf4)
);

BUFX2 BUFX2_insert219 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[23]),
    .Y(areg_23_bF$buf3)
);

FILL SFILL74040x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_459_),
    .B(_450_),
    .C(_248_),
    .Y(_460_)
);

NAND3X1 _18747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8567_),
    .B(_8571_),
    .C(_8574_),
    .Y(_8584_)
);

OAI21X1 _18327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7715_),
    .B(_7712_),
    .C(_7718_),
    .Y(_8124_)
);

FILL SFILL23640x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg_18_bF$buf5),
    .Y(_3254_)
);

DFFPOSX1 _23980_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[34]),
    .CLK(clk_bF$buf3),
    .D(_0_[34])
);

AOI21X1 _13462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2594_),
    .B(_2599_),
    .C(_2613_),
    .Y(_2794_)
);

AND2X2 _13042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_965_),
    .Y(_2337_)
);

NAND3X1 _23560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_1930_),
    .C(_1937_),
    .Y(_1946_)
);

OAI21X1 _23140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1487_),
    .B(_1486_),
    .C(_1362_),
    .Y(_1488_)
);

FILL SFILL8680x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _14667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4111_),
    .Y(_4112_)
);

OAI22X1 _14247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3130_),
    .B(_3390_),
    .C(_3388_),
    .D(_3392_),
    .Y(_3653_)
);

FILL SFILL8600x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44120x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7851_),
    .B(_7852_),
    .C(_7819_),
    .Y(_7853_)
);

AND2X2 _20685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf0),
    .B(breg_27_bF$buf5),
    .Y(_10709_)
);

OAI21X1 _20265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10247_),
    .B(_10248_),
    .C(_10246_),
    .Y(_10249_)
);

AOI21X1 _16813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6133_),
    .B(_6463_),
    .C(_6462_),
    .Y(_6464_)
);

OAI21X1 _19285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8369_),
    .B(_9173_),
    .C(_9174_),
    .Y(_9175_)
);

FILL SFILL44040x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _12733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11350_),
    .B(_11329_),
    .C(_11318_),
    .Y(_11384_)
);

NAND3X1 _12313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6703_),
    .B(_6769_),
    .C(_6341_),
    .Y(_6780_)
);

XOR2X1 _22831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1137_),
    .Y(_1152_)
);

NOR2X1 _22411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_690_),
    .B(_676_),
    .Y(_693_)
);

FILL SFILL38840x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43800x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _13938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .B(breg_12_bF$buf3),
    .Y(_3315_)
);

INVX2 _13518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2854_),
    .Y(_2855_)
);

NOR2X1 _23616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6686__bF$buf1),
    .B(_6815__bF$buf3),
    .Y(_2007_)
);

FILL SFILL64200x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf3),
    .B(areg_26_bF$buf1),
    .Y(_7515_)
);

AOI21X1 _17351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6652_),
    .B(_6674_),
    .C(_6671_),
    .Y(_7055_)
);

NAND3X1 _18976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8829_),
    .B(_8831_),
    .C(_8828_),
    .Y(_8836_)
);

FILL SFILL33800x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8365_),
    .B(_8366_),
    .C(_8362_),
    .Y(_8376_)
);

OAI21X1 _18136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7908_),
    .B(_7913_),
    .C(_7914_),
    .Y(_7915_)
);

OAI21X1 _13691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3038_),
    .B(_3037_),
    .C(_3035_),
    .Y(_3045_)
);

NOR2X1 _13271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2583_),
    .Y(_2585_)
);

FILL SFILL54200x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _14896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_23_bF$buf3),
    .Y(_4363_)
);

NAND3X1 _14476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3886_),
    .B(_3893_),
    .C(_3873_),
    .Y(_3904_)
);

FILL SFILL13800x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3355_),
    .B(_3354_),
    .C(_3311_),
    .Y(_3444_)
);

FILL SFILL58920x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_17_bF$buf4),
    .B(areg_22_bF$buf3),
    .Y(_10500_)
);

NAND3X1 _20074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10003_),
    .B(_10030_),
    .C(_10027_),
    .Y(_10039_)
);

AOI21X1 _16622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5888_),
    .B(_5909_),
    .C(_5906_),
    .Y(_6255_)
);

NAND2X1 _16202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_14_bF$buf1),
    .Y(_5795_)
);

AOI21X1 _19094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8623_),
    .B(_8627_),
    .C(_8608_),
    .Y(_8965_)
);

FILL SFILL23720x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11819_),
    .B(_11818_),
    .Y(_11820_)
);

AOI21X1 _21279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11354_),
    .B(_11355_),
    .C(_11331_),
    .Y(_11359_)
);

OAI21X1 _17827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7473_),
    .B(_7474_),
    .C(_7471_),
    .Y(_7576_)
);

NAND2X1 _17407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf5),
    .B(areg_30_bF$buf0),
    .Y(_7116_)
);

NAND2X1 _12962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf0),
    .B(areg_10_bF$buf4),
    .Y(_1979_)
);

AOI21X1 _12542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9236_),
    .B(_9279_),
    .C(_8950_),
    .Y(_9290_)
);

OAI21X1 _12122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4664_),
    .B(_4675_),
    .C(_4653_),
    .Y(_4686_)
);

OAI21X1 _22640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7651_),
    .B(_924_),
    .C(_941_),
    .Y(_942_)
);

NAND2X1 _22220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_477_),
    .Y(_483_)
);

FILL SFILL48920x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3101_),
    .B(_3105_),
    .C(_3104_),
    .Y(_3106_)
);

NOR2X1 _13327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2627_),
    .B(_2437_),
    .Y(_2646_)
);

XNOR2X1 _23845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2244_),
    .Y(_2254_)
);

XOR2X1 _23425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1792_),
    .B(_1798_),
    .Y(_1799_)
);

INVX1 _23005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1268_),
    .Y(_1341_)
);

AOI21X1 _17580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7288_),
    .B(_7293_),
    .C(_7275_),
    .Y(_7304_)
);

AND2X2 _17160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6843_),
    .B(_6841_),
    .Y(_6844_)
);

NOR2X1 _18785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8614_),
    .B(_8612_),
    .Y(_8626_)
);

OAI21X1 _18365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8164_),
    .B(_8165_),
    .C(_8163_),
    .Y(_8166_)
);

AOI21X1 _13080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2312_),
    .B(_2316_),
    .C(_1902_),
    .Y(_2375_)
);

NOR3X1 _21911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_134_),
    .C(_132_),
    .Y(_145_)
);

AOI21X1 _14285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3694_),
    .B(_3689_),
    .C(_3676_),
    .Y(_3695_)
);

FILL SFILL3880x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6499_),
    .B(_6500_),
    .C(_6501_),
    .Y(_6506_)
);

NAND2X1 _16431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5732_),
    .B(_6004_),
    .Y(_6045_)
);

NAND3X1 _16011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5515_),
    .B(_5536_),
    .C(_5537_),
    .Y(_5586_)
);

FILL SFILL28840x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _21088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11150_),
    .B(_11139_),
    .C(_11146_),
    .Y(_11151_)
);

OAI21X1 _17636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7361_),
    .B(_7365_),
    .C(_7352_),
    .Y(_7366_)
);

NAND3X1 _17216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6903_),
    .B(_6904_),
    .C(_6905_),
    .Y(_6906_)
);

XNOR2X1 _12771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11789_),
    .B(_11756_),
    .Y(_11800_)
);

OAI21X1 _12351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6933_),
    .B(_6088_),
    .C(_6834_),
    .Y(_7196_)
);

NAND3X1 _13976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3353_),
    .B(_3355_),
    .C(_3354_),
    .Y(_3356_)
);

XNOR2X1 _13556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2874_),
    .B(_2895_),
    .Y(_2896_)
);

AND2X2 _13136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2426_),
    .Y(_2437_)
);

XNOR2X1 _23654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2048_),
    .B(_1995_),
    .Y(_2049_)
);

AOI21X1 _23234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1502_),
    .B(_1501_),
    .C(_1353_),
    .Y(_1591_)
);

DFFPOSX1 _24019_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[9]),
    .CLK(clk_bF$buf0),
    .D(a[9])
);

AOI21X1 _15702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5228_),
    .B(_5234_),
    .C(_5148_),
    .Y(_5247_)
);

NAND3X1 _18594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8273_),
    .B(_8275_),
    .C(_8268_),
    .Y(_8417_)
);

OAI21X1 _18174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7956_),
    .B(_7548_),
    .C(_7541_),
    .Y(_7957_)
);

FILL SFILL44200x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10602_),
    .Y(_10812_)
);

INVX1 _20359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10350_),
    .Y(_10351_)
);

NOR2X1 _16907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5842_),
    .B(_6223_),
    .Y(_6567_)
);

NAND3X1 _21720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11842_),
    .B(_11840_),
    .C(_11841_),
    .Y(_11843_)
);

NAND2X1 _21300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_21_bF$buf1),
    .Y(_11383_)
);

OAI21X1 _19799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9733_),
    .B(_9734_),
    .C(_9688_),
    .Y(_9738_)
);

NAND2X1 _19379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8979_),
    .B(_8985_),
    .Y(_9277_)
);

OAI21X1 _14094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3484_),
    .B(_3485_),
    .C(_3483_),
    .Y(_3486_)
);

FILL SFILL69080x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_9104__bF$buf1),
    .Y(_505_)
);

OAI21X1 _12407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7788_),
    .B(_7799_),
    .C(_7645_),
    .Y(_7810_)
);

NAND3X1 _22925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1098_),
    .B(_1247_),
    .C(_1251_),
    .Y(_1254_)
);

NAND3X1 _22505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_774_),
    .B(_788_),
    .C(_794_),
    .Y(_795_)
);

NOR3X1 _15299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4803_),
    .B(_4804_),
    .C(_4802_),
    .Y(_4805_)
);

NAND2X1 _16660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf2),
    .B(areg_24_bF$buf3),
    .Y(_6296_)
);

AOI21X1 _16240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5584_),
    .B(_5591_),
    .C(_5513_),
    .Y(_5836_)
);

FILL SFILL3640x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7221_),
    .B(_7611_),
    .C(_7616_),
    .Y(_7617_)
);

NAND3X1 _17445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7016_),
    .B(_7059_),
    .C(_7060_),
    .Y(_7158_)
);

AND2X2 _17025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf5),
    .B(areg_28_bF$buf3),
    .Y(_6697_)
);

NAND3X1 _12580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9641_),
    .B(_8238_),
    .C(_9696_),
    .Y(_9707_)
);

NOR2X1 _12160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3635_),
    .B(_4390_),
    .Y(_5102_)
);

OAI21X1 _13785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf0),
    .B(_3146__bF$buf3),
    .C(_3147_),
    .Y(_3148_)
);

NAND3X1 _13365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2660_),
    .B(_2674_),
    .C(_2671_),
    .Y(_2688_)
);

BUFX2 _23883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[1]),
    .Y(y[1])
);

AOI21X1 _23463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1840_),
    .C(_1741_),
    .Y(_1841_)
);

AOI21X1 _23043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1372_),
    .B(_1373_),
    .C(_1226_),
    .Y(_1383_)
);

FILL SFILL28920x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5496_),
    .B(_5174_),
    .C(_5166_),
    .Y(_5498_)
);

NAND3X1 _15511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5032_),
    .B(_5031_),
    .C(_5019_),
    .Y(_5037_)
);

NOR3X1 _20588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10250_),
    .B(_10265_),
    .C(_10254_),
    .Y(_10603_)
);

OAI21X1 _20168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9826_),
    .B(_9793_),
    .C(_9819_),
    .Y(_10142_)
);

OAI21X1 _16716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6256_),
    .B(_6251_),
    .C(_6258_),
    .Y(_6358_)
);

OAI21X1 _19188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9057_),
    .B(_9058_),
    .C(_9055_),
    .Y(_9068_)
);

FILL SFILL63960x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18920x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10299_),
    .B(_10255_),
    .C(_10310_),
    .Y(_10321_)
);

AOI21X1 _12216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4226_),
    .B(_4632_),
    .C(_4664_),
    .Y(_5716_)
);

OAI21X1 _22734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf2),
    .B(_8759_),
    .C(_852_),
    .Y(_1046_)
);

NAND2X1 _22314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_320_),
    .B(_324_),
    .Y(_586_)
);

FILL SFILL18840x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 _23939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[57]),
    .Y(y[57])
);

NAND2X1 _23519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1898_),
    .B(_1899_),
    .Y(_1900_)
);

AOI21X1 _17674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6960_),
    .B(_6983_),
    .C(_6986_),
    .Y(_7408_)
);

NAND3X1 _17254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6941_),
    .B(_6943_),
    .C(_6942_),
    .Y(_6948_)
);

FILL SFILL74360x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10477_),
    .B(_10479_),
    .C(_10486_),
    .Y(_10835_)
);

OAI21X1 _18879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8723_),
    .B(_8727_),
    .C(_8728_),
    .Y(_8729_)
);

NAND3X1 _18459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8263_),
    .B(_8265_),
    .C(_8264_),
    .Y(_8269_)
);

AOI21X1 _18039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7800_),
    .B(_7798_),
    .C(_7795_),
    .Y(_7808_)
);

AOI21X1 _13594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2919_),
    .B(_2923_),
    .C(_2840_),
    .Y(_2939_)
);

OAI21X1 _13174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2478_),
    .C(_2476_),
    .Y(_2479_)
);

AND2X2 _23692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2087_),
    .Y(_2090_)
);

NAND2X1 _23272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1513_),
    .Y(_1633_)
);

AND2X2 _19820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9702_),
    .B(_9759_),
    .Y(_9761_)
);

AOI21X1 _19400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9291_),
    .B(_9289_),
    .C(_9286_),
    .Y(_9300_)
);

FILL SFILL69080x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4248_),
    .B(_4246_),
    .C(_4244_),
    .Y(_4256_)
);

NAND3X1 _14379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3794_),
    .B(_3796_),
    .C(_3795_),
    .Y(_3797_)
);

DFFPOSX1 _24057_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[15]),
    .CLK(clk_bF$buf8),
    .D(b[15])
);

AOI21X1 _15740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5286_),
    .B(_5287_),
    .C(_5280_),
    .Y(_5288_)
);

NAND3X1 _15320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4826_),
    .B(_4827_),
    .C(_4825_),
    .Y(_4828_)
);

FILL SFILL3640x46050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10059_),
    .B(_10065_),
    .Y(_10393_)
);

XNOR2X1 _16945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6608_),
    .B(_6605_),
    .Y(_6609_)
);

OAI21X1 _16525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf0),
    .B(_3529__bF$buf1),
    .C(_5768_),
    .Y(_6148_)
);

NAND2X1 _16105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf3),
    .B(breg_22_bF$buf3),
    .Y(_5688_)
);

FILL SFILL59080x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _12865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_122_),
    .B(_89_),
    .Y(_921_)
);

NAND3X1 _12445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8194_),
    .B(_8205_),
    .C(_8216_),
    .Y(_8227_)
);

NAND3X1 _22963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1146_),
    .C(_1149_),
    .Y(_1296_)
);

INVX1 _12025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3613_),
    .Y(_3624_)
);

OAI21X1 _22543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(_831_),
    .C(_662_),
    .Y(_837_)
);

INVX1 _22123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .Y(_377_)
);

FILL SFILL33880x51050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _23748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2129_),
    .B(_2149_),
    .Y(_2150_)
);

INVX2 _23328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1692_),
    .Y(_1693_)
);

NOR3X1 _17483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7193_),
    .B(_7194_),
    .C(_7192_),
    .Y(_7199_)
);

AOI21X1 _17063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6733_),
    .B(_6732_),
    .C(_6731_),
    .Y(_6739_)
);

FILL SFILL49000x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _18688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8516_),
    .B(_8517_),
    .C(_8518_),
    .Y(_8519_)
);

AOI21X1 _18268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7219_),
    .B(_7628_),
    .C(_8059_),
    .Y(_8060_)
);

NAND2X1 _23081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1420_),
    .B(_1422_),
    .Y(_1424_)
);

INVX1 _21814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_33_),
    .Y(_38_)
);

OAI21X1 _14188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3579_),
    .B(_3581_),
    .C(_3577_),
    .Y(_3588_)
);

FILL SFILL53880x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8760x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _16754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6045_),
    .Y(_6400_)
);

OAI21X1 _16334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5939_),
    .B(_5934_),
    .C(_5930_),
    .Y(_5940_)
);

BUFX2 BUFX2_insert180 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_549__bF$buf1)
);

BUFX2 BUFX2_insert181 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .Y(_549__bF$buf0)
);

BUFX2 BUFX2_insert182 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(areg_9_bF$buf4)
);

BUFX2 BUFX2_insert183 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(areg_9_bF$buf3)
);

BUFX2 BUFX2_insert184 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(areg_9_bF$buf2)
);

NAND3X1 _17959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7717_),
    .B(_7719_),
    .C(_7718_),
    .Y(_7720_)
);

BUFX2 BUFX2_insert185 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(areg_9_bF$buf1)
);

AOI21X1 _17539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7255_),
    .B(_7258_),
    .C(_7231_),
    .Y(_7259_)
);

BUFX2 BUFX2_insert186 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[9]),
    .Y(areg_9_bF$buf0)
);

NAND3X1 _17119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6787_),
    .B(_6792_),
    .C(_6794_),
    .Y(_6800_)
);

BUFX2 BUFX2_insert187 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551_),
    .Y(_4551__bF$buf4)
);

BUFX2 BUFX2_insert188 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551_),
    .Y(_4551__bF$buf3)
);

NAND2X1 _12674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_8_bF$buf4),
    .Y(_10737_)
);

BUFX2 BUFX2_insert189 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551_),
    .Y(_4551__bF$buf2)
);

NOR2X1 _12254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_5420__bF$buf2),
    .Y(_6132_)
);

NOR2X1 _22772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_1087_),
    .Y(_1088_)
);

XOR2X1 _22352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_378_),
    .B(_627_),
    .Y(_628_)
);

OAI21X1 _18900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf4),
    .B(_7520__bF$buf0),
    .C(_8743_),
    .Y(_8752_)
);

INVX1 _13879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3249_),
    .Y(_3250_)
);

AND2X2 _13459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2786_),
    .B(_2789_),
    .Y(_2790_)
);

DFFPOSX1 _23977_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[31]),
    .CLK(clk_bF$buf6),
    .D(_0_[31])
);

AOI21X1 _13039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2326_),
    .C(_1478_),
    .Y(_2334_)
);

OAI21X1 _23557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1942_),
    .B(_1938_),
    .C(_1867_),
    .Y(_1943_)
);

FILL SFILL3720x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _23137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1471_),
    .B(_1464_),
    .C(_1469_),
    .Y(_1485_)
);

FILL SFILL43960x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL74360x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4279_),
    .B(_4273_),
    .C(_4202_),
    .Y(_4280_)
);

NOR2X1 _14400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3595_),
    .B(_3596_),
    .Y(_3820_)
);

NAND3X1 _17292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6959_),
    .B(_6984_),
    .C(_6989_),
    .Y(_6990_)
);

FILL SFILL43880x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL23880x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4816_),
    .B(_4839_),
    .C(_4842_),
    .Y(_5140_)
);

FILL SFILL59080x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _18497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8287_),
    .B(_8284_),
    .Y(_8311_)
);

NAND3X1 _18077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7844_),
    .B(_7845_),
    .C(_7846_),
    .Y(_7850_)
);

FILL FILL74040x3050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64360x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _11945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2738_),
    .B(_2716_),
    .Y(_2749_)
);

NAND2X1 _21623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11731_),
    .B(_11732_),
    .Y(_11737_)
);

NOR2X1 _21203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10960_),
    .B(_11277_),
    .Y(_11278_)
);

NAND2X1 _22828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(_1039_),
    .Y(_1148_)
);

NAND3X1 _22408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_671_),
    .C(_672_),
    .Y(_688_)
);

OAI21X1 _16983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6345_),
    .B(_6649_),
    .C(_6335_),
    .Y(_6650_)
);

AOI21X1 _16563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6172_),
    .B(_6175_),
    .C(_6179_),
    .Y(_6190_)
);

NAND3X1 _16143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5726_),
    .B(_5728_),
    .C(_5729_),
    .Y(_5730_)
);

FILL SFILL49000x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18840x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _17768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7506_),
    .B(_7510_),
    .Y(_7511_)
);

NAND3X1 _17348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7050_),
    .B(_7044_),
    .C(_7049_),
    .Y(_7051_)
);

NAND2X1 _12483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7207_),
    .B(_8632_),
    .Y(_8643_)
);

NOR2X1 _12063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4030_),
    .B(_4019_),
    .Y(_0_[6])
);

OR2X2 _22581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_839_),
    .Y(_879_)
);

FILL SFILL23880x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _22161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_410_),
    .C(_414_),
    .Y(_419_)
);

FILL SFILL39080x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2988_),
    .B(_3036_),
    .C(_3040_),
    .Y(_3041_)
);

NOR2X1 _13268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf1),
    .B(_2379_),
    .Y(_2581_)
);

OR2X2 _23786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2129_),
    .B(_2149_),
    .Y(_2191_)
);

FILL SFILL23800x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1733_),
    .C(_1734_),
    .Y(_1735_)
);

AND2X2 _19914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_10_bF$buf4),
    .B(areg_27_bF$buf3),
    .Y(_9865_)
);

FILL SFILL8840x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39000x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13880x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5382_),
    .B(_5383_),
    .Y(_5391_)
);

NAND3X1 _15414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4673_),
    .B(_4931_),
    .C(_4923_),
    .Y(_4932_)
);

FILL SFILL53960x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL29080x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6244_),
    .B(_6249_),
    .C(_6250_),
    .Y(_6251_)
);

NAND3X1 _21852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_76_),
    .B(_79_),
    .C(_77_),
    .Y(_80_)
);

OAI21X1 _21432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586__bF$buf2),
    .B(_8759_),
    .C(_11228_),
    .Y(_11529_)
);

INVX1 _21012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11061_),
    .Y(_11068_)
);

OAI21X1 _12959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf5),
    .B(_5190__bF$buf1),
    .C(_177_),
    .Y(_1947_)
);

NOR3X1 _12539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9192_),
    .B(_9214_),
    .C(_9203_),
    .Y(_9257_)
);

OR2X2 _12119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4215_),
    .B(_4193_),
    .Y(_4653_)
);

AOI22X1 _22637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(_938_),
    .C(_718_),
    .D(_920_),
    .Y(_939_)
);

NAND3X1 _22217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_243_),
    .B(_474_),
    .C(_475_),
    .Y(_480_)
);

FILL SFILL19000x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3269_),
    .B(_3272_),
    .C(_3265_),
    .Y(_3273_)
);

AND2X2 _16792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6081_),
    .B(_6073_),
    .Y(_6441_)
);

NAND3X1 _16372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5978_),
    .B(_5979_),
    .C(_5980_),
    .Y(_5981_)
);

OAI21X1 _17997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7757_),
    .B(_7758_),
    .C(_7708_),
    .Y(_7762_)
);

OAI21X1 _17577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6931_),
    .B(_7300_),
    .C(_6953_),
    .Y(_7301_)
);

OAI21X1 _17157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6840_),
    .B(_6838_),
    .C(_6436_),
    .Y(_6841_)
);

OAI21X1 _12292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6538_),
    .B(_6527_),
    .C(_6516_),
    .Y(_6549_)
);

AOI21X1 _22390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_607_),
    .C(_668_),
    .Y(_669_)
);

NAND3X1 _20703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10702_),
    .B(_10727_),
    .C(_10728_),
    .Y(_10729_)
);

AOI21X1 _13497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2629_),
    .B(_2644_),
    .C(_2831_),
    .Y(_2832_)
);

OAI21X1 _13077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2371_),
    .B(_1489_),
    .C(_1762_),
    .Y(_2372_)
);

NAND3X1 _23595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1982_),
    .B(_1652_),
    .C(_1983_),
    .Y(_1984_)
);

INVX2 _23175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .Y(_1527_)
);

AND2X2 _19723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf4),
    .B(breg_28_bF$buf2),
    .Y(_9655_)
);

NAND2X1 _19303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9184_),
    .B(_9186_),
    .Y(_9195_)
);

AOI21X1 _21908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11812_),
    .B(_140_),
    .C(_11814_),
    .Y(_141_)
);

NOR2X1 _15643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4258__bF$buf1),
    .B(_3958__bF$buf2),
    .Y(_5182_)
);

NAND3X1 _15223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4712_),
    .B(_4720_),
    .C(_4721_),
    .Y(_4722_)
);

FILL SFILL18600x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6499_),
    .B(_6500_),
    .C(_6501_),
    .Y(_6502_)
);

NOR2X1 _16428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6040_),
    .B(_4962_),
    .Y(_6041_)
);

AOI21X1 _16008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5567_),
    .B(_5571_),
    .C(_5554_),
    .Y(_5582_)
);

OAI22X1 _11983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2442_),
    .B(_3055_),
    .C(_3154_),
    .D(_3077_),
    .Y(_3165_)
);

FILL SFILL23880x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11774_),
    .B(_11775_),
    .C(_11777_),
    .Y(_11779_)
);

OAI21X1 _21241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11047_),
    .B(_11017_),
    .C(_11054_),
    .Y(_11319_)
);

NAND2X1 _12768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg_10_bF$buf3),
    .Y(_11767_)
);

NAND2X1 _12348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7109_),
    .B(_7153_),
    .Y(_7164_)
);

AOI21X1 _22866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(_1052_),
    .C(_1189_),
    .Y(_1190_)
);

INVX1 _22446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .Y(_730_)
);

OAI21X1 _22026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_268_),
    .C(_258_),
    .Y(_270_)
);

OAI21X1 _16181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5770_),
    .B(_5769_),
    .C(_5754_),
    .Y(_5772_)
);

OAI21X1 _14914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4373_),
    .B(_4372_),
    .C(_4370_),
    .Y(_4383_)
);

OAI21X1 _17386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7092_),
    .B(_6717_),
    .C(_6708_),
    .Y(_7093_)
);

FILL SFILL13800x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10964_),
    .B(_10971_),
    .C(_10974_),
    .Y(_10981_)
);

AOI21X1 _20512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10239_),
    .B(_10519_),
    .C(_10517_),
    .Y(_10520_)
);

NOR2X1 _19952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9905_),
    .B(_9535_),
    .Y(_9906_)
);

NAND2X1 _19532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf4),
    .B(areg_23_bF$buf1),
    .Y(_9446_)
);

NAND3X1 _19112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8979_),
    .B(_8984_),
    .C(_8933_),
    .Y(_8985_)
);

AOI21X1 _21717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11556_),
    .B(_11554_),
    .C(_11562_),
    .Y(_11840_)
);

NOR3X1 _15872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5425_),
    .B(_5428_),
    .C(_5424_),
    .Y(_5433_)
);

INVX2 _15452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4662_),
    .Y(_4972_)
);

NAND2X1 _15032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4219_),
    .B(_4238_),
    .Y(_4513_)
);

FILL SFILL64040x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6292_),
    .B(_5950_),
    .C(_5941_),
    .Y(_6293_)
);

NAND3X1 _16237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5818_),
    .B(_5823_),
    .C(_5822_),
    .Y(_5833_)
);

XNOR2X1 _21890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_95_),
    .Y(_121_)
);

OAI21X1 _21470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11566_),
    .B(_11569_),
    .C(_11322_),
    .Y(_11570_)
);

OAI21X1 _21050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11107_),
    .B(_11108_),
    .C(_11104_),
    .Y(_11109_)
);

OAI21X1 _12997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2291_),
    .B(_2290_),
    .C(_2259_),
    .Y(_2292_)
);

AOI21X1 _12577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9609_),
    .B(_9620_),
    .C(_8511_),
    .Y(_9674_)
);

AND2X2 _12157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5036_),
    .B(_5047_),
    .Y(_5069_)
);

OAI21X1 _22675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_797_),
    .B(_796_),
    .C(_788_),
    .Y(_981_)
);

AOI21X1 _22255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_265_),
    .C(_268_),
    .Y(_521_)
);

NAND3X1 _18803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8640_),
    .B(_8645_),
    .C(_8642_),
    .Y(_8646_)
);

FILL SFILL54040x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4172_),
    .B(_4173_),
    .C(_4164_),
    .Y(_4174_)
);

OAI21X1 _14303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3714_),
    .B(_3707_),
    .C(_3639_),
    .Y(_3715_)
);

AOI21X1 _17195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6876_),
    .B(_6877_),
    .C(_6875_),
    .Y(_6883_)
);

FILL SFILL44440x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5480_),
    .B(_5484_),
    .C(_5487_),
    .Y(_5494_)
);

NAND3X1 _15508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5018_),
    .B(_5032_),
    .C(_5031_),
    .Y(_5033_)
);

NAND3X1 _20741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10767_),
    .B(_10768_),
    .C(_10769_),
    .Y(_10771_)
);

NAND3X1 _20321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10305_),
    .B(_10309_),
    .C(_9995_),
    .Y(_10311_)
);

FILL SFILL44040x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9695_),
    .B(_9694_),
    .C(_9691_),
    .Y(_9697_)
);

AOI21X1 _19341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9234_),
    .B(_9235_),
    .C(_8887_),
    .Y(_9237_)
);

NOR3X1 _21946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_170_),
    .C(_165_),
    .Y(_183_)
);

NOR3X1 _21526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11630_),
    .B(_11626_),
    .C(_11629_),
    .Y(_11631_)
);

INVX1 _21106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11170_),
    .Y(_11171_)
);

NAND3X1 _15681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5217_),
    .B(_5178_),
    .C(_5222_),
    .Y(_5223_)
);

NAND3X1 _15261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4751_),
    .B(_4753_),
    .C(_4747_),
    .Y(_4764_)
);

AOI21X1 _16886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6542_),
    .B(_6543_),
    .C(_6541_),
    .Y(_6544_)
);

INVX1 _16466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6059_),
    .Y(_6082_)
);

FILL SFILL74120x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _16046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5606_),
    .B(_5612_),
    .C(_5461_),
    .Y(_5624_)
);

INVX2 _12386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7569_),
    .Y(_7580_)
);

OAI21X1 _22484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_580_),
    .B(_771_),
    .C(_574_),
    .Y(_772_)
);

OAI22X1 _22064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11721_),
    .B(_311_),
    .C(_99_),
    .D(_95_),
    .Y(_312_)
);

OAI21X1 _18612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8429_),
    .B(_8436_),
    .C(_8078_),
    .Y(_8437_)
);

FILL SFILL74040x50 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _23689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2031_),
    .Y(_2086_)
);

AND2X2 _23269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1627_),
    .Y(_1629_)
);

NAND2X1 _19817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_14_bF$buf3),
    .B(breg_23_bF$buf1),
    .Y(_9758_)
);

AOI21X1 _14952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4413_),
    .B(_4409_),
    .C(_4391_),
    .Y(_4425_)
);

NAND2X1 _14532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3685_),
    .B(_3959_),
    .Y(_3966_)
);

NAND2X1 _14112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1206_),
    .B(_1217_),
    .Y(_3505_)
);

AOI21X1 _15737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4943_),
    .B(_4654_),
    .C(_4945_),
    .Y(_5285_)
);

INVX1 _15317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4819_),
    .Y(_4825_)
);

OAI21X1 _20970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10716_),
    .B(_10706_),
    .C(_10710_),
    .Y(_11021_)
);

OAI21X1 _20550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10227_),
    .B(_10216_),
    .C(_10220_),
    .Y(_10561_)
);

AOI21X1 _20130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9757_),
    .B(_9842_),
    .C(_9852_),
    .Y(_10100_)
);

BUFX2 BUFX2_insert95 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf5)
);

BUFX2 BUFX2_insert96 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf4)
);

BUFX2 BUFX2_insert97 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf3)
);

BUFX2 BUFX2_insert98 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf2)
);

BUFX2 BUFX2_insert99 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[19]),
    .Y(breg_19_bF$buf1)
);

NAND3X1 _19990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9743_),
    .B(_9747_),
    .C(_9749_),
    .Y(_9947_)
);

XNOR2X1 _19570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9486_),
    .B(_9484_),
    .Y(_9487_)
);

OAI21X1 _19150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9025_),
    .B(_9024_),
    .C(_9015_),
    .Y(_9026_)
);

OAI21X1 _21755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11637_),
    .B(_11606_),
    .C(_11644_),
    .Y(_11881_)
);

NAND3X1 _21335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11405_),
    .B(_11412_),
    .C(_11410_),
    .Y(_11422_)
);

NOR2X1 _15490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4679_),
    .B(_5012_),
    .Y(_5013_)
);

AOI21X1 _15070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4552_),
    .B(_4553_),
    .C(_4537_),
    .Y(_4554_)
);

OAI21X1 _13803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3149_),
    .B(_3155_),
    .C(_3157_),
    .Y(_3168_)
);

BUFX2 _23901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[19]),
    .Y(y[19])
);

NAND3X1 _16695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6293_),
    .B(_6334_),
    .C(_6329_),
    .Y(_6335_)
);

AOI21X1 _16275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5865_),
    .B(_5858_),
    .C(_5845_),
    .Y(_5875_)
);

FILL SFILL44040x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5475_),
    .B(_5431_),
    .Y(_5486_)
);

OAI21X1 _22293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf3),
    .B(_5315__bF$buf2),
    .C(_546_),
    .Y(_563_)
);

AND2X2 _18841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8269_),
    .B(_8264_),
    .Y(_8688_)
);

INVX1 _18421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8226_),
    .Y(_8228_)
);

OAI21X1 _18001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7765_),
    .B(_7344_),
    .C(_7422_),
    .Y(_7767_)
);

NAND3X1 _20606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10449_),
    .B(_10454_),
    .C(_10456_),
    .Y(_10623_)
);

NOR2X1 _23498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(_1877_),
    .Y(_1878_)
);

OAI21X1 _23078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4551__bF$buf2),
    .B(_6427_),
    .C(_1419_),
    .Y(_1420_)
);

AOI21X1 _19626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9545_),
    .B(_9548_),
    .C(_9529_),
    .Y(_9549_)
);

OAI21X1 _19206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8737_),
    .B(_8736_),
    .C(_8734_),
    .Y(_9087_)
);

OAI21X1 _14761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_2669__bF$buf0),
    .C(_4209_),
    .Y(_4216_)
);

NAND3X1 _14341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3520_),
    .B(_3751_),
    .C(_3750_),
    .Y(_3757_)
);

FILL SFILL34040x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5531_),
    .B(_5532_),
    .C(_5527_),
    .Y(_5536_)
);

OAI21X1 _15546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5060_),
    .B(_5061_),
    .C(_5057_),
    .Y(_5075_)
);

NAND3X1 _15126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4598_),
    .B(_4605_),
    .C(_4608_),
    .Y(_4616_)
);

AOI21X1 _21984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_224_),
    .B(_218_),
    .C(_11882_),
    .Y(_225_)
);

INVX1 _21564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11649_),
    .Y(_11672_)
);

NAND3X1 _21144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11205_),
    .B(_11212_),
    .C(_11210_),
    .Y(_11213_)
);

FILL SFILL23800x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL64280x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28760x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59160x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _22769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_1080_),
    .C(_946_),
    .Y(_1084_)
);

FILL SFILL64120x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3640x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_622_),
    .C(_623_),
    .Y(_624_)
);

NOR3X1 _13612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .B(_2726_),
    .C(_2724_),
    .Y(_2959_)
);

OAI21X1 _23710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2106_),
    .B(_1398_),
    .C(_1536_),
    .Y(_2108_)
);

OAI21X1 _16084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5644_),
    .B(_5305_),
    .C(_5634_),
    .Y(_5665_)
);

OAI21X1 _14817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4271_),
    .B(_4269_),
    .C(_4235_),
    .Y(_4277_)
);

NOR3X1 _17289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6980_),
    .B(_6982_),
    .C(_6979_),
    .Y(_6986_)
);

OAI21X1 _18650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8476_),
    .B(_8076_),
    .C(_8444_),
    .Y(_8477_)
);

AOI21X1 _18230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8016_),
    .B(_8017_),
    .C(_8015_),
    .Y(_8018_)
);

FILL SFILL54120x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10580_),
    .B(_10873_),
    .C(_10872_),
    .Y(_10874_)
);

NOR2X1 _20415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10056_),
    .B(_10114_),
    .Y(_10413_)
);

NAND3X1 _19855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9796_),
    .B(_9799_),
    .C(_9798_),
    .Y(_9800_)
);

OAI21X1 _19435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287__bF$buf3),
    .B(_3781__bF$buf1),
    .C(_8948_),
    .Y(_9339_)
);

NOR3X1 _19015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8865_),
    .B(_8868_),
    .C(_8871_),
    .Y(_8878_)
);

NOR2X1 _14990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4457_),
    .B(_4458_),
    .Y(_4465_)
);

NAND2X1 _14570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4006_),
    .B(_4005_),
    .Y(_4007_)
);

NOR2X1 _14150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3542_),
    .Y(_3546_)
);

FILL SFILL59400x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59320x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5319_),
    .B(_5320_),
    .C(_5309_),
    .Y(_5326_)
);

FILL SFILL39160x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4538_),
    .B(_4542_),
    .C(_4546_),
    .Y(_4867_)
);

AOI21X1 _21793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11608_),
    .B(_11633_),
    .C(_11631_),
    .Y(_15_)
);

NAND3X1 _21373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11460_),
    .B(_11462_),
    .C(_11463_),
    .Y(_11464_)
);

NAND3X1 _17921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7673_),
    .B(_7677_),
    .C(_7676_),
    .Y(_7679_)
);

NOR2X1 _17501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7204_),
    .B(_7216_),
    .Y(_7218_)
);

NAND3X1 _22998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(_1319_),
    .C(_1323_),
    .Y(_1333_)
);

XOR2X1 _22578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_864_),
    .Y(_875_)
);

OAI21X1 _22158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_410_),
    .C(_413_),
    .Y(_415_)
);

OAI21X1 _18706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf3),
    .B(_5315__bF$buf3),
    .C(_8531_),
    .Y(_8539_)
);

FILL SFILL69240x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _13841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3190_),
    .B(_3194_),
    .C(_3197_),
    .Y(_3210_)
);

NAND2X1 _13421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2748_),
    .B(_2744_),
    .Y(_2750_)
);

NOR2X1 _13001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2259_),
    .B(_2295_),
    .Y(_2296_)
);

FILL SFILL34040x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _14626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3808_),
    .B(_4066_),
    .C(_3856_),
    .Y(_4067_)
);

INVX2 _14206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3601_),
    .Y(_3607_)
);

OAI21X1 _17098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6775_),
    .B(_6776_),
    .C(_6774_),
    .Y(_6777_)
);

AOI21X1 _20644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8872_),
    .B(_8873_),
    .C(_8871_),
    .Y(_10664_)
);

NAND3X1 _20224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10201_),
    .B(_10203_),
    .C(_10202_),
    .Y(_10204_)
);

AOI21X1 _19664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9590_),
    .B(_9584_),
    .C(_9387_),
    .Y(_9591_)
);

OAI21X1 _19244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9123_),
    .B(_9128_),
    .C(_9129_),
    .Y(_9130_)
);

FILL SFILL59160x39050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _21849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_22_),
    .B(_19_),
    .Y(_76_)
);

NOR2X1 _21429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2379_),
    .B(_7520__bF$buf1),
    .Y(_11525_)
);

NOR2X1 _21009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11062_),
    .B(_11063_),
    .Y(_11064_)
);

NAND3X1 _15584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5111_),
    .B(_5116_),
    .C(_5115_),
    .Y(_5117_)
);

OAI21X1 _15164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4367_),
    .B(_4385_),
    .C(_4384_),
    .Y(_4657_)
);

FILL FILL74120x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49240x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5726_),
    .B(_6049_),
    .C(_6434_),
    .Y(_6437_)
);

NAND2X1 _16369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5976_),
    .B(_5977_),
    .Y(_5978_)
);

NAND3X1 _21182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11221_),
    .B(_11222_),
    .C(_11223_),
    .Y(_11255_)
);

FILL SFILL49160x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7467_),
    .B(_7468_),
    .C(_7466_),
    .Y(_7469_)
);

NAND3X1 _17310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6924_),
    .B(_7004_),
    .C(_7008_),
    .Y(_7009_)
);

FILL SFILL33960x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _12289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6472_),
    .Y(_6516_)
);

OAI21X1 _22387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_665_),
    .C(_663_),
    .Y(_666_)
);

AOI21X1 _18935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8389_),
    .B(_8387_),
    .C(_8396_),
    .Y(_8791_)
);

AOI21X1 _18515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7983_),
    .B(_7982_),
    .C(_7957_),
    .Y(_8331_)
);

OAI21X1 _13650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2763_),
    .C(_2998_),
    .Y(_2999_)
);

INVX1 _13230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2538_),
    .Y(_2539_)
);

FILL SFILL39160x35050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4301_),
    .B(_4308_),
    .C(_4311_),
    .Y(_4319_)
);

OAI21X1 _14435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3856_),
    .B(_3857_),
    .C(_3858_),
    .Y(_3859_)
);

AND2X2 _14015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf3),
    .B(areg_18_bF$buf3),
    .Y(_3399_)
);

OAI21X1 _20873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10567_),
    .B(_10563_),
    .C(_10566_),
    .Y(_10916_)
);

NAND3X1 _20453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10349_),
    .B(_10449_),
    .C(_10454_),
    .Y(_10455_)
);

AOI21X1 _20033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9957_),
    .B(_9958_),
    .C(_9644_),
    .Y(_9994_)
);

OAI21X1 _19893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9838_),
    .B(_9830_),
    .C(_9841_),
    .Y(_9842_)
);

OAI21X1 _19473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9377_),
    .B(_9379_),
    .C(_9380_),
    .Y(_9381_)
);

OAI21X1 _19053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8915_),
    .B(_8916_),
    .C(_8912_),
    .Y(_8920_)
);

FILL SFILL69320x22050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11762_),
    .B(_11760_),
    .C(_11757_),
    .Y(_11775_)
);

NOR2X1 _21238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11312_),
    .B(_11314_),
    .Y(_11315_)
);

FILL SFILL69240x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _12921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1522_),
    .B(_1500_),
    .Y(_1533_)
);

OAI22X1 _12501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6385_),
    .B(_7591_),
    .C(_7580_),
    .D(_7623_),
    .Y(_8851_)
);

AOI21X1 _15393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4495_),
    .B(_4583_),
    .C(_4908_),
    .Y(_4909_)
);

NOR2X1 _13706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4434__bF$buf3),
    .B(_8555_),
    .Y(_3061_)
);

OAI21X1 _23804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .B(_2155_),
    .C(_2201_),
    .Y(_2210_)
);

INVX2 _16598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6227_),
    .Y(_6228_)
);

NAND2X1 _16178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_19_bF$buf1),
    .Y(_5768_)
);

FILL SFILL3800x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59240x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_1_bF$buf6),
    .B(areg_7_bF$buf1),
    .Y(_4423_)
);

NAND2X1 _22196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_455_),
    .Y(_457_)
);

NAND3X1 _18744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8572_),
    .B(_8580_),
    .C(_8525_),
    .Y(_8581_)
);

AND2X2 _18324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8116_),
    .B(_8120_),
    .Y(_8121_)
);

NAND3X1 _20929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10975_),
    .B(_10976_),
    .C(_10974_),
    .Y(_10977_)
);

AOI21X1 _20509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10505_),
    .B(_10504_),
    .C(_10501_),
    .Y(_10516_)
);

FILL FILL74200x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9149_),
    .B(_9901_),
    .C(_9539_),
    .Y(_9902_)
);

NAND3X1 _19529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9441_),
    .B(_9435_),
    .C(_9438_),
    .Y(_9442_)
);

AOI21X1 _19109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8977_),
    .B(_8976_),
    .C(_8975_),
    .Y(_8981_)
);

NOR2X1 _14664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3870_),
    .B(_3871_),
    .Y(_4109_)
);

OAI21X1 _14244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf4),
    .B(_549__bF$buf3),
    .C(_3644_),
    .Y(_3650_)
);

FILL FILL74120x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5424_),
    .B(_5425_),
    .C(_5428_),
    .Y(_5429_)
);

AOI21X1 _15449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4915_),
    .B(_4922_),
    .C(_4676_),
    .Y(_4968_)
);

OAI21X1 _15029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4116__bF$buf3),
    .B(_2669__bF$buf0),
    .C(_4504_),
    .Y(_4509_)
);

NAND2X1 _20682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_11_bF$buf4),
    .B(breg_29_bF$buf0),
    .Y(_10706_)
);

AOI21X1 _20262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9536_),
    .B(_9539_),
    .C(_9911_),
    .Y(_10246_)
);

AOI21X1 _16810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6449_),
    .B(_6448_),
    .C(_6445_),
    .Y(_6460_)
);

AOI21X1 _19282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9169_),
    .B(_9171_),
    .C(_9168_),
    .Y(_9172_)
);

FILL SFILL33960x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_106_),
    .C(_104_),
    .Y(_118_)
);

NAND3X1 _21467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11564_),
    .B(_11561_),
    .C(_11325_),
    .Y(_11567_)
);

OAI21X1 _21047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11092_),
    .B(_11093_),
    .C(_11090_),
    .Y(_11106_)
);

NOR3X1 _12730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11329_),
    .B(_11318_),
    .C(_11350_),
    .Y(_11361_)
);

AOI21X1 _12310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6736_),
    .B(_6725_),
    .C(_6659_),
    .Y(_6747_)
);

NOR2X1 _13935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2825__bF$buf1),
    .B(_2379_),
    .Y(_3312_)
);

OAI21X1 _13515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5420__bF$buf0),
    .B(_6582__bF$buf3),
    .C(_2851_),
    .Y(_2852_)
);

INVX1 _23613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .Y(_2004_)
);

FILL SFILL23960x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69400x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8825_),
    .B(_8832_),
    .C(_8601_),
    .Y(_8833_)
);

OAI21X1 _18553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8372_),
    .B(_8371_),
    .C(_8362_),
    .Y(_8373_)
);

OAI21X1 _18133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7894_),
    .B(_7899_),
    .C(_7901_),
    .Y(_7912_)
);

FILL SFILL69320x17050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10743_),
    .Y(_10767_)
);

OAI21X1 _20318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10302_),
    .B(_10303_),
    .C(_9998_),
    .Y(_10307_)
);

NAND2X1 _19758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_13_bF$buf4),
    .B(breg_24_bF$buf3),
    .Y(_9693_)
);

AOI21X1 _19338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9232_),
    .B(_9227_),
    .C(_8888_),
    .Y(_9233_)
);

AOI21X1 _14893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4287_),
    .B(_4294_),
    .C(_4154_),
    .Y(_4360_)
);

AOI21X1 _14473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3641_),
    .B(_3660_),
    .C(_3663_),
    .Y(_3901_)
);

AOI21X1 _14053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3424_),
    .B(_3429_),
    .C(_3385_),
    .Y(_3441_)
);

AOI21X1 _15678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5215_),
    .B(_5214_),
    .C(_5213_),
    .Y(_5220_)
);

NOR2X1 _15258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4424_),
    .B(_4425_),
    .Y(_4760_)
);

OAI21X1 _20491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10171_),
    .B(_10169_),
    .C(_10160_),
    .Y(_10497_)
);

NOR3X1 _20071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10032_),
    .B(_10033_),
    .C(_10034_),
    .Y(_10036_)
);

NAND3X1 _19091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8957_),
    .B(_8943_),
    .C(_8947_),
    .Y(_8962_)
);

XNOR2X1 _21696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11816_),
    .B(_11812_),
    .Y(_11817_)
);

NAND3X1 _21276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11331_),
    .B(_11354_),
    .C(_11355_),
    .Y(_11356_)
);

NAND3X1 _17824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7566_),
    .B(_7572_),
    .C(_7483_),
    .Y(_7573_)
);

AOI22X1 _17404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf2),
    .B(areg_30_bF$buf5),
    .C(breg_1_bF$buf5),
    .D(areg_29_bF$buf4),
    .Y(_7113_)
);

NAND3X1 _18609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8426_),
    .B(_8427_),
    .C(_8187_),
    .Y(_8433_)
);

AND2X2 _13744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf4),
    .B(areg_12_bF$buf0),
    .Y(_3103_)
);

INVX1 _13324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .Y(_2643_)
);

XOR2X1 _23842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2248_),
    .B(_2250_),
    .Y(_2251_)
);

OAI21X1 _23422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7100__bF$buf1),
    .B(_5668__bF$buf0),
    .C(_1679_),
    .Y(_1796_)
);

AOI21X1 _23002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(_1329_),
    .C(_1294_),
    .Y(_1338_)
);

NAND3X1 _14949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4399_),
    .B(_4407_),
    .C(_4404_),
    .Y(_4421_)
);

OAI21X1 _14529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551__bF$buf1),
    .B(_3961__bF$buf1),
    .C(_3685_),
    .Y(_3962_)
);

AND2X2 _14109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_3500_),
    .Y(_3501_)
);

NAND3X1 _18782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8609_),
    .B(_8618_),
    .C(_8617_),
    .Y(_8623_)
);

AOI21X1 _18362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7709_),
    .B(_7743_),
    .C(_7747_),
    .Y(_8163_)
);

OAI21X1 _20967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10718_),
    .B(_10703_),
    .C(_10728_),
    .Y(_11018_)
);

NAND2X1 _20547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_27_bF$buf3),
    .Y(_10558_)
);

NAND3X1 _20127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10096_),
    .B(_10095_),
    .C(_10091_),
    .Y(_10097_)
);

OAI21X1 _19987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9942_),
    .B(_9943_),
    .C(_9854_),
    .Y(_9944_)
);

NAND2X1 _19567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_14_bF$buf1),
    .B(areg_22_bF$buf3),
    .Y(_9484_)
);

NAND2X1 _19147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf3),
    .B(breg_18_bF$buf1),
    .Y(_9023_)
);

NAND3X1 _14282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3684_),
    .B(_3687_),
    .C(_3686_),
    .Y(_3692_)
);

FILL SFILL8680x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _15487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_2_bF$buf3),
    .B(breg_23_bF$buf3),
    .Y(_5010_)
);

INVX8 _15067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_22_bF$buf0),
    .Y(_4551_)
);

NAND2X1 _21085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11144_),
    .B(_11141_),
    .Y(_11148_)
);

NAND2X1 _17633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7357_),
    .B(_7358_),
    .Y(_7363_)
);

NAND2X1 _17213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6841_),
    .B(_6843_),
    .Y(_6903_)
);

FILL SFILL74280x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28680x50 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8327_),
    .B(_8325_),
    .C(_8323_),
    .Y(_8684_)
);

AND2X2 _18418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_16_bF$buf3),
    .B(areg_17_bF$buf3),
    .Y(_8224_)
);

AOI21X1 _13973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3058_),
    .B(_3076_),
    .C(_3352_),
    .Y(_3353_)
);

OAI21X1 _13553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2891_),
    .B(_2892_),
    .C(_2876_),
    .Y(_2893_)
);

NAND2X1 _13133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2433_),
    .B(_2430_),
    .Y(_2434_)
);

XNOR2X1 _23651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2044_),
    .B(_1923_),
    .Y(_2046_)
);

OAI22X1 _23231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1348_),
    .B(_1496_),
    .C(_1498_),
    .D(_1495_),
    .Y(_1588_)
);

OAI22X1 _14758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_2669__bF$buf0),
    .C(_4116__bF$buf4),
    .D(_2465__bF$buf0),
    .Y(_4212_)
);

OAI21X1 _14338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3752_),
    .B(_3749_),
    .C(_3519_),
    .Y(_3753_)
);

FILL SFILL64200x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

DFFPOSX1 _24016_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[6]),
    .CLK(clk_bF$buf0),
    .D(a[6])
);

FILL SFILL64200x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8411_),
    .B(_8412_),
    .C(_8410_),
    .Y(_8414_)
);

NAND3X1 _18171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7950_),
    .B(_7951_),
    .C(_7952_),
    .Y(_7954_)
);

OAI21X1 _20776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10802_),
    .B(_10801_),
    .C(_10799_),
    .Y(_10809_)
);

OAI21X1 _20356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10294_),
    .B(_10347_),
    .C(_10283_),
    .Y(_10348_)
);

NAND3X1 _16904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6556_),
    .B(_6559_),
    .C(_6563_),
    .Y(_6564_)
);

OAI21X1 _19796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9733_),
    .B(_9734_),
    .C(_9730_),
    .Y(_9735_)
);

INVX2 _19376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9273_),
    .Y(_9274_)
);

AOI21X1 _14091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2984_),
    .B(_3221_),
    .C(_3481_),
    .Y(_3483_)
);

XNOR2X1 _12824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_418_),
    .Y(_473_)
);

NAND3X1 _12404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7766_),
    .B(_7733_),
    .C(_7656_),
    .Y(_7777_)
);

NAND3X1 _22922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1251_),
    .C(_1246_),
    .Y(_1252_)
);

NOR2X1 _22502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_610_),
    .B(_611_),
    .Y(_792_)
);

AOI21X1 _15296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4798_),
    .B(_4797_),
    .C(_4795_),
    .Y(_4802_)
);

NAND3X1 _13609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2941_),
    .B(_2945_),
    .C(_2949_),
    .Y(_2955_)
);

XNOR2X1 _23707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2105_),
    .Y(_0_[57])
);

AOI21X1 _17862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7609_),
    .B(_7608_),
    .C(_7607_),
    .Y(_7614_)
);

OAI21X1 _17442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7152_),
    .B(_7154_),
    .C(_7151_),
    .Y(_7155_)
);

OAI21X1 _17022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6309_),
    .B(_6314_),
    .C(_6313_),
    .Y(_6694_)
);

OAI21X1 _22099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_346_),
    .C(_295_),
    .Y(_350_)
);

OAI21X1 _18647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8111_),
    .B(_8081_),
    .C(_8119_),
    .Y(_8474_)
);

NAND2X1 _18227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8014_),
    .B(_8013_),
    .Y(_8015_)
);

OAI21X1 _13782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3220_),
    .B(_2884__bF$buf0),
    .C(_3144_),
    .Y(_3145_)
);

AOI21X1 _13362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2679_),
    .B(_2684_),
    .C(_2652_),
    .Y(_2685_)
);

XOR2X1 _23880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3285_),
    .B(_3274_),
    .Y(_0_[3])
);

AOI21X1 _23460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(_1836_),
    .C(_1830_),
    .Y(_1837_)
);

OAI21X1 _23040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(_1378_),
    .C(_1265_),
    .Y(_1379_)
);

NAND3X1 _14987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4456_),
    .B(_4461_),
    .C(_4459_),
    .Y(_4462_)
);

AOI21X1 _14567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4003_),
    .B(_3998_),
    .C(_3913_),
    .Y(_4004_)
);

OR2X2 _14147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3266_),
    .B(_3542_),
    .Y(_3543_)
);

FILL SFILL13640x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _20585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10596_),
    .Y(_10600_)
);

OAI21X1 _20165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10125_),
    .B(_10129_),
    .C(_10131_),
    .Y(_10139_)
);

OAI21X1 _16713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6353_),
    .B(_6354_),
    .C(_6351_),
    .Y(_6355_)
);

INVX1 _19185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8641_),
    .Y(_9065_)
);

FILL SFILL74200x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _17918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_5_bF$buf2),
    .B(breg_27_bF$buf3),
    .Y(_7675_)
);

FILL SFILL44040x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10145_),
    .B(_10079_),
    .C(_10167_),
    .Y(_10288_)
);

NAND2X1 _12213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5596_),
    .B(_5629_),
    .Y(_5683_)
);

AND2X2 _22731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_857_),
    .B(_1041_),
    .Y(_1043_)
);

OAI21X1 _22311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_576_),
    .C(_573_),
    .Y(_583_)
);

FILL SFILL38840x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL43800x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2988_),
    .B(_3043_),
    .C(_3045_),
    .Y(_3206_)
);

NAND3X1 _13418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2527_),
    .B(_2733_),
    .C(_2739_),
    .Y(_2746_)
);

BUFX2 _23936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11909_[54]),
    .Y(y[54])
);

NAND2X1 _23516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1806_),
    .B(_1818_),
    .Y(_1897_)
);

FILL SFILL64200x47050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _17671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7388_),
    .B(_7391_),
    .C(_7394_),
    .Y(_7405_)
);

AOI21X1 _17251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6943_),
    .B(_6942_),
    .C(_6941_),
    .Y(_6945_)
);

OAI21X1 _18876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8708_),
    .B(_8713_),
    .C(_8715_),
    .Y(_8726_)
);

FILL SFILL33800x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8265_),
    .B(_8264_),
    .C(_8263_),
    .Y(_8266_)
);

OAI21X1 _18036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7804_),
    .B(_7803_),
    .C(_7794_),
    .Y(_7805_)
);

NOR3X1 _13591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2699_),
    .B(_2700_),
    .C(_2701_),
    .Y(_2936_)
);

XNOR2X1 _13171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2449_),
    .Y(_2476_)
);

FILL SFILL54200x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4252_),
    .B(_4249_),
    .C(_4242_),
    .Y(_4253_)
);

INVX1 _14376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3789_),
    .Y(_3794_)
);

DFFPOSX1 _24054_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(breg[12]),
    .CLK(clk_bF$buf0),
    .D(b[12])
);

FILL SFILL13720x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _20394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10350_),
    .B(_10389_),
    .C(_10388_),
    .Y(_10390_)
);

NAND2X1 _16942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_17_bF$buf4),
    .Y(_6606_)
);

NOR3X1 _16522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6138_),
    .B(_6140_),
    .C(_6144_),
    .Y(_6145_)
);

NAND2X1 _16102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf3),
    .B(breg_25_bF$buf3),
    .Y(_5685_)
);

FILL SFILL23720x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11709_),
    .B(_11427_),
    .Y(_11710_)
);

NAND3X1 _21179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11249_),
    .B(_11244_),
    .C(_11250_),
    .Y(_11251_)
);

XNOR2X1 _17727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7441_),
    .B(_7465_),
    .Y(_7466_)
);

AOI21X1 _17307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6990_),
    .B(_6996_),
    .C(_6957_),
    .Y(_7006_)
);

NOR3X1 _12862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_385_),
    .C(_790_),
    .Y(_889_)
);

INVX2 _12442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7185_),
    .Y(_8194_)
);

NAND3X1 _22960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1291_),
    .B(_1288_),
    .C(_1285_),
    .Y(_1292_)
);

AOI21X1 _12022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2803_),
    .B(_2836_),
    .C(_3580_),
    .Y(_3591_)
);

AOI21X1 _22540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_832_),
    .C(_732_),
    .Y(_833_)
);

XNOR2X1 _22120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_367_),
    .Y(_372_)
);

NAND2X1 _13647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_16_bF$buf1),
    .Y(_2996_)
);

XNOR2X1 _13227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2356_),
    .B(_2536_),
    .Y(_0_[15])
);

XOR2X1 _23745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2146_),
    .B(_2130_),
    .Y(_2147_)
);

NAND2X1 _23325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1684_),
    .B(_1671_),
    .Y(_1690_)
);

FILL SFILL48840x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL13720x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _17480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7193_),
    .B(_7194_),
    .C(_7192_),
    .Y(_7195_)
);

NAND3X1 _17060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6728_),
    .B(_6734_),
    .C(_6650_),
    .Y(_6735_)
);

FILL SFILL34120x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8083_),
    .B(_8108_),
    .C(_8105_),
    .Y(_8516_)
);

AOI21X1 _18265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8056_),
    .B(_8055_),
    .C(_7655_),
    .Y(_8057_)
);

OAI21X1 _21811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .B(_33_),
    .C(_29_),
    .Y(_35_)
);

FILL SFILL38840x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _14185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3286_),
    .Y(_3585_)
);

NAND2X1 _12918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .B(breg_14_bF$buf2),
    .Y(_1500_)
);

AOI21X1 _16751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6378_),
    .B(_6383_),
    .C(_6127_),
    .Y(_6397_)
);

NAND3X1 _16331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5931_),
    .B(_5935_),
    .C(_5933_),
    .Y(_5937_)
);

FILL SFILL28840x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert150 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .Y(_2376__bF$buf0)
);

BUFX2 BUFX2_insert151 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf5)
);

BUFX2 BUFX2_insert152 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf4)
);

BUFX2 BUFX2_insert153 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf3)
);

INVX1 _17956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7712_),
    .Y(_7717_)
);

BUFX2 BUFX2_insert154 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf2)
);

OAI21X1 _17536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7252_),
    .B(_7253_),
    .C(_7248_),
    .Y(_7256_)
);

BUFX2 BUFX2_insert155 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf1)
);

BUFX2 BUFX2_insert156 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(breg_10_bF$buf0)
);

OAI21X1 _17116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6795_),
    .B(_6796_),
    .C(_6794_),
    .Y(_6797_)
);

BUFX2 BUFX2_insert157 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf5)
);

BUFX2 BUFX2_insert158 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf4)
);

BUFX2 BUFX2_insert159 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5668_),
    .Y(_5668__bF$buf3)
);

OAI21X1 _12671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9247_),
    .B(_9268_),
    .C(_9181_),
    .Y(_10704_)
);

INVX2 _12251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6088_),
    .Y(_6099_)
);

AOI21X1 _13876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3199_),
    .B(_3202_),
    .C(_3049_),
    .Y(_3247_)
);

NAND2X1 _13456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2780_),
    .B(_2783_),
    .Y(_2787_)
);

DFFPOSX1 _23974_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(_11909_[28]),
    .CLK(clk_bF$buf4),
    .D(_0_[28])
);

OAI21X1 _13036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_2330_),
    .C(_2328_),
    .Y(_2331_)
);

AOI21X1 _23554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1934_),
    .B(_1935_),
    .C(_1931_),
    .Y(_1940_)
);

OAI21X1 _23134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1480_),
    .B(_1481_),
    .C(_1479_),
    .Y(_1482_)
);

FILL SFILL18840x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5129_),
    .B(_5134_),
    .C(_5136_),
    .Y(_5137_)
);

OAI21X1 _18494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8307_),
    .B(_8306_),
    .C(_8290_),
    .Y(_8308_)
);

AOI21X1 _18074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7845_),
    .B(_7846_),
    .C(_7844_),
    .Y(_7847_)
);

FILL SFILL44200x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _20679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7711__bF$buf3),
    .B(_6815__bF$buf2),
    .Y(_10702_)
);

NAND3X1 _20259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10230_),
    .B(_10224_),
    .C(_10228_),
    .Y(_10242_)
);

OAI22X1 _16807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5750_),
    .B(_6455_),
    .C(_6456_),
    .D(_6131_),
    .Y(_6457_)
);

NAND2X1 _11942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_5_bF$buf1),
    .B(areg[0]),
    .Y(_2716_)
);

NOR2X1 _21620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11731_),
    .B(_11732_),
    .Y(_11733_)
);

AOI21X1 _21200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11272_),
    .B(_11273_),
    .C(_11269_),
    .Y(_11274_)
);

NAND2X1 _19699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9628_),
    .B(_9623_),
    .Y(_9629_)
);

OAI21X1 _19279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8765_),
    .B(_9167_),
    .C(_8750_),
    .Y(_9168_)
);

FILL SFILL69080x30050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL48920x15050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _12727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8698_),
    .B(_9466_),
    .C(_11308_),
    .Y(_11318_)
);

AOI21X1 _12307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5091_),
    .B(_5278_),
    .C(_5310_),
    .Y(_6714_)
);

OR2X2 _22825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_984_),
    .B(_1144_),
    .Y(_1145_)
);

NOR3X1 _22405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_452_),
    .B(_449_),
    .C(_446_),
    .Y(_685_)
);

OAI21X1 _15199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4371_),
    .B(_4694_),
    .C(_4692_),
    .Y(_4695_)
);

NAND3X1 _16980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6644_),
    .B(_6645_),
    .C(_6646_),
    .Y(_6647_)
);

NAND3X1 _16560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6164_),
    .B(_6180_),
    .C(_6185_),
    .Y(_6186_)
);

INVX2 _16140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5669_),
    .Y(_5726_)
);

FILL SFILL3640x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _17765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7502_),
    .B(_7504_),
    .C(_7501_),
    .Y(_7508_)
);

NAND3X1 _17345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7039_),
    .B(_7033_),
    .C(_7037_),
    .Y(_7048_)
);

OAI21X1 _12480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519__bF$buf3),
    .B(_6044__bF$buf2),
    .C(_8599_),
    .Y(_8610_)
);

NAND3X1 _12060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3350_),
    .B(_3964_),
    .C(_3997_),
    .Y(_4008_)
);

FILL SFILL38920x13050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR3X1 _13685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2990_),
    .B(_3020_),
    .C(_3028_),
    .Y(_3038_)
);

AOI21X1 _13265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2488_),
    .B(_2494_),
    .C(_2423_),
    .Y(_2578_)
);

NAND2X1 _23783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2184_),
    .B(_2170_),
    .Y(_2188_)
);

NAND3X1 _23363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1730_),
    .B(_1731_),
    .C(_1728_),
    .Y(_1732_)
);

FILL SFILL3560x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9500_),
    .B(_9490_),
    .C(_9494_),
    .Y(_9862_)
);

NAND3X1 _15831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5381_),
    .B(_5386_),
    .C(_5384_),
    .Y(_5388_)
);

AOI21X1 _15411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4926_),
    .B(_4927_),
    .C(_4919_),
    .Y(_4929_)
);

FILL SFILL28840x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _20488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10476_),
    .B(_10480_),
    .C(_10482_),
    .Y(_10493_)
);

AOI21X1 _20068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9649_),
    .B(_9673_),
    .C(_9671_),
    .Y(_10032_)
);

FILL SFILL18920x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6239_),
    .B(_6233_),
    .C(_6237_),
    .Y(_6248_)
);

OAI21X1 _19088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8954_),
    .B(_8953_),
    .C(_8957_),
    .Y(_8958_)
);

OR2X2 _12956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_286_),
    .B(_1913_),
    .Y(_1914_)
);

OAI21X1 _12536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9203_),
    .B(_9214_),
    .C(_9192_),
    .Y(_9225_)
);

AOI21X1 _12116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4478_),
    .B(_4522_),
    .C(_4325_),
    .Y(_4621_)
);

NOR2X1 _22634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_904_),
    .B(_907_),
    .Y(_936_)
);

OAI21X1 _22214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_472_),
    .B(_476_),
    .C(_241_),
    .Y(_477_)
);

FILL SFILL18840x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _23839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .Y(_2247_)
);

NOR2X1 _23419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1790_),
    .B(_1791_),
    .Y(_1792_)
);

BUFX2 BUFX2_insert530 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465_),
    .Y(_2465__bF$buf0)
);

BUFX2 BUFX2_insert531 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf5)
);

BUFX2 BUFX2_insert532 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf4)
);

BUFX2 BUFX2_insert533 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf3)
);

OAI21X1 _17994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7757_),
    .B(_7758_),
    .C(_7753_),
    .Y(_7759_)
);

BUFX2 BUFX2_insert534 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf2)
);

OAI21X1 _17574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7289_),
    .B(_7290_),
    .C(_7287_),
    .Y(_7298_)
);

BUFX2 BUFX2_insert535 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf1)
);

BUFX2 BUFX2_insert536 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[30]),
    .Y(areg_30_bF$buf0)
);

NOR3X1 _17154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6817_),
    .B(_6832_),
    .C(_6837_),
    .Y(_6838_)
);

OAI21X1 _20700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10724_),
    .B(_10718_),
    .C(_10703_),
    .Y(_10725_)
);

AOI21X1 _18779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8618_),
    .B(_8617_),
    .C(_8609_),
    .Y(_8619_)
);

OAI21X1 _18359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8153_),
    .B(_8152_),
    .C(_8149_),
    .Y(_8159_)
);

AOI21X1 _13494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2822_),
    .B(_2823_),
    .C(_2821_),
    .Y(_2829_)
);

INVX1 _13074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2368_),
    .Y(_2369_)
);

OAI21X1 _23592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10684_),
    .B(_1974_),
    .C(_1980_),
    .Y(_1981_)
);

NAND3X1 _23172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .B(_1509_),
    .C(_1514_),
    .Y(_1524_)
);

OAI21X1 _19720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9295_),
    .B(_9285_),
    .C(_9289_),
    .Y(_9651_)
);

NAND2X1 _19300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9190_),
    .B(_9189_),
    .Y(_9191_)
);

FILL SFILL69080x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

OR2X2 _21905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11764_),
    .B(_131_),
    .Y(_138_)
);

NAND2X1 _14699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3838_),
    .B(_3848_),
    .Y(_4147_)
);

AOI21X1 _14279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3687_),
    .B(_3686_),
    .C(_3684_),
    .Y(_3688_)
);

FILL SFILL38600x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _15640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5173_),
    .B(_5177_),
    .Y(_5178_)
);

NAND3X1 _15220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4713_),
    .B(_4717_),
    .C(_4716_),
    .Y(_4718_)
);

FILL SFILL3640x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9935_),
    .B(_9933_),
    .C(_9942_),
    .Y(_10284_)
);

NAND3X1 _16845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6492_),
    .B(_6493_),
    .C(_6495_),
    .Y(_6499_)
);

OAI21X1 _16425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6035_),
    .B(_5298_),
    .C(_6037_),
    .Y(_6038_)
);

NOR3X1 _16005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5208_),
    .B(_5207_),
    .C(_5209_),
    .Y(_5579_)
);

NAND2X1 _11980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3131_),
    .B(_2486_),
    .Y(_3142_)
);

FILL SFILL69320x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL59000x21050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _12765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg_12_bF$buf3),
    .C(areg[0]),
    .D(breg_13_bF$buf0),
    .Y(_11734_)
);

NAND3X1 _12345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7043_),
    .B(_5859_),
    .C(_7020_),
    .Y(_7131_)
);

OAI21X1 _22863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1181_),
    .B(_1180_),
    .C(_1059_),
    .Y(_1187_)
);

INVX1 _22443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .Y(_727_)
);

NAND2X1 _22023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_18_bF$buf1),
    .B(breg_28_bF$buf1),
    .Y(_267_)
);

FILL SFILL33880x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _23648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2040_),
    .B(_2041_),
    .Y(_2042_)
);

OR2X2 _23228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1578_),
    .Y(_1583_)
);

OAI21X1 _14911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4374_),
    .B(_4378_),
    .C(_4369_),
    .Y(_4380_)
);

OAI21X1 _17383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7088_),
    .B(_7089_),
    .C(_7086_),
    .Y(_7090_)
);

FILL SFILL18920x49050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _18588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8001_),
    .B(_8003_),
    .C(_8409_),
    .Y(_8410_)
);

AOI21X1 _18168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7070_),
    .B(_7934_),
    .C(_7501_),
    .Y(_7950_)
);

FILL SFILL63960x44050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11826_),
    .B(_11821_),
    .C(_11716_),
    .Y(_11837_)
);

NAND3X1 _14088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3476_),
    .B(_3477_),
    .C(_3478_),
    .Y(_3479_)
);

NOR3X1 _22919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1235_),
    .B(_1233_),
    .C(_1230_),
    .Y(_1248_)
);

FILL SFILL8760x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _16654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6288_),
    .B(_6287_),
    .C(_6289_),
    .Y(_6290_)
);

OAI21X1 _16234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5829_),
    .B(_5824_),
    .C(_5746_),
    .Y(_5830_)
);

FILL SFILL53960x42050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7604_),
    .B(_7610_),
    .C(_7223_),
    .Y(_7611_)
);

AOI21X1 _17439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6677_),
    .B(_6727_),
    .C(_7150_),
    .Y(_7151_)
);

AND2X2 _17019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6683_),
    .B(_6684_),
    .Y(_6690_)
);

NAND3X1 _12994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2270_),
    .B(_2288_),
    .C(_2286_),
    .Y(_2289_)
);

NAND3X1 _12574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9598_),
    .B(_9631_),
    .C(_8500_),
    .Y(_9641_)
);

NAND2X1 _12154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf4),
    .B(breg_4_bF$buf5),
    .Y(_5036_)
);

NAND3X1 _22672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .B(_977_),
    .C(_975_),
    .Y(_978_)
);

OAI21X1 _22252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3402__bF$buf2),
    .B(_5668__bF$buf2),
    .C(_267_),
    .Y(_518_)
);

NAND2X1 _18800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8637_),
    .B(_8641_),
    .Y(_8642_)
);

OAI21X1 _13779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2888_),
    .B(_2878_),
    .C(_2883_),
    .Y(_3140_)
);

NOR3X1 _13359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2676_),
    .B(_2660_),
    .C(_2677_),
    .Y(_2681_)
);

XNOR2X1 _23877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3231_),
    .B(_3055_),
    .Y(_0_[1])
);

NAND3X1 _23457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1779_),
    .B(_1829_),
    .C(_1833_),
    .Y(_1834_)
);

FILL SFILL3720x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _23037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1371_),
    .B(_1364_),
    .C(_1368_),
    .Y(_1376_)
);

FILL SFILL74360x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4165_),
    .B(_4169_),
    .C(_4168_),
    .Y(_4170_)
);

NAND3X1 _14300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3704_),
    .B(_3705_),
    .C(_3669_),
    .Y(_3711_)
);

AOI21X1 _17192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6532_),
    .B(_6536_),
    .C(_6518_),
    .Y(_6880_)
);

FILL SFILL48840x7050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5485_),
    .B(_5490_),
    .C(_5471_),
    .Y(_5491_)
);

OAI21X1 _15505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5029_),
    .B(_5024_),
    .C(_5019_),
    .Y(_5030_)
);

FILL SFILL59080x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _18397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2465__bF$buf3),
    .B(_3529__bF$buf4),
    .C(_8200_),
    .Y(_8201_)
);

FILL SFILL59000x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _21943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_178_),
    .B(_11528_),
    .C(_179_),
    .Y(_180_)
);

OAI21X1 _21523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669__bF$buf2),
    .B(_5668__bF$buf5),
    .C(_11613_),
    .Y(_11628_)
);

OAI21X1 _21103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10879_),
    .B(_10877_),
    .C(_10868_),
    .Y(_11168_)
);

FILL SFILL33880x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

XOR2X1 _22728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_1038_),
    .Y(_1039_)
);

NAND3X1 _22308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_543_),
    .B(_574_),
    .C(_578_),
    .Y(_579_)
);

FILL SFILL49080x16050 (
    .gnd(gnd),
    .vdd(vdd)
);

XNOR2X1 _16883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6515_),
    .B(_6540_),
    .Y(_6541_)
);

AOI21X1 _16463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5748_),
    .B(_6078_),
    .C(_6077_),
    .Y(_6079_)
);

NAND3X1 _16043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5613_),
    .B(_5620_),
    .C(_5367_),
    .Y(_5621_)
);

FILL SFILL49000x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _17668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7380_),
    .B(_7395_),
    .C(_7400_),
    .Y(_7401_)
);

INVX2 _17248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6934_),
    .Y(_6941_)
);

NAND2X1 _12383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7492_),
    .B(_7536_),
    .Y(_7547_)
);

NAND3X1 _22481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_733_),
    .B(_766_),
    .C(_767_),
    .Y(_769_)
);

OAI21X1 _22061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3961__bF$buf3),
    .B(_5315__bF$buf1),
    .C(_302_),
    .Y(_309_)
);

FILL SFILL54280x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x14050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _13588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2909_),
    .B(_2918_),
    .C(_2920_),
    .Y(_2932_)
);

AOI21X1 _13168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2466_),
    .B(_2463_),
    .C(_2460_),
    .Y(_2472_)
);

XNOR2X1 _23686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2082_),
    .B(_2064_),
    .Y(_2083_)
);

FILL SFILL23800x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .B(_1623_),
    .C(_1625_),
    .Y(_1626_)
);

AOI21X1 _19814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9574_),
    .B(_9573_),
    .C(_9482_),
    .Y(_9755_)
);

FILL SFILL8840x40050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL44280x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _15734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5264_),
    .B(_5269_),
    .C(_4969_),
    .Y(_5282_)
);

NAND2X1 _15314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4820_),
    .B(_4821_),
    .Y(_4822_)
);

FILL SFILL53960x37050 (
    .gnd(gnd),
    .vdd(vdd)
);

BUFX2 BUFX2_insert60 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf2)
);

BUFX2 BUFX2_insert61 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf1)
);

BUFX2 BUFX2_insert62 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[15]),
    .Y(areg_15_bF$buf0)
);

BUFX2 BUFX2_insert63 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf5)
);

BUFX2 BUFX2_insert64 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf4)
);

BUFX2 BUFX2_insert65 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf3)
);

BUFX2 BUFX2_insert66 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf2)
);

BUFX2 BUFX2_insert67 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf1)
);

BUFX2 BUFX2_insert68 (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[25]),
    .Y(breg_25_bF$buf0)
);

BUFX2 BUFX2_insert69 (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6815_),
    .Y(_6815__bF$buf4)
);

OAI21X1 _16939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6359_),
    .B(_6601_),
    .C(_6349_),
    .Y(_6602_)
);

AND2X2 _16519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_19_bF$buf1),
    .Y(_6141_)
);

FILL SFILL74040x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _21752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10688_),
    .B(_11877_),
    .Y(_11878_)
);

NAND3X1 _21332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11411_),
    .B(_11418_),
    .C(_11368_),
    .Y(_11419_)
);

FILL SFILL29000x10050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL28680x2050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _12859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_144_),
    .B(_801_),
    .C(_845_),
    .Y(_856_)
);

AOI21X1 _12439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8073_),
    .B(_8008_),
    .C(_7283_),
    .Y(_8161_)
);

NAND2X1 _22957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1288_),
    .B(_1285_),
    .Y(_1289_)
);

FILL SFILL3720x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX2 _12019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3547_),
    .Y(_3558_)
);

AOI21X1 _22537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_826_),
    .B(_825_),
    .C(_824_),
    .Y(_830_)
);

NOR2X1 _22117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_368_),
    .Y(_369_)
);

FILL SFILL74360x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _13800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3156_),
    .B(_3163_),
    .C(_3139_),
    .Y(_3164_)
);

OAI21X1 _16692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6327_),
    .B(_6326_),
    .C(_6307_),
    .Y(_6332_)
);

OAI21X1 _16272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5529_),
    .B(_5535_),
    .C(_5537_),
    .Y(_5872_)
);

INVX2 _17897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7651_),
    .Y(_7652_)
);

AOI21X1 _17477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6509_),
    .B(_6770_),
    .C(_6775_),
    .Y(_7192_)
);

OAI21X1 _17057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6724_),
    .B(_6726_),
    .C(_6679_),
    .Y(_6732_)
);

INVX8 _12192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_6_bF$buf0),
    .Y(_5453_)
);

NAND3X1 _22290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_555_),
    .C(_558_),
    .Y(_559_)
);

OAI21X1 _20603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10612_),
    .B(_10613_),
    .C(_10608_),
    .Y(_10620_)
);

NOR3X1 _13397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2511_),
    .C(_2509_),
    .Y(_2723_)
);

AOI21X1 _23495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1820_),
    .B(_1802_),
    .C(_1874_),
    .Y(_1875_)
);

NAND2X1 _23075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_24_bF$buf0),
    .B(breg_28_bF$buf3),
    .Y(_1417_)
);

AOI21X1 _19623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9540_),
    .B(_9542_),
    .C(_9533_),
    .Y(_9546_)
);

OAI21X1 _19203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9082_),
    .B(_9078_),
    .C(_9083_),
    .Y(_9084_)
);

NAND2X1 _21808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_20_bF$buf4),
    .B(breg_24_bF$buf0),
    .Y(_31_)
);

NOR3X1 _15963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5532_),
    .B(_5527_),
    .C(_5531_),
    .Y(_5533_)
);

NAND3X1 _15543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5041_),
    .B(_5066_),
    .C(_5071_),
    .Y(_5072_)
);

NAND3X1 _15123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4359_),
    .B(_4606_),
    .C(_4612_),
    .Y(_4613_)
);

NOR3X1 _16748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5999_),
    .B(_6000_),
    .C(_5998_),
    .Y(_6393_)
);

NAND2X1 _16328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5558_),
    .B(_5932_),
    .Y(_5933_)
);

NAND3X1 _21981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11885_),
    .B(_215_),
    .C(_216_),
    .Y(_222_)
);

AOI21X1 _21561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11466_),
    .B(_11443_),
    .C(_11667_),
    .Y(_11669_)
);

FILL SFILL54280x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _21141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11207_),
    .B(_11208_),
    .C(_11206_),
    .Y(_11210_)
);

OAI21X1 _12668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10595_),
    .B(_10584_),
    .C(_10562_),
    .Y(_10671_)
);

INVX1 _12248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5585_),
    .Y(_6076_)
);

OAI21X1 _22766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1078_),
    .B(_1077_),
    .C(_1076_),
    .Y(_1081_)
);

INVX1 _22346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .Y(_621_)
);

INVX1 _16081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5658_),
    .Y(_5662_)
);

FILL SFILL13880x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _14814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4205_),
    .B(_4228_),
    .C(_4222_),
    .Y(_4274_)
);

OAI21X1 _17286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6979_),
    .B(_6980_),
    .C(_6982_),
    .Y(_6983_)
);

FILL SFILL13800x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10859_),
    .B(_10857_),
    .C(_10854_),
    .Y(_10871_)
);

NAND3X1 _20412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10401_),
    .B(_10405_),
    .C(_10409_),
    .Y(_10410_)
);

AND2X2 _19852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_15_bF$buf4),
    .B(areg_22_bF$buf3),
    .Y(_9797_)
);

NAND3X1 _19432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9328_),
    .B(_9332_),
    .C(_9335_),
    .Y(_9336_)
);

NAND2X1 _19012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8875_),
    .B(_8869_),
    .Y(_8876_)
);

OAI21X1 _11939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2398_),
    .B(_2419_),
    .C(_2672_),
    .Y(_2683_)
);

NOR2X1 _21617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11448_),
    .B(_11729_),
    .Y(_11730_)
);

OR2X2 _15772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4679_),
    .B(_5012_),
    .Y(_5323_)
);

NOR2X1 _15352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4545_),
    .B(_4863_),
    .Y(_4864_)
);

FILL SFILL64040x43050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _16977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6244_),
    .B(_6238_),
    .Y(_6644_)
);

NOR2X1 _16557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5468_),
    .B(_6177_),
    .Y(_6183_)
);

AOI21X1 _16137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5707_),
    .B(_5711_),
    .C(_5673_),
    .Y(_5723_)
);

NAND3X1 _21790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11904_),
    .B(_11895_),
    .C(_11908_),
    .Y(_11_)
);

AOI21X1 _21370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11147_),
    .B(_11149_),
    .C(_11156_),
    .Y(_11460_)
);

NAND2X1 _12897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1250_),
    .B(_1260_),
    .Y(_1271_)
);

INVX1 _12477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8566_),
    .Y(_8577_)
);

NAND3X1 _22995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(_1329_),
    .C(_1294_),
    .Y(_1330_)
);

NAND2X1 _12057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3942_),
    .B(_3909_),
    .Y(_3975_)
);

INVX1 _22575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_871_),
    .Y(_872_)
);

NAND3X1 _22155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .B(_409_),
    .C(_411_),
    .Y(_412_)
);

OAI21X1 _18703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8535_),
    .B(_8534_),
    .C(_8530_),
    .Y(_8536_)
);

FILL SFILL54040x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _19908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf2),
    .B(areg_25_bF$buf4),
    .Y(_9858_)
);

AOI21X1 _14623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4014_),
    .B(_4015_),
    .C(_3867_),
    .Y(_4064_)
);

AND2X2 _14203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_10_bF$buf0),
    .B(breg_10_bF$buf5),
    .Y(_3604_)
);

NAND2X1 _17095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6772_),
    .B(_6773_),
    .Y(_6774_)
);

NAND2X1 _15828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5382_),
    .B(_5383_),
    .Y(_5384_)
);

AOI21X1 _15408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4444_),
    .B(_4597_),
    .C(_4924_),
    .Y(_4925_)
);

XOR2X1 _20641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10337_),
    .B(_10660_),
    .Y(_0_[39])
);

AND2X2 _20221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9843_),
    .B(_9836_),
    .Y(_10201_)
);

NAND3X1 _19661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9581_),
    .B(_9582_),
    .C(_9580_),
    .Y(_9588_)
);

OAI21X1 _19241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9112_),
    .B(_9117_),
    .C(_9119_),
    .Y(_9127_)
);

FILL SFILL8920x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _21846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_62_),
    .B(_57_),
    .C(_27_),
    .Y(_73_)
);

NAND3X1 _21426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11519_),
    .B(_11521_),
    .C(_11520_),
    .Y(_11522_)
);

NAND2X1 _21006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_15_bF$buf4),
    .B(breg_26_bF$buf4),
    .Y(_11061_)
);

AND2X2 _15581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_16_bF$buf4),
    .Y(_5114_)
);

INVX2 _15161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4652_),
    .Y(_4654_)
);

FILL SFILL69160x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX1 _16786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6433_),
    .Y(_6434_)
);

NAND3X1 _16366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5968_),
    .B(_5884_),
    .C(_5974_),
    .Y(_5975_)
);

FILL SFILL74120x33050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_9_bF$buf1),
    .Y(_6483_)
);

AOI21X1 _22384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_399_),
    .B(_422_),
    .C(_431_),
    .Y(_663_)
);

NAND3X1 _18932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8779_),
    .B(_8374_),
    .C(_8777_),
    .Y(_8788_)
);

NOR3X1 _18512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8314_),
    .B(_8317_),
    .C(_8310_),
    .Y(_8328_)
);

FILL SFILL64520x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _23589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_917_),
    .B(_1976_),
    .C(_935_),
    .Y(_1977_)
);

OAI21X1 _23169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1519_),
    .B(_1515_),
    .C(_1406_),
    .Y(_1520_)
);

FILL SFILL64120x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _19717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9297_),
    .B(_9283_),
    .C(_9305_),
    .Y(_9648_)
);

NAND3X1 _14852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4063_),
    .B(_4309_),
    .C(_4315_),
    .Y(_4316_)
);

AOI21X1 _14432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3850_),
    .B(_3851_),
    .C(_3849_),
    .Y(_3856_)
);

OAI21X1 _14012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3161_),
    .B(_3141_),
    .C(_3151_),
    .Y(_3396_)
);

NAND3X1 _15637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5171_),
    .B(_5160_),
    .C(_5163_),
    .Y(_5175_)
);

AND2X2 _15217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_9_bF$buf3),
    .B(breg_15_bF$buf5),
    .Y(_4715_)
);

NAND2X1 _20870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_12_bF$buf0),
    .B(areg_28_bF$buf0),
    .Y(_10912_)
);

AOI21X1 _20450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10435_),
    .B(_10442_),
    .C(_10391_),
    .Y(_10451_)
);

NOR3X1 _20030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9961_),
    .B(_9964_),
    .C(_9966_),
    .Y(_9990_)
);

AOI21X1 _19890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9837_),
    .B(_9836_),
    .C(_9835_),
    .Y(_9838_)
);

AOI21X1 _19470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9372_),
    .B(_9373_),
    .C(_9371_),
    .Y(_9377_)
);

AOI21X1 _19050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8904_),
    .B(_8903_),
    .C(_8900_),
    .Y(_8916_)
);

NOR2X1 _11977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2376__bF$buf0),
    .Y(_3099_)
);

OAI21X1 _21655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2560__bF$buf3),
    .B(_7100__bF$buf0),
    .C(_11759_),
    .Y(_11772_)
);

AND2X2 _21235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11311_),
    .B(_11309_),
    .Y(_11312_)
);

FILL SFILL54040x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4903_),
    .B(_4904_),
    .C(_4902_),
    .Y(_4905_)
);

XNOR2X1 _13703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3057_),
    .B(_3052_),
    .Y(_3058_)
);

NAND2X1 _23801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2206_),
    .B(_2204_),
    .Y(_0_[59])
);

XNOR2X1 _16595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6224_),
    .B(_6222_),
    .Y(_6225_)
);

OAI21X1 _16175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5759_),
    .B(_5764_),
    .C(_5753_),
    .Y(_5765_)
);

OR2X2 _14908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4076_),
    .B(_4371_),
    .Y(_4376_)
);

FILL SFILL44040x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _12095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf3),
    .B(areg_7_bF$buf1),
    .Y(_4390_)
);

AOI21X1 _22193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_359_),
    .C(_250_),
    .Y(_454_)
);

AOI21X1 _18741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8576_),
    .B(_8575_),
    .C(_8568_),
    .Y(_8578_)
);

OAI21X1 _18321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8114_),
    .B(_8113_),
    .C(_8112_),
    .Y(_8118_)
);

AOI21X1 _20926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10625_),
    .B(_10627_),
    .C(_10973_),
    .Y(_10974_)
);

OAI22X1 _20506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9858_),
    .B(_10511_),
    .C(_10512_),
    .D(_10211_),
    .Y(_10513_)
);

FILL SFILL69640x52050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _23398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .B(_1654_),
    .Y(_1769_)
);

OAI21X1 _19946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9892_),
    .B(_9893_),
    .C(_9890_),
    .Y(_9899_)
);

NOR2X1 _19526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9059_),
    .B(_9100_),
    .Y(_9439_)
);

NAND3X1 _19106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8975_),
    .B(_8977_),
    .C(_8976_),
    .Y(_8978_)
);

NAND3X1 _14661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4100_),
    .B(_4104_),
    .C(_4103_),
    .Y(_4106_)
);

OAI22X1 _14241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf1),
    .B(_2287__bF$buf2),
    .C(_4116__bF$buf4),
    .D(_549__bF$buf4),
    .Y(_3647_)
);

FILL SFILL38760x54050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL69160x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL34040x32050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _15866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5055_),
    .B(_5106_),
    .Y(_5426_)
);

OAI21X1 _15446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4946_),
    .B(_4652_),
    .C(_4937_),
    .Y(_4965_)
);

OAI21X1 _15026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5453__bF$buf0),
    .B(_2884__bF$buf0),
    .C(_4498_),
    .Y(_4506_)
);

OAI21X1 _21884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_114_),
    .C(_103_),
    .Y(_115_)
);

OAI21X1 _21464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11562_),
    .B(_11563_),
    .C(_11438_),
    .Y(_11564_)
);

NAND3X1 _21044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11097_),
    .B(_11102_),
    .C(_11058_),
    .Y(_11103_)
);

FILL SFILL23800x4050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_973_),
    .B(_971_),
    .C(_953_),
    .Y(_974_)
);

FILL SFILL64120x26050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_513_),
    .B(_511_),
    .C(_509_),
    .Y(_514_)
);

NAND2X1 _13932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3308_),
    .B(_3304_),
    .Y(_3309_)
);

NAND2X1 _13512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf0),
    .B(areg_11_bF$buf1),
    .Y(_2849_)
);

OAI21X1 _23610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1916_),
    .B(_1917_),
    .C(_1999_),
    .Y(_2000_)
);

AND2X2 _14717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_9_bF$buf4),
    .B(areg_13_bF$buf0),
    .Y(_4167_)
);

NAND3X1 _17189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6859_),
    .B(_6872_),
    .C(_6862_),
    .Y(_6876_)
);

FILL SFILL18760x50050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x41050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _18970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8805_),
    .B(_8823_),
    .C(_8694_),
    .Y(_8829_)
);

NAND2X1 _18550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_4_bF$buf1),
    .B(areg_30_bF$buf3),
    .Y(_8369_)
);

AOI21X1 _18130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7900_),
    .B(_7907_),
    .C(_7886_),
    .Y(_7908_)
);

FILL SFILL54120x24050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _20735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10465_),
    .B(_10763_),
    .C(_10762_),
    .Y(_10764_)
);

OAI21X1 _20315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10302_),
    .B(_10303_),
    .C(_10301_),
    .Y(_10304_)
);

OAI21X1 _19755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9327_),
    .B(_9322_),
    .C(_9330_),
    .Y(_9690_)
);

NAND3X1 _19335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9223_),
    .B(_9224_),
    .C(_9222_),
    .Y(_9230_)
);

AOI21X1 _14890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4096_),
    .B(_4355_),
    .C(_4354_),
    .Y(_4356_)
);

NAND3X1 _14470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3889_),
    .B(_3874_),
    .C(_3892_),
    .Y(_3897_)
);

OAI21X1 _14050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3428_),
    .B(_3426_),
    .C(_3386_),
    .Y(_3437_)
);

FILL SFILL33960x6050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL18680x12050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND3X1 _15675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5216_),
    .B(_5181_),
    .C(_5211_),
    .Y(_5217_)
);

AOI21X1 _15255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4448_),
    .B(_4492_),
    .C(_4488_),
    .Y(_4757_)
);

FILL SFILL44040x29050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _21693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11528_),
    .B(_11813_),
    .Y(_11814_)
);

OAI21X1 _21273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11352_),
    .B(_11345_),
    .C(_11332_),
    .Y(_11353_)
);

AOI21X1 _17821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7564_),
    .B(_7563_),
    .C(_7562_),
    .Y(_7570_)
);

INVX2 _17401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7108_),
    .Y(_7110_)
);

AOI21X1 _22898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1224_),
    .C(_1072_),
    .Y(_1225_)
);

OAI21X1 _22478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_761_),
    .B(_764_),
    .C(_734_),
    .Y(_765_)
);

OAI21X1 _22058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_301_),
    .C(_299_),
    .Y(_305_)
);

NAND3X1 _18606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8174_),
    .B(_8180_),
    .C(_8178_),
    .Y(_8430_)
);

NAND2X1 _13741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .B(areg_10_bF$buf4),
    .Y(_3100_)
);

XOR2X1 _13321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2427_),
    .B(_2638_),
    .Y(_2640_)
);

FILL SFILL34040x27050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _14946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4416_),
    .B(_4417_),
    .C(_4415_),
    .Y(_4418_)
);

FILL SFILL29240x9050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_0_bF$buf1),
    .B(areg_21_bF$buf1),
    .Y(_3959_)
);

XOR2X1 _14106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3242_),
    .B(_3498_),
    .Y(_0_[19])
);

FILL SFILL69160x1050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL3800x53050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL8840x8050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10786_),
    .B(_10794_),
    .Y(_11015_)
);

FILL SFILL59240x31050 (
    .gnd(gnd),
    .vdd(vdd)
);

NAND2X1 _20544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10549_),
    .B(_10554_),
    .Y(_10555_)
);

NAND3X1 _20124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10084_),
    .B(_10077_),
    .C(_10082_),
    .Y(_10094_)
);

NAND3X1 _19984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9934_),
    .B(_9935_),
    .C(_9933_),
    .Y(_9941_)
);

NAND2X1 _19564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9475_),
    .B(_9480_),
    .Y(_9481_)
);

NAND2X1 _19144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9018_),
    .B(_9019_),
    .Y(_9020_)
);

FILL SFILL59160x38050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL24040x25050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI22X1 _21749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11584_),
    .B(_11589_),
    .C(_11859_),
    .D(_11864_),
    .Y(_11874_)
);

AOI21X1 _21329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11413_),
    .B(_11414_),
    .C(_11407_),
    .Y(_11415_)
);

NAND2X1 _15484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5002_),
    .B(_5006_),
    .Y(_5007_)
);

OAI21X1 _15064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4547_),
    .B(_4546_),
    .C(_4537_),
    .Y(_4548_)
);

FILL FILL74120x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _16689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6327_),
    .B(_6326_),
    .C(_6323_),
    .Y(_6328_)
);

OAI21X1 _16269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5863_),
    .B(_5864_),
    .C(_5846_),
    .Y(_5868_)
);

OAI21X1 _21082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3529__bF$buf3),
    .B(_4541__bF$buf4),
    .C(_11144_),
    .Y(_11145_)
);

FILL SFILL18760x45050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL49160x36050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL14040x23050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _17630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7357_),
    .B(_7358_),
    .Y(_7359_)
);

AOI21X1 _17210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6882_),
    .B(_6887_),
    .C(_6848_),
    .Y(_6899_)
);

FILL SFILL54120x19050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL39080x5050 (
    .gnd(gnd),
    .vdd(vdd)
);

FILL SFILL33960x20050 (
    .gnd(gnd),
    .vdd(vdd)
);

INVX8 _12189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(_5420_)
);

OAI21X1 _22287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3781__bF$buf0),
    .B(_5921__bF$buf3),
    .C(_311_),
    .Y(_556_)
);

OAI21X1 _18835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8674_),
    .B(_8679_),
    .C(_8680_),
    .Y(_8681_)
);

AOI21X1 _18415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8219_),
    .B(_8220_),
    .C(_8218_),
    .Y(_8221_)
);

NOR3X1 _13970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3346_),
    .B(_3348_),
    .C(_3347_),
    .Y(_3349_)
);

NAND3X1 _13550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2886_),
    .B(_2889_),
    .C(_2877_),
    .Y(_2890_)
);

XNOR2X1 _13130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2429_),
    .B(_2426_),
    .Y(_2430_)
);

FILL SFILL39160x34050 (
    .gnd(gnd),
    .vdd(vdd)
);

AND2X2 _14755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_7_bF$buf2),
    .B(areg_15_bF$buf1),
    .Y(_4209_)
);

NAND3X1 _14335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3746_),
    .B(_3747_),
    .C(_3522_),
    .Y(_3750_)
);

DFFPOSX1 _24013_ (
    .gnd(gnd),
    .vdd(vdd),
    .Q(areg[3]),
    .CLK(clk_bF$buf5),
    .D(a[3])
);

NAND3X1 _20773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10698_),
    .B(_10800_),
    .C(_10805_),
    .Y(_10806_)
);

NAND2X1 _20353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10097_),
    .B(_10292_),
    .Y(_10345_)
);

NAND2X1 _16901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg_13_bF$buf1),
    .B(areg_16_bF$buf4),
    .Y(_6561_)
);

OAI21X1 _19793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9720_),
    .B(_9719_),
    .C(_9716_),
    .Y(_9732_)
);

AOI21X1 _19373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9231_),
    .B(_9230_),
    .C(_8890_),
    .Y(_9271_)
);

OAI21X1 _21978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_217_),
    .C(_11884_),
    .Y(_218_)
);

AOI21X1 _21558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11659_),
    .B(_11658_),
    .C(_11656_),
    .Y(_11665_)
);

OR2X2 _21138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_11160_),
    .B(_11166_),
    .Y(_11206_)
);

FILL SFILL69240x28050 (
    .gnd(gnd),
    .vdd(vdd)
);

NOR2X1 _12821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_429_),
    .Y(_440_)
);

NOR2X1 _12401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6571_),
    .B(_7689_),
    .Y(_7744_)
);

NAND3X1 _15293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4798_),
    .B(_4797_),
    .C(_4795_),
    .Y(_4799_)
);

OAI21X1 _13606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2950_),
    .B(_2951_),
    .C(_2949_),
    .Y(_2952_)
);

NAND2X1 _23704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2056_),
    .B(_2102_),
    .Y(_2103_)
);

AOI21X1 _16498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_6109_),
    .B(_6102_),
    .C(_6054_),
    .Y(_6118_)
);

XNOR2X1 _16078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5302_),
    .B(_5658_),
    .Y(_0_[26])
);

FILL SFILL3800x48050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _22096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_345_),
    .B(_346_),
    .C(_344_),
    .Y(_347_)
);

AOI21X1 _18644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8470_),
    .B(_7652_),
    .C(_8469_),
    .Y(_8471_)
);

AOI21X1 _18224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8005_),
    .B(_8011_),
    .C(_7878_),
    .Y(_8012_)
);

OAI22X1 _20829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10212_),
    .B(_10865_),
    .C(_10866_),
    .D(_10557_),
    .Y(_10867_)
);

NAND2X1 _20409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_17_bF$buf2),
    .B(breg_22_bF$buf1),
    .Y(_10406_)
);

FILL FILL74200x11050 (
    .gnd(gnd),
    .vdd(vdd)
);

AOI21X1 _19849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9045_),
    .B(_9792_),
    .C(_9443_),
    .Y(_9793_)
);

NAND3X1 _19429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9329_),
    .B(_9331_),
    .C(_9330_),
    .Y(_9332_)
);

NAND3X1 _19009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8474_),
    .B(_8866_),
    .C(_8867_),
    .Y(_8872_)
);

NAND2X1 _14984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4457_),
    .B(_4458_),
    .Y(_4459_)
);

NAND3X1 _14564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_3994_),
    .B(_3993_),
    .C(_3995_),
    .Y(_4001_)
);

NAND2X1 _14144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_3_bF$buf0),
    .B(breg_17_bF$buf4),
    .Y(_3540_)
);

FILL FILL74120x18050 (
    .gnd(gnd),
    .vdd(vdd)
);

OAI21X1 _15769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_5318_),
    .C(_5313_),
    .Y(_5319_)
);

INVX2 _15349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4859_),
    .Y(_4860_)
);

AOI21X1 _20582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10594_),
    .B(_10590_),
    .C(_10596_),
    .Y(_10597_)
);

AOI21X1 _20162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10135_),
    .B(_10130_),
    .C(_10116_),
    .Y(_10136_)
);

AOI21X1 _16710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_5912_),
    .B(_5960_),
    .C(_6350_),
    .Y(_6351_)
);

OAI22X1 _19182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8286_),
    .B(_9059_),
    .C(_9061_),
    .D(_8696_),
    .Y(_9062_)
);

endmodule
