/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module multiplierCarry(
    input [7:0] a,
    input [7:0] b,
    input clk,
    output [15:0] y
);

wire [7:0] a ;
wire [7:0] b ;
wire [15:0] y ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _512_ ;
wire _321_ ;
wire _57_ ;
wire _130_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _127_ ;
wire _356_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire _488_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _115_ ;
wire _344_ ;
wire [7:0] \partialss[5]  ;
wire _153_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire _285_ ;
wire [15:0] _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire [15:0] _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire [14:0] psreg ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _141_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _176_ ;
wire _499_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _517_ ;
wire _270_ ;
wire _326_ ;
wire _135_ ;
wire _364_ ;
wire [7:0] \partialss[7]  ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _420_ ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _132_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire _493_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _167_ ;
wire _396_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire _126_ ;
wire _355_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire [7:0] breg ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _314_ ;
wire [7:0] \partialss[2]  ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire [7:0] areg ;
wire _311_ ;
wire _47_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire _308_ ;
wire _481_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire [6:0] _0_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _431_ ;
wire _240_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire [7:0] \partialss[4]  ;
wire _143_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire _140_ ;
wire _425_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _272_ ;
wire _328_ ;
wire _137_ ;
wire _366_ ;
wire _175_ ;
wire _269_ ;
wire _498_ ;
wire _26_ ;
wire _64_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _172_ ;
wire _228_ ;
wire _457_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire [7:0] \partialsb[0]  ;
wire _398_ ;
wire _513_ ;
wire _322_ ;
wire _58_ ;
wire _131_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire _454_ ;
wire _263_ ;
wire _319_ ;
wire _492_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire [7:0] \partialsco[7]  ;
wire _451_ ;
wire [7:0] \partialsb[7]  ;
wire _507_ ;
wire _260_ ;
wire _316_ ;
wire _125_ ;
wire _354_ ;
wire [7:0] \partialss[6]  ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _313_ ;
wire _49_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _116_ ;
wire _345_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire [7:0] \partialss[1]  ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _145_ ;
wire [7:0] pcreg ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _430_ ;
wire _524_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _142_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _177_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _518_ ;
wire _271_ ;
wire _327_ ;
wire _136_ ;
wire _365_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _421_ ;
wire _230_ ;
wire _515_ ;
wire _324_ ;
wire [7:0] \partialss[3]  ;
wire _133_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

CLKBUF1 CLKBUF1_insert6 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert5 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf6)
);

INVX1 _1000_ (
    .A(_210_),
    .Y(_419_)
);

NAND2X1 _1001_ (
    .A(_419_),
    .B(_181_),
    .Y(_420_)
);

XNOR2X1 _1002_ (
    .A(_420_),
    .B(_208_),
    .Y(\partialss[5] [0])
);

INVX1 _1003_ (
    .A(_176_),
    .Y(_421_)
);

NAND2X1 _1004_ (
    .A(_212_),
    .B(_421_),
    .Y(_422_)
);

XOR2X1 _1005_ (
    .A(_422_),
    .B(_211_),
    .Y(\partialss[6] [0])
);

INVX1 _1006_ (
    .A(_495_),
    .Y(_423_)
);

NAND3X1 _1007_ (
    .A(_499_),
    .B(_169_),
    .C(_170_),
    .Y(_424_)
);

OAI21X1 _1008_ (
    .A(_148_),
    .B(_167_),
    .C(_498_),
    .Y(_425_)
);

AOI21X1 _1009_ (
    .A(_424_),
    .B(_425_),
    .C(_423_),
    .Y(_426_)
);

OAI21X1 _1010_ (
    .A(_172_),
    .B(_426_),
    .C(_213_),
    .Y(_427_)
);

NAND3X1 _1011_ (
    .A(_423_),
    .B(_424_),
    .C(_425_),
    .Y(_428_)
);

NAND3X1 _1012_ (
    .A(_214_),
    .B(_428_),
    .C(_215_),
    .Y(_429_)
);

NAND2X1 _1013_ (
    .A(_429_),
    .B(_427_),
    .Y(\partialss[7] [0])
);

NAND2X1 _1014_ (
    .A(_266_),
    .B(_262_),
    .Y(_430_)
);

OAI21X1 _1015_ (
    .A(_430_),
    .B(_273_),
    .C(_270_),
    .Y(_431_)
);

OAI21X1 _1016_ (
    .A(_274_),
    .B(_268_),
    .C(_269_),
    .Y(_432_)
);

OAI21X1 _1017_ (
    .A(_268_),
    .B(_431_),
    .C(_432_),
    .Y(\partialss[7] [1])
);

NOR2X1 _1018_ (
    .A(_308_),
    .B(_279_),
    .Y(_433_)
);

OAI21X1 _1019_ (
    .A(_433_),
    .B(_365_),
    .C(_363_),
    .Y(_434_)
);

NAND2X1 _1020_ (
    .A(_308_),
    .B(_279_),
    .Y(_435_)
);

NAND3X1 _1021_ (
    .A(_362_),
    .B(_364_),
    .C(_435_),
    .Y(_436_)
);

INVX1 _1022_ (
    .A(_318_),
    .Y(_437_)
);

AOI21X1 _1023_ (
    .A(_436_),
    .B(_434_),
    .C(_437_),
    .Y(_438_)
);

OAI21X1 _1024_ (
    .A(_438_),
    .B(_319_),
    .C(_321_),
    .Y(_439_)
);

NAND3X1 _1025_ (
    .A(_436_),
    .B(_437_),
    .C(_434_),
    .Y(_440_)
);

NAND3X1 _1026_ (
    .A(_322_),
    .B(_323_),
    .C(_440_),
    .Y(_441_)
);

NAND2X1 _1027_ (
    .A(_441_),
    .B(_439_),
    .Y(\partialss[7] [2])
);

INVX1 _1028_ (
    .A(_366_),
    .Y(_442_)
);

AND2X2 _1029_ (
    .A(_357_),
    .B(_325_),
    .Y(_443_)
);

NOR2X1 _1030_ (
    .A(_325_),
    .B(_357_),
    .Y(_444_)
);

INVX1 _1031_ (
    .A(_360_),
    .Y(_445_)
);

NOR3X1 _1032_ (
    .A(_444_),
    .B(_445_),
    .C(_443_),
    .Y(_446_)
);

OAI21X1 _1033_ (
    .A(_446_),
    .B(_361_),
    .C(_442_),
    .Y(_447_)
);

OAI21X1 _1034_ (
    .A(_443_),
    .B(_444_),
    .C(_445_),
    .Y(_448_)
);

NAND3X1 _1035_ (
    .A(_366_),
    .B(_448_),
    .C(_367_),
    .Y(_449_)
);

NAND2X1 _1036_ (
    .A(_449_),
    .B(_447_),
    .Y(\partialss[7] [3])
);

NAND2X1 _1037_ (
    .A(_392_),
    .B(_387_),
    .Y(_450_)
);

XOR2X1 _1038_ (
    .A(_450_),
    .B(_390_),
    .Y(\partialss[7] [4])
);

XNOR2X1 _1039_ (
    .A(_401_),
    .B(_402_),
    .Y(_451_)
);

XOR2X1 _1040_ (
    .A(_451_),
    .B(_406_),
    .Y(\partialss[7] [5])
);

OR2X2 _1041_ (
    .A(\partialsco[7] [6]),
    .B(_413_),
    .Y(_452_)
);

AOI22X1 _1042_ (
    .A(_408_),
    .B(\partialsco[7] [6]),
    .C(_452_),
    .D(_412_),
    .Y(\partialss[7] [6])
);

NOR2X1 _1043_ (
    .A(_525_),
    .B(_485_),
    .Y(\partialsb[0] [0])
);

INVX1 _1044_ (
    .A(_199_),
    .Y(_453_)
);

NAND2X1 _1045_ (
    .A(_198_),
    .B(_453_),
    .Y(_454_)
);

XNOR2X1 _1046_ (
    .A(_454_),
    .B(_200_),
    .Y(\partialss[2] [0])
);

NAND2X1 _1047_ (
    .A(psreg[8]),
    .B(pcreg[0]),
    .Y(_455_)
);

INVX2 _1048_ (
    .A(_455_),
    .Y(_456_)
);

NOR2X1 _1049_ (
    .A(psreg[8]),
    .B(pcreg[0]),
    .Y(_457_)
);

NOR2X1 _1050_ (
    .A(_457_),
    .B(_456_),
    .Y(_1_[8])
);

NAND2X1 _1051_ (
    .A(psreg[9]),
    .B(pcreg[1]),
    .Y(_458_)
);

NOR2X1 _1052_ (
    .A(psreg[9]),
    .B(pcreg[1]),
    .Y(_459_)
);

INVX1 _1053_ (
    .A(_459_),
    .Y(_460_)
);

NAND2X1 _1054_ (
    .A(_458_),
    .B(_460_),
    .Y(_461_)
);

XNOR2X1 _1055_ (
    .A(_461_),
    .B(_456_),
    .Y(_1_[9])
);

AOI21X1 _1056_ (
    .A(_455_),
    .B(_458_),
    .C(_459_),
    .Y(_462_)
);

XNOR2X1 _1057_ (
    .A(psreg[10]),
    .B(pcreg[2]),
    .Y(_463_)
);

XNOR2X1 _1058_ (
    .A(_462_),
    .B(_463_),
    .Y(_1_[10])
);

INVX1 _1059_ (
    .A(psreg[11]),
    .Y(_464_)
);

NAND2X1 _1060_ (
    .A(psreg[10]),
    .B(_462_),
    .Y(_465_)
);

OAI21X1 _1061_ (
    .A(_462_),
    .B(psreg[10]),
    .C(pcreg[2]),
    .Y(_466_)
);

AND2X2 _1062_ (
    .A(_466_),
    .B(_465_),
    .Y(_467_)
);

NOR2X1 _1063_ (
    .A(_464_),
    .B(_467_),
    .Y(_468_)
);

NAND2X1 _1064_ (
    .A(pcreg[3]),
    .B(_468_),
    .Y(_469_)
);

NAND2X1 _1065_ (
    .A(_464_),
    .B(_467_),
    .Y(_470_)
);

OAI21X1 _1066_ (
    .A(_468_),
    .B(pcreg[3]),
    .C(_470_),
    .Y(_471_)
);

OAI21X1 _1067_ (
    .A(pcreg[3]),
    .B(_470_),
    .C(_471_),
    .Y(_472_)
);

NAND2X1 _1068_ (
    .A(_469_),
    .B(_472_),
    .Y(_1_[11])
);

INVX1 _1069_ (
    .A(pcreg[4]),
    .Y(_473_)
);

INVX1 _1070_ (
    .A(_471_),
    .Y(_474_)
);

NAND2X1 _1071_ (
    .A(psreg[12]),
    .B(_474_),
    .Y(_475_)
);

INVX1 _1072_ (
    .A(psreg[12]),
    .Y(_476_)
);

NAND2X1 _1073_ (
    .A(_476_),
    .B(_471_),
    .Y(_477_)
);

OAI21X1 _1074_ (
    .A(_471_),
    .B(_476_),
    .C(_473_),
    .Y(_478_)
);

OAI21X1 _1075_ (
    .A(psreg[12]),
    .B(_474_),
    .C(_478_),
    .Y(_479_)
);

OAI21X1 _1076_ (
    .A(pcreg[4]),
    .B(_477_),
    .C(_479_),
    .Y(_480_)
);

OAI21X1 _1077_ (
    .A(_473_),
    .B(_475_),
    .C(_480_),
    .Y(_1_[12])
);

INVX1 _1078_ (
    .A(pcreg[5]),
    .Y(_481_)
);

INVX1 _1079_ (
    .A(_479_),
    .Y(_482_)
);

NAND2X1 _1080_ (
    .A(psreg[13]),
    .B(_482_),
    .Y(_483_)
);

INVX1 _1081_ (
    .A(psreg[13]),
    .Y(_484_)
);

NAND2X1 _1082_ (
    .A(_484_),
    .B(_479_),
    .Y(_486_)
);

OAI21X1 _1083_ (
    .A(_479_),
    .B(_484_),
    .C(_481_),
    .Y(_487_)
);

OAI21X1 _1084_ (
    .A(psreg[13]),
    .B(_482_),
    .C(_487_),
    .Y(_488_)
);

OAI21X1 _1085_ (
    .A(pcreg[5]),
    .B(_486_),
    .C(_488_),
    .Y(_489_)
);

OAI21X1 _1086_ (
    .A(_481_),
    .B(_483_),
    .C(_489_),
    .Y(_1_[13])
);

XOR2X1 _1087_ (
    .A(psreg[14]),
    .B(pcreg[6]),
    .Y(_490_)
);

XNOR2X1 _1088_ (
    .A(_488_),
    .B(_490_),
    .Y(_1_[14])
);

INVX1 _1089_ (
    .A(psreg[14]),
    .Y(_491_)
);

INVX1 _1090_ (
    .A(_488_),
    .Y(_492_)
);

OAI21X1 _1091_ (
    .A(_492_),
    .B(psreg[14]),
    .C(pcreg[6]),
    .Y(_493_)
);

OAI21X1 _1092_ (
    .A(_491_),
    .B(_488_),
    .C(_493_),
    .Y(_0_[6])
);

BUFX2 _1093_ (
    .A(_532_[0]),
    .Y(y[0])
);

BUFX2 _1094_ (
    .A(_532_[1]),
    .Y(y[1])
);

BUFX2 _1095_ (
    .A(_532_[2]),
    .Y(y[2])
);

BUFX2 _1096_ (
    .A(_532_[3]),
    .Y(y[3])
);

BUFX2 _1097_ (
    .A(_532_[4]),
    .Y(y[4])
);

BUFX2 _1098_ (
    .A(_532_[5]),
    .Y(y[5])
);

BUFX2 _1099_ (
    .A(_532_[6]),
    .Y(y[6])
);

BUFX2 _1100_ (
    .A(_532_[7]),
    .Y(y[7])
);

BUFX2 _1101_ (
    .A(_532_[8]),
    .Y(y[8])
);

BUFX2 _1102_ (
    .A(_532_[9]),
    .Y(y[9])
);

BUFX2 _1103_ (
    .A(_532_[10]),
    .Y(y[10])
);

BUFX2 _1104_ (
    .A(_532_[11]),
    .Y(y[11])
);

BUFX2 _1105_ (
    .A(_532_[12]),
    .Y(y[12])
);

BUFX2 _1106_ (
    .A(_532_[13]),
    .Y(y[13])
);

BUFX2 _1107_ (
    .A(_532_[14]),
    .Y(y[14])
);

BUFX2 _1108_ (
    .A(_532_[15]),
    .Y(y[15])
);

DFFPOSX1 _1109_ (
    .CLK(clk_bF$buf6),
    .D(psreg[0]),
    .Q(_532_[0])
);

DFFPOSX1 _1110_ (
    .CLK(clk_bF$buf5),
    .D(psreg[1]),
    .Q(_532_[1])
);

DFFPOSX1 _1111_ (
    .CLK(clk_bF$buf4),
    .D(psreg[2]),
    .Q(_532_[2])
);

DFFPOSX1 _1112_ (
    .CLK(clk_bF$buf3),
    .D(psreg[3]),
    .Q(_532_[3])
);

DFFPOSX1 _1113_ (
    .CLK(clk_bF$buf2),
    .D(psreg[4]),
    .Q(_532_[4])
);

DFFPOSX1 _1114_ (
    .CLK(clk_bF$buf1),
    .D(psreg[5]),
    .Q(_532_[5])
);

DFFPOSX1 _1115_ (
    .CLK(clk_bF$buf0),
    .D(psreg[6]),
    .Q(_532_[6])
);

DFFPOSX1 _1116_ (
    .CLK(clk_bF$buf6),
    .D(psreg[7]),
    .Q(_532_[7])
);

DFFPOSX1 _1117_ (
    .CLK(clk_bF$buf5),
    .D(_1_[8]),
    .Q(_532_[8])
);

DFFPOSX1 _1118_ (
    .CLK(clk_bF$buf4),
    .D(_1_[9]),
    .Q(_532_[9])
);

DFFPOSX1 _1119_ (
    .CLK(clk_bF$buf3),
    .D(_1_[10]),
    .Q(_532_[10])
);

DFFPOSX1 _1120_ (
    .CLK(clk_bF$buf2),
    .D(_1_[11]),
    .Q(_532_[11])
);

DFFPOSX1 _1121_ (
    .CLK(clk_bF$buf1),
    .D(_1_[12]),
    .Q(_532_[12])
);

DFFPOSX1 _1122_ (
    .CLK(clk_bF$buf0),
    .D(_1_[13]),
    .Q(_532_[13])
);

DFFPOSX1 _1123_ (
    .CLK(clk_bF$buf6),
    .D(_1_[14]),
    .Q(_532_[14])
);

DFFPOSX1 _1124_ (
    .CLK(clk_bF$buf5),
    .D(_0_[6]),
    .Q(_532_[15])
);

DFFPOSX1 _1125_ (
    .CLK(clk_bF$buf4),
    .D(\partialsb[0] [0]),
    .Q(psreg[0])
);

DFFPOSX1 _1126_ (
    .CLK(clk_bF$buf3),
    .D(\partialss[1] [0]),
    .Q(psreg[1])
);

DFFPOSX1 _1127_ (
    .CLK(clk_bF$buf2),
    .D(\partialss[2] [0]),
    .Q(psreg[2])
);

DFFPOSX1 _1128_ (
    .CLK(clk_bF$buf1),
    .D(\partialss[3] [0]),
    .Q(psreg[3])
);

DFFPOSX1 _1129_ (
    .CLK(clk_bF$buf0),
    .D(\partialss[4] [0]),
    .Q(psreg[4])
);

DFFPOSX1 _1130_ (
    .CLK(clk_bF$buf6),
    .D(\partialss[5] [0]),
    .Q(psreg[5])
);

DFFPOSX1 _1131_ (
    .CLK(clk_bF$buf5),
    .D(\partialss[6] [0]),
    .Q(psreg[6])
);

DFFPOSX1 _1132_ (
    .CLK(clk_bF$buf4),
    .D(\partialss[7] [0]),
    .Q(psreg[7])
);

DFFPOSX1 _1133_ (
    .CLK(clk_bF$buf3),
    .D(\partialss[7] [1]),
    .Q(psreg[8])
);

DFFPOSX1 _1134_ (
    .CLK(clk_bF$buf2),
    .D(\partialss[7] [2]),
    .Q(psreg[9])
);

DFFPOSX1 _1135_ (
    .CLK(clk_bF$buf1),
    .D(\partialss[7] [3]),
    .Q(psreg[10])
);

DFFPOSX1 _1136_ (
    .CLK(clk_bF$buf0),
    .D(\partialss[7] [4]),
    .Q(psreg[11])
);

DFFPOSX1 _1137_ (
    .CLK(clk_bF$buf6),
    .D(\partialss[7] [5]),
    .Q(psreg[12])
);

DFFPOSX1 _1138_ (
    .CLK(clk_bF$buf5),
    .D(\partialss[7] [6]),
    .Q(psreg[13])
);

DFFPOSX1 _1139_ (
    .CLK(clk_bF$buf4),
    .D(\partialsb[7] [7]),
    .Q(psreg[14])
);

DFFPOSX1 _1140_ (
    .CLK(clk_bF$buf3),
    .D(\partialsco[7] [0]),
    .Q(pcreg[0])
);

DFFPOSX1 _1141_ (
    .CLK(clk_bF$buf2),
    .D(\partialsco[7] [1]),
    .Q(pcreg[1])
);

DFFPOSX1 _1142_ (
    .CLK(clk_bF$buf1),
    .D(\partialsco[7] [2]),
    .Q(pcreg[2])
);

DFFPOSX1 _1143_ (
    .CLK(clk_bF$buf0),
    .D(\partialsco[7] [3]),
    .Q(pcreg[3])
);

DFFPOSX1 _1144_ (
    .CLK(clk_bF$buf6),
    .D(\partialsco[7] [4]),
    .Q(pcreg[4])
);

DFFPOSX1 _1145_ (
    .CLK(clk_bF$buf5),
    .D(\partialsco[7] [5]),
    .Q(pcreg[5])
);

DFFPOSX1 _1146_ (
    .CLK(clk_bF$buf4),
    .D(\partialsco[7] [6]),
    .Q(pcreg[6])
);

DFFPOSX1 _1147_ (
    .CLK(clk_bF$buf3),
    .D(a[0]),
    .Q(areg[0])
);

DFFPOSX1 _1148_ (
    .CLK(clk_bF$buf2),
    .D(a[1]),
    .Q(areg[1])
);

DFFPOSX1 _1149_ (
    .CLK(clk_bF$buf1),
    .D(a[2]),
    .Q(areg[2])
);

DFFPOSX1 _1150_ (
    .CLK(clk_bF$buf0),
    .D(a[3]),
    .Q(areg[3])
);

DFFPOSX1 _1151_ (
    .CLK(clk_bF$buf6),
    .D(a[4]),
    .Q(areg[4])
);

DFFPOSX1 _1152_ (
    .CLK(clk_bF$buf5),
    .D(a[5]),
    .Q(areg[5])
);

DFFPOSX1 _1153_ (
    .CLK(clk_bF$buf4),
    .D(a[6]),
    .Q(areg[6])
);

DFFPOSX1 _1154_ (
    .CLK(clk_bF$buf3),
    .D(a[7]),
    .Q(areg[7])
);

DFFPOSX1 _1155_ (
    .CLK(clk_bF$buf2),
    .D(b[0]),
    .Q(breg[0])
);

DFFPOSX1 _1156_ (
    .CLK(clk_bF$buf1),
    .D(b[1]),
    .Q(breg[1])
);

DFFPOSX1 _1157_ (
    .CLK(clk_bF$buf0),
    .D(b[2]),
    .Q(breg[2])
);

DFFPOSX1 _1158_ (
    .CLK(clk_bF$buf6),
    .D(b[3]),
    .Q(breg[3])
);

DFFPOSX1 _1159_ (
    .CLK(clk_bF$buf5),
    .D(b[4]),
    .Q(breg[4])
);

DFFPOSX1 _1160_ (
    .CLK(clk_bF$buf4),
    .D(b[5]),
    .Q(breg[5])
);

DFFPOSX1 _1161_ (
    .CLK(clk_bF$buf3),
    .D(b[6]),
    .Q(breg[6])
);

DFFPOSX1 _1162_ (
    .CLK(clk_bF$buf2),
    .D(b[7]),
    .Q(breg[7])
);

INVX4 _533_ (
    .A(breg[0]),
    .Y(_485_)
);

INVX4 _534_ (
    .A(areg[7]),
    .Y(_494_)
);

NOR2X1 _535_ (
    .A(_485_),
    .B(_494_),
    .Y(_495_)
);

INVX4 _536_ (
    .A(areg[6]),
    .Y(_496_)
);

INVX4 _537_ (
    .A(breg[1]),
    .Y(_497_)
);

NOR2X1 _538_ (
    .A(_496_),
    .B(_497_),
    .Y(_498_)
);

INVX2 _539_ (
    .A(_498_),
    .Y(_499_)
);

NAND2X1 _540_ (
    .A(breg[2]),
    .B(areg[2]),
    .Y(_500_)
);

NAND2X1 _541_ (
    .A(breg[3]),
    .B(areg[0]),
    .Y(_501_)
);

NAND2X1 _542_ (
    .A(breg[2]),
    .B(areg[1]),
    .Y(_502_)
);

NOR2X1 _543_ (
    .A(_501_),
    .B(_502_),
    .Y(_503_)
);

AND2X2 _544_ (
    .A(breg[3]),
    .B(areg[0]),
    .Y(_504_)
);

AND2X2 _545_ (
    .A(areg[1]),
    .B(breg[4]),
    .Y(_505_)
);

NAND2X1 _546_ (
    .A(_504_),
    .B(_505_),
    .Y(_506_)
);

INVX4 _547_ (
    .A(breg[3]),
    .Y(_507_)
);

INVX2 _548_ (
    .A(areg[1]),
    .Y(_508_)
);

NAND2X1 _549_ (
    .A(areg[0]),
    .B(breg[4]),
    .Y(_509_)
);

OAI21X1 _550_ (
    .A(_507_),
    .B(_508_),
    .C(_509_),
    .Y(_510_)
);

AOI21X1 _551_ (
    .A(_510_),
    .B(_506_),
    .C(_503_),
    .Y(_511_)
);

AND2X2 _552_ (
    .A(breg[3]),
    .B(areg[1]),
    .Y(_512_)
);

NAND2X1 _553_ (
    .A(breg[2]),
    .B(areg[0]),
    .Y(_513_)
);

INVX1 _554_ (
    .A(_513_),
    .Y(_514_)
);

NAND3X1 _555_ (
    .A(_509_),
    .B(_512_),
    .C(_514_),
    .Y(_515_)
);

INVX1 _556_ (
    .A(_515_),
    .Y(_516_)
);

OAI21X1 _557_ (
    .A(_516_),
    .B(_511_),
    .C(_500_),
    .Y(_517_)
);

INVX1 _558_ (
    .A(_500_),
    .Y(_518_)
);

INVX1 _559_ (
    .A(_512_),
    .Y(_519_)
);

NAND2X1 _560_ (
    .A(areg[1]),
    .B(breg[4]),
    .Y(_520_)
);

OAI21X1 _561_ (
    .A(_501_),
    .B(_520_),
    .C(_510_),
    .Y(_521_)
);

OAI21X1 _562_ (
    .A(_519_),
    .B(_513_),
    .C(_521_),
    .Y(_522_)
);

NAND3X1 _563_ (
    .A(_518_),
    .B(_515_),
    .C(_522_),
    .Y(_523_)
);

INVX2 _564_ (
    .A(_502_),
    .Y(_524_)
);

INVX2 _565_ (
    .A(areg[0]),
    .Y(_525_)
);

NOR2X1 _566_ (
    .A(_525_),
    .B(_497_),
    .Y(_526_)
);

NAND2X1 _567_ (
    .A(_524_),
    .B(_526_),
    .Y(_527_)
);

NOR2X1 _568_ (
    .A(_504_),
    .B(_524_),
    .Y(_528_)
);

OAI21X1 _569_ (
    .A(_528_),
    .B(_503_),
    .C(_527_),
    .Y(_529_)
);

INVX4 _570_ (
    .A(areg[2]),
    .Y(_530_)
);

NAND3X1 _571_ (
    .A(_501_),
    .B(_524_),
    .C(_526_),
    .Y(_531_)
);

OAI21X1 _572_ (
    .A(_530_),
    .B(_497_),
    .C(_531_),
    .Y(_2_)
);

AND2X2 _573_ (
    .A(_529_),
    .B(_2_),
    .Y(_3_)
);

NAND3X1 _574_ (
    .A(_517_),
    .B(_523_),
    .C(_3_),
    .Y(_4_)
);

AOI21X1 _575_ (
    .A(_517_),
    .B(_523_),
    .C(_3_),
    .Y(_5_)
);

INVX4 _576_ (
    .A(areg[3]),
    .Y(_6_)
);

NOR2X1 _577_ (
    .A(_6_),
    .B(_497_),
    .Y(_7_)
);

INVX1 _578_ (
    .A(_7_),
    .Y(_8_)
);

OAI21X1 _579_ (
    .A(_5_),
    .B(_8_),
    .C(_4_),
    .Y(_9_)
);

INVX4 _580_ (
    .A(breg[2]),
    .Y(_10_)
);

NOR2X1 _581_ (
    .A(_6_),
    .B(_10_),
    .Y(_11_)
);

INVX2 _582_ (
    .A(_11_),
    .Y(_12_)
);

OAI21X1 _583_ (
    .A(_511_),
    .B(_500_),
    .C(_515_),
    .Y(_13_)
);

NOR2X1 _584_ (
    .A(_507_),
    .B(_530_),
    .Y(_14_)
);

INVX2 _585_ (
    .A(_14_),
    .Y(_15_)
);

INVX1 _586_ (
    .A(_509_),
    .Y(_16_)
);

AND2X2 _587_ (
    .A(areg[0]),
    .B(breg[5]),
    .Y(_17_)
);

NAND2X1 _588_ (
    .A(_505_),
    .B(_17_),
    .Y(_18_)
);

INVX4 _589_ (
    .A(breg[4]),
    .Y(_19_)
);

NAND2X1 _590_ (
    .A(areg[0]),
    .B(breg[5]),
    .Y(_20_)
);

OAI21X1 _591_ (
    .A(_508_),
    .B(_19_),
    .C(_20_),
    .Y(_21_)
);

AOI22X1 _592_ (
    .A(_512_),
    .B(_16_),
    .C(_18_),
    .D(_21_),
    .Y(_22_)
);

NAND3X1 _593_ (
    .A(_20_),
    .B(_504_),
    .C(_505_),
    .Y(_23_)
);

INVX1 _594_ (
    .A(_23_),
    .Y(_24_)
);

OAI21X1 _595_ (
    .A(_22_),
    .B(_24_),
    .C(_15_),
    .Y(_25_)
);

NOR2X1 _596_ (
    .A(_520_),
    .B(_20_),
    .Y(_26_)
);

NOR2X1 _597_ (
    .A(_505_),
    .B(_17_),
    .Y(_27_)
);

OAI21X1 _598_ (
    .A(_27_),
    .B(_26_),
    .C(_506_),
    .Y(_28_)
);

NAND3X1 _599_ (
    .A(_14_),
    .B(_23_),
    .C(_28_),
    .Y(_29_)
);

AOI21X1 _600_ (
    .A(_25_),
    .B(_29_),
    .C(_13_),
    .Y(_30_)
);

OAI21X1 _601_ (
    .A(_10_),
    .B(_530_),
    .C(_515_),
    .Y(_31_)
);

NAND2X1 _602_ (
    .A(_31_),
    .B(_522_),
    .Y(_32_)
);

NAND3X1 _603_ (
    .A(_15_),
    .B(_23_),
    .C(_28_),
    .Y(_33_)
);

OAI21X1 _604_ (
    .A(_22_),
    .B(_24_),
    .C(_14_),
    .Y(_34_)
);

AOI21X1 _605_ (
    .A(_34_),
    .B(_33_),
    .C(_32_),
    .Y(_35_)
);

OAI21X1 _606_ (
    .A(_35_),
    .B(_30_),
    .C(_12_),
    .Y(_36_)
);

NAND3X1 _607_ (
    .A(_33_),
    .B(_34_),
    .C(_32_),
    .Y(_37_)
);

NAND3X1 _608_ (
    .A(_13_),
    .B(_25_),
    .C(_29_),
    .Y(_38_)
);

NAND3X1 _609_ (
    .A(_11_),
    .B(_38_),
    .C(_37_),
    .Y(_39_)
);

NAND3X1 _610_ (
    .A(_36_),
    .B(_39_),
    .C(_9_),
    .Y(_40_)
);

AOI21X1 _611_ (
    .A(_36_),
    .B(_39_),
    .C(_9_),
    .Y(_41_)
);

INVX4 _612_ (
    .A(areg[4]),
    .Y(_42_)
);

NOR2X1 _613_ (
    .A(_42_),
    .B(_497_),
    .Y(_43_)
);

INVX1 _614_ (
    .A(_43_),
    .Y(_44_)
);

OAI21X1 _615_ (
    .A(_41_),
    .B(_44_),
    .C(_40_),
    .Y(_45_)
);

NOR2X1 _616_ (
    .A(_10_),
    .B(_42_),
    .Y(_46_)
);

INVX2 _617_ (
    .A(_46_),
    .Y(_47_)
);

OAI21X1 _618_ (
    .A(_30_),
    .B(_12_),
    .C(_38_),
    .Y(_48_)
);

NOR2X1 _619_ (
    .A(_6_),
    .B(_507_),
    .Y(_49_)
);

INVX2 _620_ (
    .A(_49_),
    .Y(_50_)
);

OAI21X1 _621_ (
    .A(_22_),
    .B(_15_),
    .C(_23_),
    .Y(_51_)
);

NOR2X1 _622_ (
    .A(_530_),
    .B(_19_),
    .Y(_52_)
);

INVX2 _623_ (
    .A(_52_),
    .Y(_53_)
);

AND2X2 _624_ (
    .A(areg[1]),
    .B(breg[5]),
    .Y(_54_)
);

AND2X2 _625_ (
    .A(areg[0]),
    .B(breg[6]),
    .Y(_55_)
);

NAND2X1 _626_ (
    .A(_54_),
    .B(_55_),
    .Y(_56_)
);

INVX4 _627_ (
    .A(breg[5]),
    .Y(_57_)
);

NAND2X1 _628_ (
    .A(areg[0]),
    .B(breg[6]),
    .Y(_58_)
);

OAI21X1 _629_ (
    .A(_508_),
    .B(_57_),
    .C(_58_),
    .Y(_59_)
);

AOI21X1 _630_ (
    .A(_59_),
    .B(_56_),
    .C(_26_),
    .Y(_60_)
);

NAND3X1 _631_ (
    .A(_54_),
    .B(_58_),
    .C(_16_),
    .Y(_61_)
);

INVX2 _632_ (
    .A(_61_),
    .Y(_62_)
);

OAI21X1 _633_ (
    .A(_62_),
    .B(_60_),
    .C(_53_),
    .Y(_63_)
);

NAND2X1 _634_ (
    .A(areg[1]),
    .B(breg[5]),
    .Y(_64_)
);

NOR2X1 _635_ (
    .A(_64_),
    .B(_58_),
    .Y(_65_)
);

AND2X2 _636_ (
    .A(_64_),
    .B(_58_),
    .Y(_66_)
);

OAI21X1 _637_ (
    .A(_66_),
    .B(_65_),
    .C(_18_),
    .Y(_67_)
);

NAND3X1 _638_ (
    .A(_52_),
    .B(_61_),
    .C(_67_),
    .Y(_68_)
);

AOI21X1 _639_ (
    .A(_68_),
    .B(_63_),
    .C(_51_),
    .Y(_69_)
);

OAI21X1 _640_ (
    .A(_507_),
    .B(_530_),
    .C(_23_),
    .Y(_70_)
);

NAND2X1 _641_ (
    .A(_70_),
    .B(_28_),
    .Y(_71_)
);

NAND3X1 _642_ (
    .A(_53_),
    .B(_61_),
    .C(_67_),
    .Y(_72_)
);

OAI21X1 _643_ (
    .A(_62_),
    .B(_60_),
    .C(_52_),
    .Y(_73_)
);

AOI21X1 _644_ (
    .A(_72_),
    .B(_73_),
    .C(_71_),
    .Y(_74_)
);

OAI21X1 _645_ (
    .A(_69_),
    .B(_74_),
    .C(_50_),
    .Y(_75_)
);

NAND3X1 _646_ (
    .A(_71_),
    .B(_72_),
    .C(_73_),
    .Y(_76_)
);

NAND3X1 _647_ (
    .A(_51_),
    .B(_68_),
    .C(_63_),
    .Y(_77_)
);

NAND3X1 _648_ (
    .A(_49_),
    .B(_76_),
    .C(_77_),
    .Y(_78_)
);

AOI21X1 _649_ (
    .A(_78_),
    .B(_75_),
    .C(_48_),
    .Y(_79_)
);

AOI21X1 _650_ (
    .A(_11_),
    .B(_37_),
    .C(_35_),
    .Y(_80_)
);

NAND3X1 _651_ (
    .A(_50_),
    .B(_76_),
    .C(_77_),
    .Y(_81_)
);

OAI21X1 _652_ (
    .A(_69_),
    .B(_74_),
    .C(_49_),
    .Y(_82_)
);

AOI21X1 _653_ (
    .A(_81_),
    .B(_82_),
    .C(_80_),
    .Y(_83_)
);

OAI21X1 _654_ (
    .A(_79_),
    .B(_83_),
    .C(_47_),
    .Y(_84_)
);

NAND3X1 _655_ (
    .A(_81_),
    .B(_80_),
    .C(_82_),
    .Y(_85_)
);

NAND3X1 _656_ (
    .A(_48_),
    .B(_78_),
    .C(_75_),
    .Y(_86_)
);

NAND3X1 _657_ (
    .A(_46_),
    .B(_86_),
    .C(_85_),
    .Y(_87_)
);

NAND3X1 _658_ (
    .A(_87_),
    .B(_84_),
    .C(_45_),
    .Y(_88_)
);

AOI21X1 _659_ (
    .A(_87_),
    .B(_84_),
    .C(_45_),
    .Y(_89_)
);

INVX4 _660_ (
    .A(areg[5]),
    .Y(_90_)
);

NOR2X1 _661_ (
    .A(_90_),
    .B(_497_),
    .Y(_91_)
);

INVX1 _662_ (
    .A(_91_),
    .Y(_92_)
);

OAI21X1 _663_ (
    .A(_89_),
    .B(_92_),
    .C(_88_),
    .Y(_93_)
);

NOR2X1 _664_ (
    .A(_90_),
    .B(_10_),
    .Y(_94_)
);

INVX2 _665_ (
    .A(_94_),
    .Y(_95_)
);

OAI21X1 _666_ (
    .A(_79_),
    .B(_47_),
    .C(_86_),
    .Y(_96_)
);

NOR2X1 _667_ (
    .A(_507_),
    .B(_42_),
    .Y(_97_)
);

INVX1 _668_ (
    .A(_97_),
    .Y(_98_)
);

OAI21X1 _669_ (
    .A(_69_),
    .B(_50_),
    .C(_77_),
    .Y(_99_)
);

NOR2X1 _670_ (
    .A(_6_),
    .B(_19_),
    .Y(_100_)
);

INVX2 _671_ (
    .A(_100_),
    .Y(_101_)
);

OAI21X1 _672_ (
    .A(_60_),
    .B(_53_),
    .C(_61_),
    .Y(_102_)
);

NOR2X1 _673_ (
    .A(_530_),
    .B(_57_),
    .Y(_103_)
);

INVX2 _674_ (
    .A(_103_),
    .Y(_104_)
);

AND2X2 _675_ (
    .A(areg[1]),
    .B(breg[7]),
    .Y(_105_)
);

NAND2X1 _676_ (
    .A(_55_),
    .B(_105_),
    .Y(_106_)
);

INVX2 _677_ (
    .A(breg[7]),
    .Y(_107_)
);

NAND2X1 _678_ (
    .A(areg[1]),
    .B(breg[6]),
    .Y(_108_)
);

OAI21X1 _679_ (
    .A(_525_),
    .B(_107_),
    .C(_108_),
    .Y(_109_)
);

AOI21X1 _680_ (
    .A(_109_),
    .B(_106_),
    .C(_65_),
    .Y(_110_)
);

NAND2X1 _681_ (
    .A(areg[0]),
    .B(breg[7]),
    .Y(_111_)
);

INVX1 _682_ (
    .A(_111_),
    .Y(_112_)
);

NOR3X1 _683_ (
    .A(_20_),
    .B(_108_),
    .C(_112_),
    .Y(_113_)
);

OAI21X1 _684_ (
    .A(_110_),
    .B(_113_),
    .C(_104_),
    .Y(_114_)
);

NAND2X1 _685_ (
    .A(areg[1]),
    .B(breg[7]),
    .Y(_115_)
);

NOR2X1 _686_ (
    .A(_58_),
    .B(_115_),
    .Y(_116_)
);

AND2X2 _687_ (
    .A(_108_),
    .B(_111_),
    .Y(_117_)
);

OAI21X1 _688_ (
    .A(_117_),
    .B(_116_),
    .C(_56_),
    .Y(_118_)
);

NAND3X1 _689_ (
    .A(_65_),
    .B(_109_),
    .C(_106_),
    .Y(_119_)
);

NAND3X1 _690_ (
    .A(_103_),
    .B(_119_),
    .C(_118_),
    .Y(_120_)
);

AOI21X1 _691_ (
    .A(_120_),
    .B(_114_),
    .C(_102_),
    .Y(_121_)
);

AOI21X1 _692_ (
    .A(_52_),
    .B(_67_),
    .C(_62_),
    .Y(_122_)
);

NAND3X1 _693_ (
    .A(_104_),
    .B(_119_),
    .C(_118_),
    .Y(_123_)
);

OAI21X1 _694_ (
    .A(_110_),
    .B(_113_),
    .C(_103_),
    .Y(_124_)
);

AOI21X1 _695_ (
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_125_)
);

OAI21X1 _696_ (
    .A(_121_),
    .B(_125_),
    .C(_101_),
    .Y(_126_)
);

NAND3X1 _697_ (
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_127_)
);

NAND3X1 _698_ (
    .A(_120_),
    .B(_102_),
    .C(_114_),
    .Y(_128_)
);

NAND3X1 _699_ (
    .A(_100_),
    .B(_127_),
    .C(_128_),
    .Y(_129_)
);

AOI21X1 _700_ (
    .A(_129_),
    .B(_126_),
    .C(_99_),
    .Y(_130_)
);

AOI21X1 _701_ (
    .A(_49_),
    .B(_76_),
    .C(_74_),
    .Y(_131_)
);

NAND3X1 _702_ (
    .A(_101_),
    .B(_127_),
    .C(_128_),
    .Y(_132_)
);

OAI21X1 _703_ (
    .A(_121_),
    .B(_125_),
    .C(_100_),
    .Y(_133_)
);

AOI21X1 _704_ (
    .A(_132_),
    .B(_133_),
    .C(_131_),
    .Y(_134_)
);

OAI21X1 _705_ (
    .A(_130_),
    .B(_134_),
    .C(_98_),
    .Y(_135_)
);

NAND3X1 _706_ (
    .A(_132_),
    .B(_133_),
    .C(_131_),
    .Y(_136_)
);

NAND3X1 _707_ (
    .A(_129_),
    .B(_126_),
    .C(_99_),
    .Y(_137_)
);

NAND3X1 _708_ (
    .A(_97_),
    .B(_136_),
    .C(_137_),
    .Y(_138_)
);

AOI21X1 _709_ (
    .A(_138_),
    .B(_135_),
    .C(_96_),
    .Y(_139_)
);

AOI21X1 _710_ (
    .A(_46_),
    .B(_85_),
    .C(_83_),
    .Y(_140_)
);

NAND3X1 _711_ (
    .A(_98_),
    .B(_136_),
    .C(_137_),
    .Y(_141_)
);

OAI21X1 _712_ (
    .A(_130_),
    .B(_134_),
    .C(_97_),
    .Y(_142_)
);

AOI21X1 _713_ (
    .A(_141_),
    .B(_142_),
    .C(_140_),
    .Y(_143_)
);

OAI21X1 _714_ (
    .A(_139_),
    .B(_143_),
    .C(_95_),
    .Y(_144_)
);

NAND3X1 _715_ (
    .A(_141_),
    .B(_142_),
    .C(_140_),
    .Y(_145_)
);

NAND3X1 _716_ (
    .A(_138_),
    .B(_135_),
    .C(_96_),
    .Y(_146_)
);

NAND3X1 _717_ (
    .A(_94_),
    .B(_145_),
    .C(_146_),
    .Y(_147_)
);

AOI21X1 _718_ (
    .A(_147_),
    .B(_144_),
    .C(_93_),
    .Y(_148_)
);

NAND3X1 _719_ (
    .A(_500_),
    .B(_515_),
    .C(_522_),
    .Y(_149_)
);

OAI21X1 _720_ (
    .A(_516_),
    .B(_511_),
    .C(_518_),
    .Y(_150_)
);

NAND2X1 _721_ (
    .A(_2_),
    .B(_529_),
    .Y(_151_)
);

AOI21X1 _722_ (
    .A(_150_),
    .B(_149_),
    .C(_151_),
    .Y(_152_)
);

NAND3X1 _723_ (
    .A(_150_),
    .B(_151_),
    .C(_149_),
    .Y(_153_)
);

AOI21X1 _724_ (
    .A(_7_),
    .B(_153_),
    .C(_152_),
    .Y(_154_)
);

NAND3X1 _725_ (
    .A(_12_),
    .B(_38_),
    .C(_37_),
    .Y(_155_)
);

OAI21X1 _726_ (
    .A(_35_),
    .B(_30_),
    .C(_11_),
    .Y(_156_)
);

AOI21X1 _727_ (
    .A(_155_),
    .B(_156_),
    .C(_154_),
    .Y(_157_)
);

NAND3X1 _728_ (
    .A(_155_),
    .B(_156_),
    .C(_154_),
    .Y(_158_)
);

AOI21X1 _729_ (
    .A(_43_),
    .B(_158_),
    .C(_157_),
    .Y(_159_)
);

NAND3X1 _730_ (
    .A(_47_),
    .B(_86_),
    .C(_85_),
    .Y(_160_)
);

OAI21X1 _731_ (
    .A(_79_),
    .B(_83_),
    .C(_46_),
    .Y(_161_)
);

AOI21X1 _732_ (
    .A(_160_),
    .B(_161_),
    .C(_159_),
    .Y(_162_)
);

NAND3X1 _733_ (
    .A(_160_),
    .B(_161_),
    .C(_159_),
    .Y(_163_)
);

AOI21X1 _734_ (
    .A(_91_),
    .B(_163_),
    .C(_162_),
    .Y(_164_)
);

NAND3X1 _735_ (
    .A(_95_),
    .B(_145_),
    .C(_146_),
    .Y(_165_)
);

OAI21X1 _736_ (
    .A(_139_),
    .B(_143_),
    .C(_94_),
    .Y(_166_)
);

AOI21X1 _737_ (
    .A(_165_),
    .B(_166_),
    .C(_164_),
    .Y(_167_)
);

OAI21X1 _738_ (
    .A(_148_),
    .B(_167_),
    .C(_499_),
    .Y(_168_)
);

NAND3X1 _739_ (
    .A(_165_),
    .B(_166_),
    .C(_164_),
    .Y(_169_)
);

NAND3X1 _740_ (
    .A(_147_),
    .B(_144_),
    .C(_93_),
    .Y(_170_)
);

NAND3X1 _741_ (
    .A(_498_),
    .B(_169_),
    .C(_170_),
    .Y(_171_)
);

AOI21X1 _742_ (
    .A(_171_),
    .B(_168_),
    .C(_495_),
    .Y(_172_)
);

NOR2X1 _743_ (
    .A(_496_),
    .B(_485_),
    .Y(_173_)
);

OAI21X1 _744_ (
    .A(_89_),
    .B(_162_),
    .C(_92_),
    .Y(_174_)
);

NAND3X1 _745_ (
    .A(_91_),
    .B(_163_),
    .C(_88_),
    .Y(_175_)
);

AOI21X1 _746_ (
    .A(_175_),
    .B(_174_),
    .C(_173_),
    .Y(_176_)
);

NOR2X1 _747_ (
    .A(_90_),
    .B(_485_),
    .Y(_177_)
);

OAI21X1 _748_ (
    .A(_41_),
    .B(_157_),
    .C(_43_),
    .Y(_178_)
);

NAND3X1 _749_ (
    .A(_44_),
    .B(_158_),
    .C(_40_),
    .Y(_179_)
);

NAND2X1 _750_ (
    .A(_179_),
    .B(_178_),
    .Y(_180_)
);

OR2X2 _751_ (
    .A(_180_),
    .B(_177_),
    .Y(_181_)
);

NOR2X1 _752_ (
    .A(_42_),
    .B(_485_),
    .Y(_182_)
);

INVX1 _753_ (
    .A(_182_),
    .Y(_183_)
);

OAI21X1 _754_ (
    .A(_5_),
    .B(_152_),
    .C(_8_),
    .Y(_184_)
);

NAND3X1 _755_ (
    .A(_153_),
    .B(_7_),
    .C(_4_),
    .Y(_185_)
);

NAND2X1 _756_ (
    .A(_185_),
    .B(_184_),
    .Y(_186_)
);

AOI21X1 _757_ (
    .A(_185_),
    .B(_184_),
    .C(_182_),
    .Y(_187_)
);

NOR2X1 _758_ (
    .A(_530_),
    .B(_497_),
    .Y(_188_)
);

NAND2X1 _759_ (
    .A(_531_),
    .B(_529_),
    .Y(_189_)
);

XOR2X1 _760_ (
    .A(_189_),
    .B(_188_),
    .Y(_190_)
);

OAI21X1 _761_ (
    .A(_6_),
    .B(_485_),
    .C(_190_),
    .Y(_191_)
);

NOR2X1 _762_ (
    .A(_508_),
    .B(_485_),
    .Y(_192_)
);

NAND2X1 _763_ (
    .A(_526_),
    .B(_192_),
    .Y(_193_)
);

INVX2 _764_ (
    .A(_193_),
    .Y(_194_)
);

OAI21X1 _765_ (
    .A(_508_),
    .B(_497_),
    .C(_513_),
    .Y(_195_)
);

NAND2X1 _766_ (
    .A(_195_),
    .B(_527_),
    .Y(_196_)
);

INVX1 _767_ (
    .A(_196_),
    .Y(_197_)
);

NAND2X1 _768_ (
    .A(_194_),
    .B(_197_),
    .Y(_198_)
);

NOR2X1 _769_ (
    .A(_194_),
    .B(_197_),
    .Y(_199_)
);

NOR2X1 _770_ (
    .A(_530_),
    .B(_485_),
    .Y(_200_)
);

INVX1 _771_ (
    .A(_200_),
    .Y(_201_)
);

OAI21X1 _772_ (
    .A(_199_),
    .B(_201_),
    .C(_198_),
    .Y(_202_)
);

NOR2X1 _773_ (
    .A(_6_),
    .B(_485_),
    .Y(_203_)
);

INVX1 _774_ (
    .A(_203_),
    .Y(_204_)
);

NOR2X1 _775_ (
    .A(_204_),
    .B(_190_),
    .Y(_205_)
);

OAI21X1 _776_ (
    .A(_205_),
    .B(_202_),
    .C(_191_),
    .Y(_206_)
);

OR2X2 _777_ (
    .A(_206_),
    .B(_187_),
    .Y(_207_)
);

OAI21X1 _778_ (
    .A(_183_),
    .B(_186_),
    .C(_207_),
    .Y(_208_)
);

INVX1 _779_ (
    .A(_177_),
    .Y(_209_)
);

AOI21X1 _780_ (
    .A(_179_),
    .B(_178_),
    .C(_209_),
    .Y(_210_)
);

OAI21X1 _781_ (
    .A(_208_),
    .B(_210_),
    .C(_181_),
    .Y(_211_)
);

NAND3X1 _782_ (
    .A(_173_),
    .B(_175_),
    .C(_174_),
    .Y(_212_)
);

AOI21X1 _783_ (
    .A(_211_),
    .B(_212_),
    .C(_176_),
    .Y(_213_)
);

INVX1 _784_ (
    .A(_213_),
    .Y(_214_)
);

NAND3X1 _785_ (
    .A(_495_),
    .B(_171_),
    .C(_168_),
    .Y(_215_)
);

AOI21X1 _786_ (
    .A(_214_),
    .B(_215_),
    .C(_172_),
    .Y(\partialsco[7] [0])
);

OAI21X1 _787_ (
    .A(_139_),
    .B(_95_),
    .C(_146_),
    .Y(_216_)
);

AOI21X1 _788_ (
    .A(_97_),
    .B(_136_),
    .C(_134_),
    .Y(_217_)
);

AOI21X1 _789_ (
    .A(_100_),
    .B(_127_),
    .C(_125_),
    .Y(_218_)
);

AOI21X1 _790_ (
    .A(_103_),
    .B(_118_),
    .C(_113_),
    .Y(_219_)
);

NAND2X1 _791_ (
    .A(areg[2]),
    .B(breg[6]),
    .Y(_220_)
);

AOI21X1 _792_ (
    .A(_58_),
    .B(_105_),
    .C(_220_),
    .Y(_221_)
);

INVX1 _793_ (
    .A(_221_),
    .Y(_222_)
);

NAND3X1 _794_ (
    .A(_58_),
    .B(_220_),
    .C(_105_),
    .Y(_223_)
);

NOR2X1 _795_ (
    .A(_6_),
    .B(_57_),
    .Y(_224_)
);

AOI21X1 _796_ (
    .A(_223_),
    .B(_222_),
    .C(_224_),
    .Y(_225_)
);

INVX2 _797_ (
    .A(_223_),
    .Y(_226_)
);

INVX2 _798_ (
    .A(_224_),
    .Y(_227_)
);

NOR3X1 _799_ (
    .A(_221_),
    .B(_227_),
    .C(_226_),
    .Y(_228_)
);

OAI21X1 _800_ (
    .A(_228_),
    .B(_225_),
    .C(_219_),
    .Y(_229_)
);

OAI21X1 _801_ (
    .A(_110_),
    .B(_104_),
    .C(_119_),
    .Y(_230_)
);

OAI21X1 _802_ (
    .A(_226_),
    .B(_221_),
    .C(_227_),
    .Y(_231_)
);

NAND3X1 _803_ (
    .A(_223_),
    .B(_224_),
    .C(_222_),
    .Y(_232_)
);

NAND3X1 _804_ (
    .A(_231_),
    .B(_232_),
    .C(_230_),
    .Y(_233_)
);

NOR2X1 _805_ (
    .A(_42_),
    .B(_19_),
    .Y(_234_)
);

AOI21X1 _806_ (
    .A(_229_),
    .B(_233_),
    .C(_234_),
    .Y(_235_)
);

AOI21X1 _807_ (
    .A(_232_),
    .B(_231_),
    .C(_230_),
    .Y(_236_)
);

NOR3X1 _808_ (
    .A(_228_),
    .B(_225_),
    .C(_219_),
    .Y(_237_)
);

INVX2 _809_ (
    .A(_234_),
    .Y(_238_)
);

NOR3X1 _810_ (
    .A(_236_),
    .B(_238_),
    .C(_237_),
    .Y(_239_)
);

OAI21X1 _811_ (
    .A(_239_),
    .B(_235_),
    .C(_218_),
    .Y(_240_)
);

OAI21X1 _812_ (
    .A(_121_),
    .B(_101_),
    .C(_128_),
    .Y(_241_)
);

OAI21X1 _813_ (
    .A(_237_),
    .B(_236_),
    .C(_238_),
    .Y(_242_)
);

NAND3X1 _814_ (
    .A(_234_),
    .B(_229_),
    .C(_233_),
    .Y(_243_)
);

NAND3X1 _815_ (
    .A(_241_),
    .B(_243_),
    .C(_242_),
    .Y(_244_)
);

NOR2X1 _816_ (
    .A(_507_),
    .B(_90_),
    .Y(_245_)
);

AOI21X1 _817_ (
    .A(_244_),
    .B(_240_),
    .C(_245_),
    .Y(_246_)
);

AOI21X1 _818_ (
    .A(_243_),
    .B(_242_),
    .C(_241_),
    .Y(_247_)
);

NOR3X1 _819_ (
    .A(_218_),
    .B(_235_),
    .C(_239_),
    .Y(_248_)
);

INVX2 _820_ (
    .A(_245_),
    .Y(_249_)
);

NOR3X1 _821_ (
    .A(_247_),
    .B(_249_),
    .C(_248_),
    .Y(_250_)
);

OAI21X1 _822_ (
    .A(_250_),
    .B(_246_),
    .C(_217_),
    .Y(_251_)
);

INVX2 _823_ (
    .A(_217_),
    .Y(_252_)
);

OAI21X1 _824_ (
    .A(_248_),
    .B(_247_),
    .C(_249_),
    .Y(_253_)
);

NAND3X1 _825_ (
    .A(_244_),
    .B(_245_),
    .C(_240_),
    .Y(_254_)
);

NAND3X1 _826_ (
    .A(_253_),
    .B(_254_),
    .C(_252_),
    .Y(_255_)
);

NOR2X1 _827_ (
    .A(_10_),
    .B(_496_),
    .Y(_256_)
);

AOI21X1 _828_ (
    .A(_251_),
    .B(_255_),
    .C(_256_),
    .Y(_257_)
);

AOI21X1 _829_ (
    .A(_254_),
    .B(_253_),
    .C(_252_),
    .Y(_258_)
);

NOR3X1 _830_ (
    .A(_217_),
    .B(_246_),
    .C(_250_),
    .Y(_259_)
);

INVX2 _831_ (
    .A(_256_),
    .Y(_260_)
);

NOR3X1 _832_ (
    .A(_258_),
    .B(_260_),
    .C(_259_),
    .Y(_261_)
);

OAI21X1 _833_ (
    .A(_261_),
    .B(_257_),
    .C(_216_),
    .Y(_262_)
);

INVX2 _834_ (
    .A(_216_),
    .Y(_263_)
);

OAI21X1 _835_ (
    .A(_259_),
    .B(_258_),
    .C(_260_),
    .Y(_264_)
);

NAND3X1 _836_ (
    .A(_256_),
    .B(_251_),
    .C(_255_),
    .Y(_265_)
);

NAND3X1 _837_ (
    .A(_265_),
    .B(_264_),
    .C(_263_),
    .Y(_266_)
);

NOR2X1 _838_ (
    .A(_497_),
    .B(_494_),
    .Y(_267_)
);

AOI21X1 _839_ (
    .A(_266_),
    .B(_262_),
    .C(_267_),
    .Y(_268_)
);

OAI21X1 _840_ (
    .A(_148_),
    .B(_499_),
    .C(_170_),
    .Y(_269_)
);

INVX1 _841_ (
    .A(_269_),
    .Y(_270_)
);

AOI21X1 _842_ (
    .A(_265_),
    .B(_264_),
    .C(_263_),
    .Y(_271_)
);

NOR3X1 _843_ (
    .A(_216_),
    .B(_257_),
    .C(_261_),
    .Y(_272_)
);

INVX1 _844_ (
    .A(_267_),
    .Y(_273_)
);

NOR3X1 _845_ (
    .A(_271_),
    .B(_273_),
    .C(_272_),
    .Y(_274_)
);

INVX1 _846_ (
    .A(_274_),
    .Y(_275_)
);

AOI21X1 _847_ (
    .A(_270_),
    .B(_275_),
    .C(_268_),
    .Y(\partialsco[7] [1])
);

OAI21X1 _848_ (
    .A(_507_),
    .B(_90_),
    .C(_217_),
    .Y(_276_)
);

NOR2X1 _849_ (
    .A(_247_),
    .B(_248_),
    .Y(_277_)
);

OAI21X1 _850_ (
    .A(_217_),
    .B(_249_),
    .C(_277_),
    .Y(_278_)
);

AND2X2 _851_ (
    .A(_278_),
    .B(_276_),
    .Y(_279_)
);

NOR2X1 _852_ (
    .A(_236_),
    .B(_237_),
    .Y(_280_)
);

OAI21X1 _853_ (
    .A(_218_),
    .B(_238_),
    .C(_280_),
    .Y(_281_)
);

OAI21X1 _854_ (
    .A(_241_),
    .B(_234_),
    .C(_281_),
    .Y(_282_)
);

INVX1 _855_ (
    .A(_282_),
    .Y(_283_)
);

NOR2X1 _856_ (
    .A(_221_),
    .B(_226_),
    .Y(_284_)
);

OAI21X1 _857_ (
    .A(_219_),
    .B(_227_),
    .C(_284_),
    .Y(_285_)
);

OAI21X1 _858_ (
    .A(_230_),
    .B(_224_),
    .C(_285_),
    .Y(_286_)
);

AOI21X1 _859_ (
    .A(_58_),
    .B(_220_),
    .C(_115_),
    .Y(_287_)
);

NAND2X1 _860_ (
    .A(areg[2]),
    .B(breg[7]),
    .Y(_288_)
);

NAND2X1 _861_ (
    .A(areg[3]),
    .B(breg[6]),
    .Y(_289_)
);

XNOR2X1 _862_ (
    .A(_288_),
    .B(_289_),
    .Y(_290_)
);

NOR2X1 _863_ (
    .A(_287_),
    .B(_290_),
    .Y(_291_)
);

AND2X2 _864_ (
    .A(_290_),
    .B(_287_),
    .Y(_292_)
);

NOR2X1 _865_ (
    .A(_291_),
    .B(_292_),
    .Y(_293_)
);

NOR2X1 _866_ (
    .A(_42_),
    .B(_57_),
    .Y(_294_)
);

XNOR2X1 _867_ (
    .A(_293_),
    .B(_294_),
    .Y(_295_)
);

AND2X2 _868_ (
    .A(_295_),
    .B(_286_),
    .Y(_296_)
);

NOR2X1 _869_ (
    .A(_286_),
    .B(_295_),
    .Y(_297_)
);

NOR2X1 _870_ (
    .A(_90_),
    .B(_19_),
    .Y(_298_)
);

INVX1 _871_ (
    .A(_298_),
    .Y(_299_)
);

OAI21X1 _872_ (
    .A(_296_),
    .B(_297_),
    .C(_299_),
    .Y(_300_)
);

NAND2X1 _873_ (
    .A(_286_),
    .B(_295_),
    .Y(_301_)
);

OR2X2 _874_ (
    .A(_295_),
    .B(_286_),
    .Y(_302_)
);

NAND3X1 _875_ (
    .A(_301_),
    .B(_298_),
    .C(_302_),
    .Y(_303_)
);

AOI21X1 _876_ (
    .A(_300_),
    .B(_303_),
    .C(_283_),
    .Y(_304_)
);

INVX1 _877_ (
    .A(_304_),
    .Y(_305_)
);

NAND2X1 _878_ (
    .A(_300_),
    .B(_303_),
    .Y(_306_)
);

OR2X2 _879_ (
    .A(_306_),
    .B(_282_),
    .Y(_307_)
);

NOR2X1 _880_ (
    .A(_507_),
    .B(_496_),
    .Y(_308_)
);

AOI21X1 _881_ (
    .A(_305_),
    .B(_307_),
    .C(_308_),
    .Y(_309_)
);

NOR2X1 _882_ (
    .A(_282_),
    .B(_306_),
    .Y(_310_)
);

INVX2 _883_ (
    .A(_308_),
    .Y(_311_)
);

NOR3X1 _884_ (
    .A(_304_),
    .B(_311_),
    .C(_310_),
    .Y(_312_)
);

OAI21X1 _885_ (
    .A(_309_),
    .B(_312_),
    .C(_279_),
    .Y(_313_)
);

OAI21X1 _886_ (
    .A(_252_),
    .B(_245_),
    .C(_278_),
    .Y(_314_)
);

OAI21X1 _887_ (
    .A(_310_),
    .B(_304_),
    .C(_311_),
    .Y(_315_)
);

NAND3X1 _888_ (
    .A(_305_),
    .B(_308_),
    .C(_307_),
    .Y(_316_)
);

NAND3X1 _889_ (
    .A(_314_),
    .B(_315_),
    .C(_316_),
    .Y(_317_)
);

NOR2X1 _890_ (
    .A(_10_),
    .B(_494_),
    .Y(_318_)
);

AOI21X1 _891_ (
    .A(_317_),
    .B(_313_),
    .C(_318_),
    .Y(_319_)
);

OAI22X1 _892_ (
    .A(_258_),
    .B(_259_),
    .C(_216_),
    .D(_256_),
    .Y(_320_)
);

OAI21X1 _893_ (
    .A(_263_),
    .B(_260_),
    .C(_320_),
    .Y(_321_)
);

INVX1 _894_ (
    .A(_321_),
    .Y(_322_)
);

NAND3X1 _895_ (
    .A(_317_),
    .B(_318_),
    .C(_313_),
    .Y(_323_)
);

AOI21X1 _896_ (
    .A(_322_),
    .B(_323_),
    .C(_319_),
    .Y(\partialsco[7] [2])
);

OAI22X1 _897_ (
    .A(_296_),
    .B(_297_),
    .C(_283_),
    .D(_298_),
    .Y(_324_)
);

OAI21X1 _898_ (
    .A(_282_),
    .B(_299_),
    .C(_324_),
    .Y(_325_)
);

OAI21X1 _899_ (
    .A(_6_),
    .B(_57_),
    .C(_219_),
    .Y(_326_)
);

AND2X2 _900_ (
    .A(_285_),
    .B(_326_),
    .Y(_327_)
);

NAND2X1 _901_ (
    .A(_294_),
    .B(_327_),
    .Y(_328_)
);

INVX1 _902_ (
    .A(_293_),
    .Y(_329_)
);

OAI21X1 _903_ (
    .A(_327_),
    .B(_294_),
    .C(_329_),
    .Y(_330_)
);

NAND2X1 _904_ (
    .A(_328_),
    .B(_330_),
    .Y(_331_)
);

INVX1 _905_ (
    .A(_289_),
    .Y(_332_)
);

INVX1 _906_ (
    .A(_287_),
    .Y(_333_)
);

OAI21X1 _907_ (
    .A(_333_),
    .B(_289_),
    .C(_288_),
    .Y(_334_)
);

OAI21X1 _908_ (
    .A(_287_),
    .B(_332_),
    .C(_334_),
    .Y(_335_)
);

NAND2X1 _909_ (
    .A(areg[3]),
    .B(breg[7]),
    .Y(_336_)
);

NAND2X1 _910_ (
    .A(areg[4]),
    .B(breg[6]),
    .Y(_337_)
);

XOR2X1 _911_ (
    .A(_336_),
    .B(_337_),
    .Y(_338_)
);

NOR2X1 _912_ (
    .A(_338_),
    .B(_335_),
    .Y(_339_)
);

AND2X2 _913_ (
    .A(_335_),
    .B(_338_),
    .Y(_340_)
);

NOR2X1 _914_ (
    .A(_90_),
    .B(_57_),
    .Y(_341_)
);

INVX1 _915_ (
    .A(_341_),
    .Y(_342_)
);

OAI21X1 _916_ (
    .A(_340_),
    .B(_339_),
    .C(_342_),
    .Y(_343_)
);

NOR2X1 _917_ (
    .A(_339_),
    .B(_340_),
    .Y(_344_)
);

NAND2X1 _918_ (
    .A(_341_),
    .B(_344_),
    .Y(_345_)
);

NAND2X1 _919_ (
    .A(_343_),
    .B(_345_),
    .Y(_346_)
);

INVX1 _920_ (
    .A(_346_),
    .Y(_347_)
);

NOR2X1 _921_ (
    .A(_331_),
    .B(_347_),
    .Y(_348_)
);

AND2X2 _922_ (
    .A(_330_),
    .B(_328_),
    .Y(_349_)
);

NOR2X1 _923_ (
    .A(_346_),
    .B(_349_),
    .Y(_350_)
);

NOR2X1 _924_ (
    .A(_496_),
    .B(_19_),
    .Y(_351_)
);

INVX1 _925_ (
    .A(_351_),
    .Y(_352_)
);

OAI21X1 _926_ (
    .A(_348_),
    .B(_350_),
    .C(_352_),
    .Y(_353_)
);

NAND2X1 _927_ (
    .A(_346_),
    .B(_349_),
    .Y(_354_)
);

NAND2X1 _928_ (
    .A(_331_),
    .B(_347_),
    .Y(_355_)
);

NAND3X1 _929_ (
    .A(_354_),
    .B(_351_),
    .C(_355_),
    .Y(_356_)
);

NAND2X1 _930_ (
    .A(_356_),
    .B(_353_),
    .Y(_357_)
);

NAND2X1 _931_ (
    .A(_325_),
    .B(_357_),
    .Y(_358_)
);

OR2X2 _932_ (
    .A(_357_),
    .B(_325_),
    .Y(_359_)
);

NOR2X1 _933_ (
    .A(_507_),
    .B(_494_),
    .Y(_360_)
);

AOI21X1 _934_ (
    .A(_358_),
    .B(_359_),
    .C(_360_),
    .Y(_361_)
);

NOR2X1 _935_ (
    .A(_304_),
    .B(_310_),
    .Y(_362_)
);

INVX1 _936_ (
    .A(_362_),
    .Y(_363_)
);

OAI21X1 _937_ (
    .A(_507_),
    .B(_496_),
    .C(_314_),
    .Y(_364_)
);

NOR2X1 _938_ (
    .A(_311_),
    .B(_314_),
    .Y(_365_)
);

OAI21X1 _939_ (
    .A(_363_),
    .B(_365_),
    .C(_364_),
    .Y(_366_)
);

NAND3X1 _940_ (
    .A(_358_),
    .B(_360_),
    .C(_359_),
    .Y(_367_)
);

AOI21X1 _941_ (
    .A(_366_),
    .B(_367_),
    .C(_361_),
    .Y(\partialsco[7] [3])
);

OAI21X1 _942_ (
    .A(_90_),
    .B(_57_),
    .C(_349_),
    .Y(_368_)
);

OAI21X1 _943_ (
    .A(_349_),
    .B(_342_),
    .C(_344_),
    .Y(_369_)
);

INVX2 _944_ (
    .A(breg[6]),
    .Y(_370_)
);

OAI21X1 _945_ (
    .A(_42_),
    .B(_370_),
    .C(_335_),
    .Y(_371_)
);

OAI21X1 _946_ (
    .A(_335_),
    .B(_337_),
    .C(_336_),
    .Y(_372_)
);

NAND2X1 _947_ (
    .A(_371_),
    .B(_372_),
    .Y(_373_)
);

NAND2X1 _948_ (
    .A(areg[4]),
    .B(breg[7]),
    .Y(_374_)
);

NOR2X1 _949_ (
    .A(_90_),
    .B(_370_),
    .Y(_375_)
);

XNOR2X1 _950_ (
    .A(_375_),
    .B(_374_),
    .Y(_376_)
);

XNOR2X1 _951_ (
    .A(_373_),
    .B(_376_),
    .Y(_377_)
);

OAI21X1 _952_ (
    .A(_496_),
    .B(_57_),
    .C(_377_),
    .Y(_378_)
);

NOR2X1 _953_ (
    .A(_496_),
    .B(_57_),
    .Y(_379_)
);

INVX1 _954_ (
    .A(_379_),
    .Y(_380_)
);

OR2X2 _955_ (
    .A(_377_),
    .B(_380_),
    .Y(_381_)
);

NAND2X1 _956_ (
    .A(_378_),
    .B(_381_),
    .Y(_382_)
);

NAND3X1 _957_ (
    .A(_368_),
    .B(_369_),
    .C(_382_),
    .Y(_383_)
);

OAI21X1 _958_ (
    .A(_331_),
    .B(_341_),
    .C(_369_),
    .Y(_384_)
);

NAND3X1 _959_ (
    .A(_378_),
    .B(_381_),
    .C(_384_),
    .Y(_385_)
);

NAND2X1 _960_ (
    .A(_383_),
    .B(_385_),
    .Y(_386_)
);

OAI21X1 _961_ (
    .A(_494_),
    .B(_19_),
    .C(_386_),
    .Y(_387_)
);

NAND2X1 _962_ (
    .A(_351_),
    .B(_325_),
    .Y(_388_)
);

NAND3X1 _963_ (
    .A(_354_),
    .B(_355_),
    .C(_388_),
    .Y(_389_)
);

OAI21X1 _964_ (
    .A(_325_),
    .B(_351_),
    .C(_389_),
    .Y(_390_)
);

NOR2X1 _965_ (
    .A(_494_),
    .B(_19_),
    .Y(_391_)
);

NAND3X1 _966_ (
    .A(_391_),
    .B(_383_),
    .C(_385_),
    .Y(_392_)
);

NAND2X1 _967_ (
    .A(_392_),
    .B(_390_),
    .Y(_393_)
);

AND2X2 _968_ (
    .A(_393_),
    .B(_387_),
    .Y(\partialsco[7] [4])
);

NOR2X1 _969_ (
    .A(_90_),
    .B(_107_),
    .Y(_394_)
);

INVX1 _970_ (
    .A(_373_),
    .Y(_395_)
);

NOR2X1 _971_ (
    .A(_375_),
    .B(_395_),
    .Y(_396_)
);

NAND2X1 _972_ (
    .A(_375_),
    .B(_395_),
    .Y(_397_)
);

OAI21X1 _973_ (
    .A(_396_),
    .B(_374_),
    .C(_397_),
    .Y(_398_)
);

NOR2X1 _974_ (
    .A(_496_),
    .B(_370_),
    .Y(_399_)
);

XNOR2X1 _975_ (
    .A(_398_),
    .B(_399_),
    .Y(_400_)
);

XNOR2X1 _976_ (
    .A(_400_),
    .B(_394_),
    .Y(_401_)
);

NOR2X1 _977_ (
    .A(_494_),
    .B(_57_),
    .Y(_402_)
);

NOR2X1 _978_ (
    .A(_402_),
    .B(_401_),
    .Y(_403_)
);

OAI21X1 _979_ (
    .A(_496_),
    .B(_57_),
    .C(_384_),
    .Y(_404_)
);

NOR2X1 _980_ (
    .A(_380_),
    .B(_384_),
    .Y(_405_)
);

AOI21X1 _981_ (
    .A(_377_),
    .B(_404_),
    .C(_405_),
    .Y(_406_)
);

NAND2X1 _982_ (
    .A(_402_),
    .B(_401_),
    .Y(_407_)
);

AOI21X1 _983_ (
    .A(_406_),
    .B(_407_),
    .C(_403_),
    .Y(\partialsco[7] [5])
);

NOR2X1 _984_ (
    .A(_494_),
    .B(_107_),
    .Y(\partialsb[7] [7])
);

NAND2X1 _985_ (
    .A(_399_),
    .B(\partialsb[7] [7]),
    .Y(_408_)
);

NAND2X1 _986_ (
    .A(_399_),
    .B(_398_),
    .Y(_409_)
);

OAI21X1 _987_ (
    .A(_398_),
    .B(_399_),
    .C(_394_),
    .Y(_410_)
);

NAND2X1 _988_ (
    .A(_409_),
    .B(_410_),
    .Y(_411_)
);

INVX1 _989_ (
    .A(_411_),
    .Y(_412_)
);

AOI22X1 _990_ (
    .A(areg[6]),
    .B(breg[7]),
    .C(areg[7]),
    .D(breg[6]),
    .Y(_413_)
);

OAI21X1 _991_ (
    .A(_412_),
    .B(_413_),
    .C(_408_),
    .Y(\partialsco[7] [6])
);

NOR2X1 _992_ (
    .A(_526_),
    .B(_192_),
    .Y(_414_)
);

NOR2X1 _993_ (
    .A(_414_),
    .B(_194_),
    .Y(\partialss[1] [0])
);

INVX1 _994_ (
    .A(_205_),
    .Y(_415_)
);

NAND2X1 _995_ (
    .A(_191_),
    .B(_415_),
    .Y(_416_)
);

XNOR2X1 _996_ (
    .A(_416_),
    .B(_202_),
    .Y(\partialss[3] [0])
);

NOR2X1 _997_ (
    .A(_183_),
    .B(_186_),
    .Y(_417_)
);

NOR2X1 _998_ (
    .A(_187_),
    .B(_417_),
    .Y(_418_)
);

XNOR2X1 _999_ (
    .A(_418_),
    .B(_206_),
    .Y(\partialss[4] [0])
);

endmodule
