/* Verilog module written by vlog2Verilog (qflow) */
/* With explicit power connections */

module multiplier(
    inout vdd,
    inout gnd,
    input [15:0] a,
    input [15:0] b,
    input clk,
    output [31:0] y
);

wire [15:0] a ;
wire [15:0] b ;
wire _1677_ ;
wire _1257_ ;
wire [31:0] y ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _2712_ ;
wire _2521_ ;
wire _2101_ ;
wire _703_ ;
wire _1389_ ;
wire _2330_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1830_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _2615_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _2424_ ;
wire _2004_ ;
wire _606_ ;
wire _2653_ ;
wire _2233_ ;
wire _1924_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _2709_ ;
wire _95_ ;
wire _2462_ ;
wire _2042_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _2518_ ;
wire _2691_ ;
wire _2271_ ;
wire _1962_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _2327_ ;
wire _2080_ ;
wire _929_ ;
wire _509_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _2556_ ;
wire _2136_ ;
wire _1827_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _2365_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _2594_ ;
wire _2174_ ;
wire _1865_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _2459_ ;
wire _2039_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _2688_ ;
wire _2268_ ;
wire _1959_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _2497_ ;
wire _2077_ ;
wire _1768_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1997_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire areg_7_bF$buf0 ;
wire areg_7_bF$buf1 ;
wire areg_7_bF$buf2 ;
wire areg_7_bF$buf3 ;
wire _16_ ;
wire _1195_ ;
wire _2612_ ;
wire _54_ ;
wire _2421_ ;
wire _2001_ ;
wire _603_ ;
wire _1289_ ;
wire _2650_ ;
wire _2230_ ;
wire _1921_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _2706_ ;
wire _92_ ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _2515_ ;
wire _870_ ;
wire _450_ ;
wire [31:0] _2744_ ;
wire _2324_ ;
wire _926_ ;
wire _506_ ;
wire _2553_ ;
wire _2133_ ;
wire _1824_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _2609_ ;
wire _2362_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _2418_ ;
wire _2591_ ;
wire _2171_ ;
wire _1862_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _2647_ ;
wire _2227_ ;
wire _1918_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _2456_ ;
wire _2036_ ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _2685_ ;
wire _2265_ ;
wire _1956_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _2494_ ;
wire _2074_ ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1994_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _2359_ ;
wire _1383_ ;
wire _294_ ;
wire _2588_ ;
wire _2168_ ;
wire _13_ ;
wire _1859_ ;
wire _1439_ ;
wire _1019_ ;
wire _1192_ ;
wire _2397_ ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1897_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _2703_ ;
wire _1095_ ;
wire _2512_ ;
wire _2741_ ;
wire _2321_ ;
wire _7_ ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _2550_ ;
wire _2130_ ;
wire _1821_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire _2606_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _2415_ ;
wire _770_ ;
wire _350_ ;
wire _2644_ ;
wire _2224_ ;
wire _1915_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _2453_ ;
wire _2033_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _2509_ ;
wire _2682_ ;
wire _2262_ ;
wire _1953_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _2738_ ;
wire _2318_ ;
wire _2491_ ;
wire _2071_ ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _2547_ ;
wire _2127_ ;
wire _1818_ ;
wire _729_ ;
wire _309_ ;
wire _1991_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _2356_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _2585_ ;
wire _2165_ ;
wire _10_ ;
wire _1856_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _2394_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1894_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _2679_ ;
wire _2259_ ;
wire _1283_ ;
wire _194_ ;
wire _2488_ ;
wire _2068_ ;
wire _1759_ ;
wire _1339_ ;
wire _2700_ ;
wire _1092_ ;
wire _2297_ ;
wire _1988_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _1797_ ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _2603_ ;
wire _45_ ;
wire _2412_ ;
wire _2641_ ;
wire _2221_ ;
wire _1912_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _2450_ ;
wire _2030_ ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _2506_ ;
wire _1950_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _2735_ ;
wire _2315_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _2544_ ;
wire _2124_ ;
wire _1815_ ;
wire _726_ ;
wire _306_ ;
wire _2353_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _2409_ ;
wire _2582_ ;
wire _2162_ ;
wire _1853_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _2638_ ;
wire _2218_ ;
wire _2391_ ;
wire _1909_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _2447_ ;
wire _2027_ ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1891_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _2676_ ;
wire _2256_ ;
wire _1947_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _2485_ ;
wire _2065_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _2294_ ;
wire _1985_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1794_ ;
wire _1374_ ;
wire _285_ ;
wire _2579_ ;
wire _2159_ ;
wire _1_ ;
wire _1183_ ;
wire _2388_ ;
wire _1659_ ;
wire _1239_ ;
wire _2600_ ;
wire _2197_ ;
wire _42_ ;
wire _1888_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _2503_ ;
wire _2732_ ;
wire _2312_ ;
wire _914_ ;
wire _2541_ ;
wire _2121_ ;
wire _1812_ ;
wire _723_ ;
wire _303_ ;
wire _2350_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _2406_ ;
wire _1850_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _2635_ ;
wire _2215_ ;
wire clk ;
wire _1906_ ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _2444_ ;
wire _2024_ ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire _2673_ ;
wire _2253_ ;
wire _1944_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _2729_ ;
wire _2309_ ;
wire _2482_ ;
wire _2062_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _2538_ ;
wire _2118_ ;
wire _2291_ ;
wire _1809_ ;
wire _1982_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _2347_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1791_ ;
wire _1371_ ;
wire _282_ ;
wire _2576_ ;
wire _2156_ ;
wire _1847_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _2385_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _2194_ ;
wire _1885_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _2479_ ;
wire _2059_ ;
wire _1083_ ;
wire _2288_ ;
wire _1979_ ;
wire _1559_ ;
wire _1139_ ;
wire _2500_ ;
wire _2097_ ;
wire _1788_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _2403_ ;
wire _2632_ ;
wire _2212_ ;
wire _1903_ ;
wire _814_ ;
wire _74_ ;
wire _2441_ ;
wire _2021_ ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _2670_ ;
wire _2250_ ;
wire _1941_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _2726_ ;
wire _2306_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _2535_ ;
wire _2115_ ;
wire _1806_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _2344_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _2573_ ;
wire _2153_ ;
wire _1844_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _2629_ ;
wire _2209_ ;
wire _2382_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _2438_ ;
wire _2018_ ;
wire _2191_ ;
wire _1709_ ;
wire _1882_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _2667_ ;
wire _2247_ ;
wire _1938_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _2476_ ;
wire _2056_ ;
wire _1747_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _2285_ ;
wire _1976_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _2094_ ;
wire _1785_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire _2379_ ;
wire _2188_ ;
wire _33_ ;
wire _1879_ ;
wire _1459_ ;
wire _1039_ ;
wire _2400_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _1900_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _2723_ ;
wire _2303_ ;
wire _905_ ;
wire _2532_ ;
wire _2112_ ;
wire _1803_ ;
wire _714_ ;
wire _2341_ ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _2570_ ;
wire _2150_ ;
wire _1841_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _2626_ ;
wire _2206_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _2435_ ;
wire _2015_ ;
wire _1706_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _2664_ ;
wire _2244_ ;
wire _1935_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _2473_ ;
wire _2053_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _2529_ ;
wire _2109_ ;
wire _2282_ ;
wire _1973_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _2338_ ;
wire _2091_ ;
wire _1609_ ;
wire _1782_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _2567_ ;
wire _2147_ ;
wire _1838_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _2376_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _2185_ ;
wire _30_ ;
wire _1876_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire _2699_ ;
wire _2279_ ;
wire _2088_ ;
wire _1779_ ;
wire _1359_ ;
wire _2720_ ;
wire _2300_ ;
wire areg_4_bF$buf0 ;
wire areg_4_bF$buf1 ;
wire areg_4_bF$buf2 ;
wire areg_4_bF$buf3 ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _1800_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire _2623_ ;
wire _2203_ ;
wire _805_ ;
wire _65_ ;
wire _2432_ ;
wire _2012_ ;
wire _1703_ ;
wire _614_ ;
wire _2661_ ;
wire _2241_ ;
wire _1932_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _2717_ ;
wire _2470_ ;
wire _2050_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _2526_ ;
wire _2106_ ;
wire _708_ ;
wire _1970_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _2335_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _2564_ ;
wire _2144_ ;
wire _1835_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _2373_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _2429_ ;
wire _2009_ ;
wire _2182_ ;
wire _1873_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _2658_ ;
wire _2238_ ;
wire _1929_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _2467_ ;
wire _2047_ ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _2696_ ;
wire _2276_ ;
wire _1967_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _2085_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _2599_ ;
wire _2179_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _2620_ ;
wire _2200_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire _2714_ ;
wire _2523_ ;
wire _2103_ ;
wire _705_ ;
wire _2332_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _2561_ ;
wire _2141_ ;
wire _1832_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _2617_ ;
wire _2370_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _2426_ ;
wire _2006_ ;
wire _608_ ;
wire _1870_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _2655_ ;
wire _2235_ ;
wire _1926_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _2464_ ;
wire _2044_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _2693_ ;
wire _2273_ ;
wire _1964_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _2329_ ;
wire _2082_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _2558_ ;
wire _2138_ ;
wire _1829_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _2367_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _2596_ ;
wire _2176_ ;
wire _21_ ;
wire _1867_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire _2499_ ;
wire _2079_ ;
wire _2711_ ;
wire _1999_ ;
wire _1579_ ;
wire _1159_ ;
wire _2520_ ;
wire _2100_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _2614_ ;
wire _56_ ;
wire _2423_ ;
wire _2003_ ;
wire _605_ ;
wire _2652_ ;
wire _2232_ ;
wire _1923_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _2708_ ;
wire _94_ ;
wire _2461_ ;
wire _2041_ ;
wire aregp1_11_bF$buf0 ;
wire aregp1_11_bF$buf1 ;
wire aregp1_11_bF$buf2 ;
wire aregp1_11_bF$buf3 ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _2517_ ;
wire _2690_ ;
wire _2270_ ;
wire _1961_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _2326_ ;
wire _928_ ;
wire _508_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _2555_ ;
wire _2135_ ;
wire _1826_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _2364_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _2593_ ;
wire _2173_ ;
wire _1864_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _2649_ ;
wire _2229_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _2458_ ;
wire _2038_ ;
wire _1729_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _2687_ ;
wire _2267_ ;
wire _1958_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _2496_ ;
wire _2076_ ;
wire _1767_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1996_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _2399_ ;
wire _2611_ ;
wire _53_ ;
wire _1899_ ;
wire _1479_ ;
wire _1059_ ;
wire _2420_ ;
wire _2000_ ;
wire _602_ ;
wire [15:0] breg ;
wire _1288_ ;
wire _199_ ;
wire _1920_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _2705_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _2514_ ;
wire _2743_ ;
wire _2323_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire _2552_ ;
wire _2132_ ;
wire _1823_ ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _2608_ ;
wire _2361_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _2417_ ;
wire _2590_ ;
wire _2170_ ;
wire _1861_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _2646_ ;
wire _2226_ ;
wire _1917_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _2455_ ;
wire _2035_ ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _2684_ ;
wire _2264_ ;
wire _1955_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _2493_ ;
wire _2073_ ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _2549_ ;
wire _2129_ ;
wire _1993_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _2358_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _2587_ ;
wire _2167_ ;
wire _12_ ;
wire _1858_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _2396_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1896_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _2702_ ;
wire _1094_ ;
wire _2299_ ;
wire _2511_ ;
wire _1799_ ;
wire _1379_ ;
wire _2740_ ;
wire _2320_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire [15:0] areg ;
wire _1188_ ;
wire _1820_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _2605_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _2414_ ;
wire _2643_ ;
wire _2223_ ;
wire _1914_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _2452_ ;
wire _2032_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _2508_ ;
wire _2681_ ;
wire _2261_ ;
wire _1952_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _2737_ ;
wire _2317_ ;
wire _2490_ ;
wire _2070_ ;
wire _919_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _2546_ ;
wire _2126_ ;
wire _1817_ ;
wire _728_ ;
wire _308_ ;
wire _1990_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _2355_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _2584_ ;
wire _2164_ ;
wire _1855_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _2393_ ;
wire areg_6_bF$buf0 ;
wire areg_6_bF$buf1 ;
wire areg_6_bF$buf2 ;
wire areg_6_bF$buf3 ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _2449_ ;
wire _2029_ ;
wire _1893_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _2678_ ;
wire _2258_ ;
wire _1949_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _2487_ ;
wire _2067_ ;
wire _1758_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _2296_ ;
wire _1987_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1796_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _2602_ ;
wire _2199_ ;
wire _44_ ;
wire _2411_ ;
wire _1699_ ;
wire _1279_ ;
wire _2640_ ;
wire _2220_ ;
wire _1911_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _2505_ ;
wire _860_ ;
wire _440_ ;
wire _2734_ ;
wire _2314_ ;
wire _916_ ;
wire _2543_ ;
wire _2123_ ;
wire _1814_ ;
wire _725_ ;
wire _305_ ;
wire _2352_ ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _2408_ ;
wire _2581_ ;
wire _2161_ ;
wire _1852_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _2637_ ;
wire _2217_ ;
wire _2390_ ;
wire _1908_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _2446_ ;
wire _2026_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1890_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _2675_ ;
wire _2255_ ;
wire _1946_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _2484_ ;
wire _2064_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _2293_ ;
wire _1984_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _2349_ ;
wire _1793_ ;
wire _1373_ ;
wire _284_ ;
wire _2578_ ;
wire _2158_ ;
wire _0_ ;
wire [31:0] \preg[7]  ;
wire _1849_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _2387_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _2196_ ;
wire _41_ ;
wire _1887_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire areg_1_bF$buf0 ;
wire areg_1_bF$buf1 ;
wire areg_1_bF$buf2 ;
wire areg_1_bF$buf3 ;
wire areg_1_bF$buf4 ;
wire _2502_ ;
wire _2099_ ;
wire _2731_ ;
wire _2311_ ;
wire _913_ ;
wire _1599_ ;
wire _1179_ ;
wire _2540_ ;
wire _2120_ ;
wire _1811_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _2405_ ;
wire _760_ ;
wire _340_ ;
wire _2634_ ;
wire _2214_ ;
wire _1905_ ;
wire _816_ ;
wire _76_ ;
wire _2443_ ;
wire _2023_ ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire _2672_ ;
wire _2252_ ;
wire _1943_ ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _2728_ ;
wire _2308_ ;
wire _2481_ ;
wire _2061_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _2537_ ;
wire _2117_ ;
wire _2290_ ;
wire _1808_ ;
wire _719_ ;
wire _1981_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _2346_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1790_ ;
wire _1370_ ;
wire _281_ ;
wire _2575_ ;
wire _2155_ ;
wire _1846_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _2384_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _2193_ ;
wire _1884_ ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _2669_ ;
wire _2249_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _2478_ ;
wire _2058_ ;
wire _1749_ ;
wire _1329_ ;
wire _1082_ ;
wire _2287_ ;
wire _1978_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _2096_ ;
wire _1787_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire aregp1_13_bF$buf0 ;
wire aregp1_13_bF$buf1 ;
wire aregp1_13_bF$buf2 ;
wire aregp1_13_bF$buf3 ;
wire _35_ ;
wire _2402_ ;
wire _2631_ ;
wire _2211_ ;
wire _1902_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _2440_ ;
wire _2020_ ;
wire _1711_ ;
wire _622_ ;
wire _202_ ;
wire _1940_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _2725_ ;
wire _2305_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _2534_ ;
wire _2114_ ;
wire _1805_ ;
wire _716_ ;
wire _2343_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _2572_ ;
wire _2152_ ;
wire _1843_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _2628_ ;
wire _2208_ ;
wire _2381_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _2437_ ;
wire _2017_ ;
wire _2190_ ;
wire _1708_ ;
wire _619_ ;
wire _1881_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _2666_ ;
wire _2246_ ;
wire _1937_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _2475_ ;
wire _2055_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _2284_ ;
wire _1975_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _2093_ ;
wire _1784_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _2569_ ;
wire _2149_ ;
wire _1593_ ;
wire _1173_ ;
wire _2378_ ;
wire _1649_ ;
wire _1229_ ;
wire _2187_ ;
wire _32_ ;
wire _1878_ ;
wire _1458_ ;
wire _1038_ ;
wire _789_ ;
wire _369_ ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _2722_ ;
wire _2302_ ;
wire _904_ ;
wire _2531_ ;
wire _2111_ ;
wire _1802_ ;
wire _713_ ;
wire _1399_ ;
wire _2340_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1840_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _2625_ ;
wire _2205_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _2434_ ;
wire _2014_ ;
wire _1705_ ;
wire _616_ ;
wire _2663_ ;
wire _2243_ ;
wire _1934_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _2719_ ;
wire _2472_ ;
wire _2052_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _2528_ ;
wire _2108_ ;
wire _2281_ ;
wire _1972_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _2337_ ;
wire _2090_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1781_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _2566_ ;
wire _2146_ ;
wire _1837_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _2375_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _2184_ ;
wire _1875_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _2469_ ;
wire _2049_ ;
wire _1493_ ;
wire _1073_ ;
wire _2698_ ;
wire _2278_ ;
wire _1969_ ;
wire _1549_ ;
wire _1129_ ;
wire _2087_ ;
wire _1778_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire [31:0] \partials[15]  ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire _2622_ ;
wire _2202_ ;
wire _804_ ;
wire _64_ ;
wire _2431_ ;
wire _2011_ ;
wire _1702_ ;
wire _613_ ;
wire _1299_ ;
wire _2660_ ;
wire _2240_ ;
wire _1931_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _2716_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _2525_ ;
wire _2105_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _2334_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _2563_ ;
wire _2143_ ;
wire _1834_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _2619_ ;
wire _2372_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _2428_ ;
wire _2008_ ;
wire _2181_ ;
wire _1872_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _2657_ ;
wire _2237_ ;
wire _1928_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire [15:0] bregp1 ;
wire _592_ ;
wire _172_ ;
wire _2466_ ;
wire _2046_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _2695_ ;
wire _2275_ ;
wire _1966_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _2084_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _2369_ ;
wire _1393_ ;
wire _2598_ ;
wire _2178_ ;
wire _23_ ;
wire _1869_ ;
wire _1449_ ;
wire _1029_ ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _2713_ ;
wire _2522_ ;
wire _2102_ ;
wire _704_ ;
wire _2331_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _2560_ ;
wire _2140_ ;
wire _1831_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _2616_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _2425_ ;
wire _2005_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _2654_ ;
wire _2234_ ;
wire _1925_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _2463_ ;
wire _2043_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _2519_ ;
wire _2692_ ;
wire _2272_ ;
wire _1963_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _2328_ ;
wire [15:0] \partials[0]  ;
wire _2081_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _2557_ ;
wire _2137_ ;
wire _1828_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _2366_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _2595_ ;
wire _2175_ ;
wire _20_ ;
wire _1866_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _2689_ ;
wire _2269_ ;
wire _1293_ ;
wire _2498_ ;
wire _2078_ ;
wire _1769_ ;
wire _1349_ ;
wire _2710_ ;
wire _1998_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire _1196_ ;
wire _2613_ ;
wire _55_ ;
wire _2422_ ;
wire _2002_ ;
wire _604_ ;
wire _2651_ ;
wire _2231_ ;
wire _1922_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _2707_ ;
wire _93_ ;
wire _1099_ ;
wire _2460_ ;
wire _2040_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _2516_ ;
wire _1960_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _2325_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _2554_ ;
wire _2134_ ;
wire _1825_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _2363_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _2419_ ;
wire _2592_ ;
wire _2172_ ;
wire _1863_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _2648_ ;
wire _2228_ ;
wire _1919_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _2457_ ;
wire _2037_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _2686_ ;
wire _2266_ ;
wire _1957_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _2495_ ;
wire _2075_ ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1995_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _2589_ ;
wire _2169_ ;
wire _14_ ;
wire _1193_ ;
wire _2398_ ;
wire [31:0] \partials[7]  ;
wire _1669_ ;
wire _1249_ ;
wire _2610_ ;
wire _52_ ;
wire _1898_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _2704_ ;
wire _90_ ;
wire _1096_ ;
wire _2513_ ;
wire _2742_ ;
wire _2322_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _2551_ ;
wire _2131_ ;
wire _1822_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _2607_ ;
wire _2360_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _2416_ ;
wire _1860_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _2645_ ;
wire _2225_ ;
wire _1916_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _2454_ ;
wire _2034_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _2683_ ;
wire _2263_ ;
wire _1954_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _2739_ ;
wire _2319_ ;
wire _2492_ ;
wire _2072_ ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _2548_ ;
wire _2128_ ;
wire _1819_ ;
wire _1992_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _2357_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _2586_ ;
wire _2166_ ;
wire _11_ ;
wire _1857_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _2395_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1895_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _2489_ ;
wire _2069_ ;
wire _2701_ ;
wire _1093_ ;
wire _2298_ ;
wire _1989_ ;
wire _1569_ ;
wire _1149_ ;
wire _2510_ ;
wire aregp1_10_bF$buf0 ;
wire aregp1_10_bF$buf1 ;
wire aregp1_10_bF$buf2 ;
wire aregp1_10_bF$buf3 ;
wire _1798_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _2604_ ;
wire _46_ ;
wire _2413_ ;
wire _2642_ ;
wire _2222_ ;
wire _1913_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _2451_ ;
wire _2031_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _2507_ ;
wire _2680_ ;
wire _2260_ ;
wire _1951_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _2736_ ;
wire _2316_ ;
wire _918_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _2545_ ;
wire _2125_ ;
wire _1816_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _2354_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _2583_ ;
wire _2163_ ;
wire _1854_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _2639_ ;
wire _2219_ ;
wire _2392_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _2448_ ;
wire _2028_ ;
wire _1719_ ;
wire _1892_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _2677_ ;
wire _2257_ ;
wire _1948_ ;
wire _1528_ ;
wire _1108_ ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _2486_ ;
wire _2066_ ;
wire _1757_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _2295_ ;
wire _1986_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1795_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _2389_ ;
wire _2601_ ;
wire _2198_ ;
wire _43_ ;
wire _1889_ ;
wire _1469_ ;
wire _1049_ ;
wire _2410_ ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _1910_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire _630_ ;
wire _210_ ;
wire _2504_ ;
wire _2733_ ;
wire _2313_ ;
wire _915_ ;
wire _2542_ ;
wire _2122_ ;
wire _1813_ ;
wire _724_ ;
wire _304_ ;
wire _2351_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _2407_ ;
wire _2580_ ;
wire _2160_ ;
wire _1851_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _2636_ ;
wire _2216_ ;
wire _1907_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _2445_ ;
wire _2025_ ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _2674_ ;
wire _2254_ ;
wire _1945_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _2483_ ;
wire _2063_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _2539_ ;
wire _2119_ ;
wire _2292_ ;
wire _1983_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _2348_ ;
wire _1619_ ;
wire _1792_ ;
wire _1372_ ;
wire _283_ ;
wire _2577_ ;
wire _2157_ ;
wire _1848_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _2386_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _2195_ ;
wire _40_ ;
wire _1886_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire aregp1_8_bF$buf0 ;
wire aregp1_8_bF$buf1 ;
wire aregp1_8_bF$buf2 ;
wire aregp1_8_bF$buf3 ;
wire aregp1_8_bF$buf4 ;
wire _1084_ ;
wire _2289_ ;
wire _2501_ ;
wire _2098_ ;
wire _1789_ ;
wire _1369_ ;
wire _2730_ ;
wire _2310_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _1810_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _2404_ ;
wire _2633_ ;
wire _2213_ ;
wire _1904_ ;
wire _815_ ;
wire _75_ ;
wire _2442_ ;
wire _2022_ ;
wire _1713_ ;
wire _624_ ;
wire _204_ ;
wire _2671_ ;
wire _2251_ ;
wire _1942_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _2727_ ;
wire _2307_ ;
wire _2480_ ;
wire _2060_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _2536_ ;
wire _2116_ ;
wire _1807_ ;
wire _718_ ;
wire _1980_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _2345_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _2574_ ;
wire _2154_ ;
wire _1845_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _2383_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _2439_ ;
wire _2019_ ;
wire _2192_ ;
wire _1883_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _2668_ ;
wire _2248_ ;
wire _1939_ ;
wire _1519_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _2477_ ;
wire _2057_ ;
wire _1748_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _2286_ ;
wire _1977_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _2095_ ;
wire _1786_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _2189_ ;
wire _34_ ;
wire _2401_ ;
wire _1689_ ;
wire _1269_ ;
wire _2630_ ;
wire _2210_ ;
wire _1901_ ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _2724_ ;
wire _2304_ ;
wire _906_ ;
wire _2533_ ;
wire _2113_ ;
wire _1804_ ;
wire _715_ ;
wire _2342_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _2571_ ;
wire _2151_ ;
wire _1842_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _2627_ ;
wire _2207_ ;
wire _2380_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _2436_ ;
wire _2016_ ;
wire _1707_ ;
wire _618_ ;
wire _1880_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _2665_ ;
wire _2245_ ;
wire _1936_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _2474_ ;
wire _2054_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _2283_ ;
wire _1974_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _2339_ ;
wire _2092_ ;
wire areg_0_bF$buf0 ;
wire areg_0_bF$buf1 ;
wire areg_0_bF$buf2 ;
wire areg_0_bF$buf3 ;
wire areg_0_bF$buf4 ;
wire _1783_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _2568_ ;
wire _2148_ ;
wire _1839_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _2377_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _2186_ ;
wire _31_ ;
wire _1877_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _2089_ ;
wire _2721_ ;
wire _2301_ ;
wire _903_ ;
wire _1589_ ;
wire _1169_ ;
wire _2530_ ;
wire _2110_ ;
wire _1801_ ;
wire _712_ ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _2624_ ;
wire _2204_ ;
wire _806_ ;
wire _66_ ;
wire _2433_ ;
wire _2013_ ;
wire _1704_ ;
wire _615_ ;
wire _2662_ ;
wire _2242_ ;
wire _1933_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _2718_ ;
wire _2471_ ;
wire _2051_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _2527_ ;
wire _2107_ ;
wire _2280_ ;
wire _709_ ;
wire _1971_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _2336_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1780_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _2565_ ;
wire _2145_ ;
wire _1836_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _2374_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _2183_ ;
wire _1874_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _2659_ ;
wire _2239_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _2468_ ;
wire _2048_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire _2697_ ;
wire _2277_ ;
wire _1968_ ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _2086_ ;
wire _1777_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _2621_ ;
wire _2201_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _2430_ ;
wire _2010_ ;
wire _1701_ ;
wire _612_ ;
wire _1298_ ;
wire _1930_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _2715_ ;
wire _650_ ;
wire _230_ ;
wire _2524_ ;
wire _2104_ ;
wire _706_ ;
wire _2333_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _2562_ ;
wire _2142_ ;
wire _1833_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _2618_ ;
wire _2371_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _2427_ ;
wire _2007_ ;
wire _2180_ ;
wire _609_ ;
wire _1871_ ;
wire _1451_ ;
wire _1031_ ;
wire [15:0] aregp1 ;
wire _782_ ;
wire _362_ ;
wire _2656_ ;
wire _2236_ ;
wire _1927_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _2465_ ;
wire _2045_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _2694_ ;
wire _2274_ ;
wire _1965_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _2083_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _2559_ ;
wire _2139_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _2368_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _2597_ ;
wire _2177_ ;
wire _22_ ;
wire _1868_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert48 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[10]),
    .Y(aregp1_10_bF$buf0)
);

BUFX2 BUFX2_insert47 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[10]),
    .Y(aregp1_10_bF$buf1)
);

BUFX2 BUFX2_insert46 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[10]),
    .Y(aregp1_10_bF$buf2)
);

BUFX2 BUFX2_insert45 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[10]),
    .Y(aregp1_10_bF$buf3)
);

BUFX2 BUFX2_insert44 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf0)
);

BUFX2 BUFX2_insert43 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf1)
);

BUFX2 BUFX2_insert42 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf2)
);

BUFX2 BUFX2_insert41 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf3)
);

BUFX2 BUFX2_insert40 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[0]),
    .Y(areg_0_bF$buf4)
);

BUFX2 BUFX2_insert39 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[13]),
    .Y(aregp1_13_bF$buf0)
);

BUFX2 BUFX2_insert38 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[13]),
    .Y(aregp1_13_bF$buf1)
);

BUFX2 BUFX2_insert37 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[13]),
    .Y(aregp1_13_bF$buf2)
);

BUFX2 BUFX2_insert36 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[13]),
    .Y(aregp1_13_bF$buf3)
);

BUFX2 BUFX2_insert35 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf0)
);

BUFX2 BUFX2_insert34 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf1)
);

BUFX2 BUFX2_insert33 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf2)
);

BUFX2 BUFX2_insert32 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[6]),
    .Y(areg_6_bF$buf3)
);

BUFX2 BUFX2_insert31 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[8]),
    .Y(aregp1_8_bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[8]),
    .Y(aregp1_8_bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[8]),
    .Y(aregp1_8_bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[8]),
    .Y(aregp1_8_bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[8]),
    .Y(aregp1_8_bF$buf4)
);

CLKBUF1 CLKBUF1_insert26 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert25 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert24 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert23 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert22 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert21 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert20 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert19 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert18 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert17 (
    .gnd(gnd),
    .vdd(vdd),
    .A(clk),
    .Y(clk_bF$buf9)
);

BUFX2 BUFX2_insert16 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[11]),
    .Y(aregp1_11_bF$buf0)
);

BUFX2 BUFX2_insert15 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[11]),
    .Y(aregp1_11_bF$buf1)
);

BUFX2 BUFX2_insert14 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[11]),
    .Y(aregp1_11_bF$buf2)
);

BUFX2 BUFX2_insert13 (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[11]),
    .Y(aregp1_11_bF$buf3)
);

BUFX2 BUFX2_insert12 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf1)
);

BUFX2 BUFX2_insert10 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[1]),
    .Y(areg_1_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[4]),
    .Y(areg_4_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf0)
);

BUFX2 BUFX2_insert2 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf1)
);

BUFX2 BUFX2_insert1 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf2)
);

BUFX2 BUFX2_insert0 (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[7]),
    .Y(areg_7_bF$buf3)
);

INVX4 _2745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .Y(_129_)
);

INVX2 _2746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .Y(_140_)
);

NOR2X1 _2747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_140_),
    .Y(\partials[0] [0])
);

INVX1 _2748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .Y(_160_)
);

INVX4 _2749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[0]),
    .Y(_171_)
);

NOR2X1 _2750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_171_),
    .Y(_182_)
);

NAND2X1 _2751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\preg[7] [8]),
    .B(_182_),
    .Y(_193_)
);

INVX2 _2752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_193_),
    .Y(_204_)
);

NOR2X1 _2753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\preg[7] [8]),
    .B(_182_),
    .Y(_215_)
);

NOR2X1 _2754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_215_),
    .B(_204_),
    .Y(\partials[15] [8])
);

INVX1 _2755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .Y(_236_)
);

NOR2X1 _2756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_236_),
    .Y(_246_)
);

NAND3X1 _2757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[1]),
    .C(\preg[7] [9]),
    .Y(_257_)
);

INVX2 _2758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .Y(_268_)
);

INVX1 _2759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(\preg[7] [9]),
    .Y(_279_)
);

OAI21X1 _2760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_160_),
    .B(_268_),
    .C(_279_),
    .Y(_290_)
);

NAND2X1 _2761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_257_),
    .B(_290_),
    .Y(_301_)
);

XNOR2X1 _2762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_301_),
    .B(_246_),
    .Y(_312_)
);

NAND2X1 _2763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_312_),
    .Y(_323_)
);

INVX1 _2764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_323_),
    .Y(_343_)
);

NOR2X1 _2765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_204_),
    .B(_312_),
    .Y(_344_)
);

NOR2X1 _2766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_344_),
    .B(_343_),
    .Y(\partials[15] [9])
);

INVX4 _2767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf3),
    .Y(_365_)
);

NOR2X1 _2768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_365_),
    .Y(_376_)
);

INVX1 _2769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .Y(_386_)
);

INVX1 _2770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_246_),
    .Y(_397_)
);

OAI21X1 _2771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_301_),
    .B(_397_),
    .C(_257_),
    .Y(_408_)
);

NAND2X1 _2772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .B(aregp1[9]),
    .Y(_419_)
);

NAND3X1 _2773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[2]),
    .C(\preg[7] [10]),
    .Y(_430_)
);

AOI21X1 _2774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[2]),
    .C(\preg[7] [10]),
    .Y(_441_)
);

INVX1 _2775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .Y(_452_)
);

NAND2X1 _2776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_452_),
    .Y(_462_)
);

NOR2X1 _2777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .B(_462_),
    .Y(_473_)
);

INVX1 _2778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_419_),
    .Y(_494_)
);

AOI21X1 _2779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_430_),
    .B(_452_),
    .C(_494_),
    .Y(_505_)
);

NOR2X1 _2780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_505_),
    .B(_473_),
    .Y(_506_)
);

NAND2X1 _2781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_506_),
    .Y(_526_)
);

INVX1 _2782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .Y(_527_)
);

OAI21X1 _2783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_473_),
    .B(_505_),
    .C(_527_),
    .Y(_538_)
);

NAND3X1 _2784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_386_),
    .B(_538_),
    .C(_526_),
    .Y(_549_)
);

XNOR2X1 _2785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_462_),
    .B(_419_),
    .Y(_560_)
);

NOR2X1 _2786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_560_),
    .B(_527_),
    .Y(_570_)
);

NOR2X1 _2787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_408_),
    .B(_506_),
    .Y(_581_)
);

OAI21X1 _2788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_570_),
    .C(_376_),
    .Y(_591_)
);

AOI21X1 _2789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_591_),
    .C(_323_),
    .Y(_602_)
);

NAND2X1 _2790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_549_),
    .B(_591_),
    .Y(_612_)
);

NOR2X1 _2791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_343_),
    .B(_612_),
    .Y(_621_)
);

NOR2X1 _2792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_602_),
    .B(_621_),
    .Y(\partials[15] [10])
);

OAI21X1 _2793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_581_),
    .B(_386_),
    .C(_526_),
    .Y(_641_)
);

INVX2 _2794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf3),
    .Y(_652_)
);

NOR2X1 _2795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_652_),
    .Y(_662_)
);

NAND2X1 _2796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_662_),
    .Y(_673_)
);

NAND2X1 _2797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .B(aregp1_10_bF$buf2),
    .Y(_684_)
);

OAI21X1 _2798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_652_),
    .C(_684_),
    .Y(_695_)
);

NAND2X1 _2799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_695_),
    .B(_673_),
    .Y(_705_)
);

OAI21X1 _2800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_441_),
    .B(_419_),
    .C(_430_),
    .Y(_716_)
);

NAND2X1 _2801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[2]),
    .Y(_727_)
);

INVX1 _2802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .Y(_738_)
);

NAND3X1 _2803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[3]),
    .C(\preg[7] [11]),
    .Y(_758_)
);

AOI21X1 _2804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .B(bregp1[3]),
    .C(\preg[7] [11]),
    .Y(_759_)
);

INVX1 _2805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .Y(_770_)
);

NAND3X1 _2806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_738_),
    .B(_758_),
    .C(_770_),
    .Y(_781_)
);

INVX1 _2807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_),
    .Y(_792_)
);

OAI21X1 _2808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_792_),
    .B(_759_),
    .C(_727_),
    .Y(_803_)
);

NAND3X1 _2809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .B(_781_),
    .C(_803_),
    .Y(_814_)
);

INVX1 _2810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_716_),
    .Y(_825_)
);

NOR3X1 _2811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_727_),
    .B(_759_),
    .C(_792_),
    .Y(_835_)
);

AOI21X1 _2812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_758_),
    .B(_770_),
    .C(_738_),
    .Y(_846_)
);

OAI21X1 _2813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_835_),
    .B(_846_),
    .C(_825_),
    .Y(_857_)
);

NAND2X1 _2814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .B(_857_),
    .Y(_868_)
);

NOR2X1 _2815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .B(_868_),
    .Y(_879_)
);

INVX1 _2816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_879_),
    .Y(_890_)
);

INVX1 _2817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_814_),
    .Y(_901_)
);

AOI21X1 _2818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_781_),
    .B(_803_),
    .C(_716_),
    .Y(_912_)
);

OAI21X1 _2819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_901_),
    .B(_912_),
    .C(_705_),
    .Y(_922_)
);

NAND3X1 _2820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .B(_890_),
    .C(_641_),
    .Y(_933_)
);

AOI21X1 _2821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_376_),
    .B(_538_),
    .C(_570_),
    .Y(_944_)
);

INVX1 _2822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_922_),
    .Y(_955_)
);

OAI21X1 _2823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_879_),
    .C(_944_),
    .Y(_976_)
);

NAND3X1 _2824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(_933_),
    .C(_602_),
    .Y(_987_)
);

INVX1 _2825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_987_),
    .Y(_988_)
);

AOI21X1 _2826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_976_),
    .B(_933_),
    .C(_602_),
    .Y(_1009_)
);

NOR2X1 _2827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1009_),
    .B(_988_),
    .Y(\partials[15] [11])
);

INVX2 _2828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .Y(_1019_)
);

OAI21X1 _2829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_912_),
    .B(_705_),
    .C(_814_),
    .Y(_1030_)
);

NAND2X1 _2830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[0]),
    .B(aregp1[12]),
    .Y(_1041_)
);

NAND2X1 _2831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[2]),
    .B(aregp1_11_bF$buf2),
    .Y(_1052_)
);

NOR2X1 _2832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_1052_),
    .Y(_1063_)
);

AOI22X1 _2833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .B(aregp1_11_bF$buf1),
    .C(bregp1[2]),
    .D(aregp1_10_bF$buf1),
    .Y(_1074_)
);

NOR2X1 _2834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1074_),
    .B(_1063_),
    .Y(_1085_)
);

XNOR2X1 _2835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_1041_),
    .Y(_1096_)
);

OAI21X1 _2836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_759_),
    .B(_727_),
    .C(_758_),
    .Y(_1107_)
);

NAND2X1 _2837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[3]),
    .Y(_1117_)
);

INVX1 _2838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1117_),
    .Y(_1128_)
);

NAND3X1 _2839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[4]),
    .C(\preg[7] [12]),
    .Y(_1139_)
);

AOI21X1 _2840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[4]),
    .C(\preg[7] [12]),
    .Y(_1150_)
);

INVX1 _2841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .Y(_1161_)
);

NAND3X1 _2842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1128_),
    .B(_1139_),
    .C(_1161_),
    .Y(_1172_)
);

INVX1 _2843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .Y(_1183_)
);

OAI21X1 _2844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1183_),
    .B(_1150_),
    .C(_1117_),
    .Y(_1194_)
);

NAND3X1 _2845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1107_),
    .B(_1172_),
    .C(_1194_),
    .Y(_1205_)
);

INVX1 _2846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1107_),
    .Y(_1216_)
);

NOR3X1 _2847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1117_),
    .B(_1150_),
    .C(_1183_),
    .Y(_1226_)
);

AOI21X1 _2848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1139_),
    .B(_1161_),
    .C(_1128_),
    .Y(_1237_)
);

OAI21X1 _2849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1237_),
    .C(_1216_),
    .Y(_1248_)
);

NAND3X1 _2850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1248_),
    .C(_1096_),
    .Y(_1259_)
);

XOR2X1 _2851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1085_),
    .B(_1041_),
    .Y(_1270_)
);

INVX1 _2852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .Y(_1281_)
);

AOI21X1 _2853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1172_),
    .B(_1194_),
    .C(_1107_),
    .Y(_1292_)
);

OAI21X1 _2854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1281_),
    .B(_1292_),
    .C(_1270_),
    .Y(_1303_)
);

NAND3X1 _2855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1030_),
    .B(_1259_),
    .C(_1303_),
    .Y(_1314_)
);

INVX1 _2856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_705_),
    .Y(_1324_)
);

AOI21X1 _2857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1324_),
    .B(_857_),
    .C(_901_),
    .Y(_1335_)
);

OAI21X1 _2858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1226_),
    .B(_1237_),
    .C(_1107_),
    .Y(_1346_)
);

NAND3X1 _2859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1172_),
    .B(_1194_),
    .C(_1216_),
    .Y(_1357_)
);

AOI21X1 _2860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1346_),
    .B(_1357_),
    .C(_1270_),
    .Y(_1368_)
);

AOI21X1 _2861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1205_),
    .B(_1248_),
    .C(_1096_),
    .Y(_1379_)
);

OAI21X1 _2862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1368_),
    .B(_1379_),
    .C(_1335_),
    .Y(_1390_)
);

NAND3X1 _2863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(_1390_),
    .C(_1314_),
    .Y(_1401_)
);

OAI21X1 _2864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1368_),
    .B(_1379_),
    .C(_1030_),
    .Y(_1412_)
);

NAND3X1 _2865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1335_),
    .B(_1259_),
    .C(_1303_),
    .Y(_1422_)
);

NAND3X1 _2866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_1412_),
    .C(_1422_),
    .Y(_1433_)
);

NAND2X1 _2867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1401_),
    .B(_1433_),
    .Y(_1444_)
);

NAND2X1 _2868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_933_),
    .B(_987_),
    .Y(_1455_)
);

XNOR2X1 _2869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1455_),
    .B(_1444_),
    .Y(\partials[15] [12])
);

NOR2X1 _2870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1444_),
    .B(_987_),
    .Y(_1476_)
);

INVX2 _2871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .Y(_1497_)
);

NOR3X1 _2872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_955_),
    .B(_879_),
    .C(_944_),
    .Y(_1508_)
);

NAND3X1 _2873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1401_),
    .B(_1508_),
    .C(_1433_),
    .Y(_1509_)
);

AOI21X1 _2874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1259_),
    .B(_1303_),
    .C(_1030_),
    .Y(_1529_)
);

OAI21X1 _2875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1529_),
    .B(_673_),
    .C(_1314_),
    .Y(_1530_)
);

NAND2X1 _2876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[0]),
    .B(aregp1_13_bF$buf3),
    .Y(_1541_)
);

INVX1 _2877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .Y(_1552_)
);

OAI22X1 _2878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_684_),
    .B(_1052_),
    .C(_1074_),
    .D(_1041_),
    .Y(_1563_)
);

NAND2X1 _2879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_1563_),
    .Y(_1574_)
);

INVX2 _2880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .Y(_1585_)
);

NOR2X1 _2881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1552_),
    .B(_1563_),
    .Y(_1596_)
);

NOR2X1 _2882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1596_),
    .B(_1585_),
    .Y(_1606_)
);

INVX2 _2883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .Y(_1617_)
);

OAI21X1 _2884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1270_),
    .B(_1292_),
    .C(_1205_),
    .Y(_1628_)
);

INVX4 _2885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .Y(_1639_)
);

NOR2X1 _2886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_1639_),
    .Y(_1650_)
);

NAND3X1 _2887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf0),
    .B(bregp1[3]),
    .C(_1052_),
    .Y(_1661_)
);

NAND2X1 _2888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf3),
    .B(bregp1[3]),
    .Y(_1672_)
);

NAND3X1 _2889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[2]),
    .B(aregp1_11_bF$buf0),
    .C(_1672_),
    .Y(_1683_)
);

NAND2X1 _2890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1661_),
    .B(_1683_),
    .Y(_1693_)
);

XNOR2X1 _2891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1693_),
    .B(_1650_),
    .Y(_1704_)
);

OAI21X1 _2892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1150_),
    .B(_1117_),
    .C(_1139_),
    .Y(_1715_)
);

NAND2X1 _2893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[4]),
    .Y(_1726_)
);

NAND3X1 _2894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[5]),
    .C(\preg[7] [13]),
    .Y(_1737_)
);

INVX1 _2895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1737_),
    .Y(_1748_)
);

AOI21X1 _2896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[5]),
    .C(\preg[7] [13]),
    .Y(_1759_)
);

NOR3X1 _2897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .B(_1759_),
    .C(_1748_),
    .Y(_1770_)
);

INVX1 _2898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1726_),
    .Y(_1780_)
);

INVX1 _2899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1759_),
    .Y(_1791_)
);

AOI21X1 _2900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1737_),
    .B(_1791_),
    .C(_1780_),
    .Y(_1802_)
);

OAI21X1 _2901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(_1802_),
    .C(_1715_),
    .Y(_1813_)
);

INVX2 _2902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1715_),
    .Y(_1824_)
);

NAND3X1 _2903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1780_),
    .B(_1737_),
    .C(_1791_),
    .Y(_1835_)
);

OAI21X1 _2904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1748_),
    .B(_1759_),
    .C(_1726_),
    .Y(_1846_)
);

NAND3X1 _2905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(_1846_),
    .C(_1824_),
    .Y(_1856_)
);

AOI21X1 _2906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1813_),
    .B(_1856_),
    .C(_1704_),
    .Y(_1867_)
);

INVX2 _2907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1650_),
    .Y(_1878_)
);

XNOR2X1 _2908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1693_),
    .B(_1878_),
    .Y(_1889_)
);

NAND3X1 _2909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1715_),
    .B(_1835_),
    .C(_1846_),
    .Y(_1900_)
);

OAI21X1 _2910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1770_),
    .B(_1802_),
    .C(_1824_),
    .Y(_1910_)
);

AOI21X1 _2911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .B(_1910_),
    .C(_1889_),
    .Y(_1921_)
);

OAI21X1 _2912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1921_),
    .C(_1628_),
    .Y(_1932_)
);

AOI21X1 _2913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1248_),
    .B(_1096_),
    .C(_1281_),
    .Y(_1943_)
);

NAND3X1 _2914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1900_),
    .B(_1910_),
    .C(_1889_),
    .Y(_1954_)
);

NOR3X1 _2915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1802_),
    .B(_1824_),
    .C(_1770_),
    .Y(_1965_)
);

AOI21X1 _2916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1835_),
    .B(_1846_),
    .C(_1715_),
    .Y(_1975_)
);

OAI21X1 _2917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1965_),
    .B(_1975_),
    .C(_1704_),
    .Y(_1995_)
);

NAND3X1 _2918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(_1995_),
    .C(_1943_),
    .Y(_2006_)
);

AOI21X1 _2919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1932_),
    .B(_2006_),
    .C(_1617_),
    .Y(_2007_)
);

NAND3X1 _2920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(_1995_),
    .C(_1628_),
    .Y(_2027_)
);

OAI21X1 _2921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1921_),
    .C(_1943_),
    .Y(_2028_)
);

AOI21X1 _2922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2028_),
    .B(_2027_),
    .C(_1606_),
    .Y(_2039_)
);

OAI21X1 _2923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2039_),
    .B(_2007_),
    .C(_1530_),
    .Y(_2043_)
);

NOR3X1 _2924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1368_),
    .B(_1379_),
    .C(_1335_),
    .Y(_2044_)
);

AOI21X1 _2925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1019_),
    .B(_1390_),
    .C(_2044_),
    .Y(_2045_)
);

NAND3X1 _2926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(_2028_),
    .C(_2027_),
    .Y(_2046_)
);

NAND3X1 _2927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1617_),
    .B(_1932_),
    .C(_2006_),
    .Y(_2047_)
);

NAND3X1 _2928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2046_),
    .B(_2047_),
    .C(_2045_),
    .Y(_2048_)
);

AOI21X1 _2929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2048_),
    .B(_2043_),
    .C(_1509_),
    .Y(_2049_)
);

NAND3X1 _2930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_673_),
    .B(_1390_),
    .C(_1314_),
    .Y(_2050_)
);

OAI21X1 _2931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2044_),
    .B(_1529_),
    .C(_1019_),
    .Y(_2051_)
);

NAND2X1 _2932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2050_),
    .B(_2051_),
    .Y(_2052_)
);

NAND3X1 _2933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2047_),
    .B(_2046_),
    .C(_1530_),
    .Y(_2053_)
);

OAI21X1 _2934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2039_),
    .B(_2007_),
    .C(_2045_),
    .Y(_2054_)
);

AOI22X1 _2935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1508_),
    .B(_2052_),
    .C(_2054_),
    .D(_2053_),
    .Y(_2055_)
);

NOR2X1 _2936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .B(_2055_),
    .Y(_2056_)
);

XNOR2X1 _2937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2056_),
    .B(_1497_),
    .Y(\partials[15] [13])
);

INVX1 _2938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2049_),
    .Y(_2057_)
);

OAI21X1 _2939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1497_),
    .B(_2055_),
    .C(_2057_),
    .Y(_2058_)
);

INVX1 _2940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .Y(_2059_)
);

AOI21X1 _2941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1954_),
    .B(_1995_),
    .C(_1628_),
    .Y(_2060_)
);

OAI21X1 _2942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2060_),
    .B(_1617_),
    .C(_2027_),
    .Y(_2061_)
);

NAND2X1 _2943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .B(aregp1[14]),
    .Y(_2062_)
);

NOR2X1 _2944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1541_),
    .B(_2062_),
    .Y(_2063_)
);

INVX2 _2945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2063_),
    .Y(_2064_)
);

INVX4 _2946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .Y(_2065_)
);

NAND2X1 _2947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[1]),
    .B(aregp1_13_bF$buf2),
    .Y(_2066_)
);

OAI21X1 _2948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_2065_),
    .C(_2066_),
    .Y(_2067_)
);

AND2X2 _2949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2067_),
    .Y(_2068_)
);

OR2X2 _2950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .B(_1672_),
    .Y(_2069_)
);

AND2X2 _2951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1052_),
    .B(_1672_),
    .Y(_2070_)
);

OAI21X1 _2952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1878_),
    .B(_2070_),
    .C(_2069_),
    .Y(_2071_)
);

NAND2X1 _2953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(_2068_),
    .Y(_2072_)
);

INVX2 _2954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2072_),
    .Y(_2073_)
);

NOR2X1 _2955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2071_),
    .B(_2068_),
    .Y(_2074_)
);

NOR2X1 _2956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2074_),
    .B(_2073_),
    .Y(_2075_)
);

OAI21X1 _2957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1704_),
    .B(_1975_),
    .C(_1900_),
    .Y(_2076_)
);

INVX2 _2958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[2]),
    .Y(_2077_)
);

NOR2X1 _2959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_1639_),
    .Y(_2078_)
);

NAND2X1 _2960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf3),
    .B(bregp1[4]),
    .Y(_2079_)
);

INVX2 _2961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[4]),
    .Y(_2080_)
);

NAND2X1 _2962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[3]),
    .B(aregp1_11_bF$buf2),
    .Y(_2081_)
);

OAI21X1 _2963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2080_),
    .C(_2081_),
    .Y(_2082_)
);

OAI21X1 _2964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1672_),
    .B(_2079_),
    .C(_2082_),
    .Y(_2083_)
);

XNOR2X1 _2965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2083_),
    .B(_2078_),
    .Y(_2084_)
);

OAI21X1 _2966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1759_),
    .B(_1726_),
    .C(_1737_),
    .Y(_2085_)
);

NAND2X1 _2967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[5]),
    .Y(_2086_)
);

INVX1 _2968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2086_),
    .Y(_2087_)
);

NAND3X1 _2969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .B(bregp1[6]),
    .C(\preg[7] [14]),
    .Y(_2088_)
);

AOI21X1 _2970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[6]),
    .C(\preg[7] [14]),
    .Y(_2089_)
);

INVX1 _2971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .Y(_2090_)
);

NAND3X1 _2972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2087_),
    .B(_2088_),
    .C(_2090_),
    .Y(_2091_)
);

INVX1 _2973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2088_),
    .Y(_2092_)
);

OAI21X1 _2974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2092_),
    .B(_2089_),
    .C(_2086_),
    .Y(_2093_)
);

NAND3X1 _2975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .B(_2091_),
    .C(_2093_),
    .Y(_2094_)
);

INVX1 _2976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2085_),
    .Y(_2095_)
);

NOR3X1 _2977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2086_),
    .B(_2089_),
    .C(_2092_),
    .Y(_2096_)
);

AOI21X1 _2978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2088_),
    .B(_2090_),
    .C(_2087_),
    .Y(_2097_)
);

OAI21X1 _2979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_2097_),
    .C(_2095_),
    .Y(_2098_)
);

NAND3X1 _2980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .B(_2098_),
    .C(_2084_),
    .Y(_2099_)
);

INVX1 _2981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2078_),
    .Y(_2100_)
);

XNOR2X1 _2982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2083_),
    .B(_2100_),
    .Y(_2101_)
);

OAI21X1 _2983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2096_),
    .B(_2097_),
    .C(_2085_),
    .Y(_2102_)
);

NAND3X1 _2984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2093_),
    .C(_2095_),
    .Y(_2103_)
);

NAND3X1 _2985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2102_),
    .B(_2103_),
    .C(_2101_),
    .Y(_2104_)
);

NAND3X1 _2986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_2104_),
    .C(_2076_),
    .Y(_2105_)
);

AOI21X1 _2987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1910_),
    .B(_1889_),
    .C(_1965_),
    .Y(_2106_)
);

AOI21X1 _2988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2102_),
    .B(_2103_),
    .C(_2101_),
    .Y(_2107_)
);

AOI21X1 _2989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .B(_2098_),
    .C(_2084_),
    .Y(_2108_)
);

OAI21X1 _2990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2108_),
    .C(_2106_),
    .Y(_2109_)
);

NAND3X1 _2991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2109_),
    .C(_2105_),
    .Y(_2110_)
);

OR2X2 _2992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2074_),
    .Y(_2111_)
);

OAI21X1 _2993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2108_),
    .C(_2076_),
    .Y(_2112_)
);

NAND3X1 _2994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_2104_),
    .C(_2106_),
    .Y(_2113_)
);

NAND3X1 _2995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2111_),
    .B(_2112_),
    .C(_2113_),
    .Y(_2114_)
);

NAND3X1 _2996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_2114_),
    .C(_2061_),
    .Y(_2115_)
);

NOR3X1 _2997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1867_),
    .B(_1921_),
    .C(_1943_),
    .Y(_2116_)
);

AOI21X1 _2998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1606_),
    .B(_2028_),
    .C(_2116_),
    .Y(_2117_)
);

AOI21X1 _2999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2112_),
    .B(_2113_),
    .C(_2111_),
    .Y(_2118_)
);

AOI21X1 _3000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2109_),
    .B(_2105_),
    .C(_2075_),
    .Y(_2119_)
);

OAI21X1 _3001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2118_),
    .B(_2119_),
    .C(_2117_),
    .Y(_2120_)
);

NAND3X1 _3002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_2115_),
    .C(_2120_),
    .Y(_2121_)
);

OAI21X1 _3003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2118_),
    .B(_2119_),
    .C(_2061_),
    .Y(_2122_)
);

NAND3X1 _3004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_2114_),
    .C(_2117_),
    .Y(_2123_)
);

NAND3X1 _3005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .B(_2122_),
    .C(_2123_),
    .Y(_2124_)
);

NAND3X1 _3006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2059_),
    .B(_2121_),
    .C(_2124_),
    .Y(_2125_)
);

NAND3X1 _3007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1574_),
    .B(_2115_),
    .C(_2120_),
    .Y(_2126_)
);

NAND3X1 _3008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1585_),
    .B(_2122_),
    .C(_2123_),
    .Y(_2127_)
);

NAND3X1 _3009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2053_),
    .B(_2126_),
    .C(_2127_),
    .Y(_2128_)
);

NAND3X1 _3010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2128_),
    .C(_2058_),
    .Y(_2129_)
);

NAND3X1 _3011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1509_),
    .B(_2048_),
    .C(_2043_),
    .Y(_2130_)
);

AOI21X1 _3012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1476_),
    .B(_2130_),
    .C(_2049_),
    .Y(_2131_)
);

AOI21X1 _3013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2126_),
    .B(_2127_),
    .C(_2053_),
    .Y(_2132_)
);

AOI21X1 _3014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2121_),
    .B(_2124_),
    .C(_2059_),
    .Y(_2133_)
);

OAI21X1 _3015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2132_),
    .B(_2133_),
    .C(_2131_),
    .Y(_2134_)
);

AND2X2 _3016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2129_),
    .B(_2134_),
    .Y(\partials[15] [14])
);

OAI21X1 _3017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2131_),
    .B(_2133_),
    .C(_2125_),
    .Y(_2135_)
);

AOI21X1 _3018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2110_),
    .B(_2114_),
    .C(_2061_),
    .Y(_2136_)
);

OAI21X1 _3019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2136_),
    .B(_1574_),
    .C(_2115_),
    .Y(_2137_)
);

AOI21X1 _3020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2099_),
    .B(_2104_),
    .C(_2076_),
    .Y(_2138_)
);

OAI21X1 _3021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2138_),
    .B(_2111_),
    .C(_2105_),
    .Y(_2139_)
);

NAND2X1 _3022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[0]),
    .B(aregp1[15]),
    .Y(_2140_)
);

NAND2X1 _3023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[2]),
    .B(aregp1[14]),
    .Y(_2141_)
);

INVX4 _3024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf1),
    .Y(_2142_)
);

OAI21X1 _3025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2142_),
    .C(_2062_),
    .Y(_2143_)
);

OAI21X1 _3026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2066_),
    .B(_2141_),
    .C(_2143_),
    .Y(_2144_)
);

OR2X2 _3027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .B(_2140_),
    .Y(_2145_)
);

INVX8 _3028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .Y(_2146_)
);

OAI21X1 _3029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_171_),
    .B(_2146_),
    .C(_2144_),
    .Y(_2147_)
);

NAND2X1 _3030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf2),
    .B(bregp1[4]),
    .Y(_2148_)
);

NOR2X1 _3031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2081_),
    .B(_2148_),
    .Y(_2149_)
);

AOI21X1 _3032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2078_),
    .B(_2082_),
    .C(_2149_),
    .Y(_2150_)
);

INVX1 _3033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2150_),
    .Y(_2151_)
);

NAND3X1 _3034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2151_),
    .B(_2147_),
    .C(_2145_),
    .Y(_2152_)
);

NOR2X1 _3035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2140_),
    .B(_2144_),
    .Y(_2153_)
);

AND2X2 _3036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2144_),
    .B(_2140_),
    .Y(_2154_)
);

OAI21X1 _3037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(_2153_),
    .C(_2150_),
    .Y(_2155_)
);

NAND3X1 _3038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2063_),
    .B(_2155_),
    .C(_2152_),
    .Y(_2156_)
);

NAND3X1 _3039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2150_),
    .B(_2147_),
    .C(_2145_),
    .Y(_2157_)
);

OAI21X1 _3040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2154_),
    .B(_2153_),
    .C(_2151_),
    .Y(_2158_)
);

NAND3X1 _3041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2158_),
    .C(_2157_),
    .Y(_2159_)
);

NAND2X1 _3042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2156_),
    .B(_2159_),
    .Y(_2160_)
);

AOI21X1 _3043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2091_),
    .B(_2093_),
    .C(_2085_),
    .Y(_2161_)
);

OAI21X1 _3044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2101_),
    .B(_2161_),
    .C(_2094_),
    .Y(_2162_)
);

INVX2 _3045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[3]),
    .Y(_2163_)
);

NOR2X1 _3046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_1639_),
    .Y(_2164_)
);

INVX1 _3047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .Y(_2165_)
);

NAND2X1 _3048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf1),
    .B(bregp1[5]),
    .Y(_2166_)
);

INVX2 _3049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[5]),
    .Y(_2167_)
);

OAI21X1 _3050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2167_),
    .C(_2079_),
    .Y(_2168_)
);

OAI21X1 _3051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2148_),
    .B(_2166_),
    .C(_2168_),
    .Y(_2169_)
);

XNOR2X1 _3052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2169_),
    .B(_2165_),
    .Y(_2170_)
);

OAI21X1 _3053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2089_),
    .B(_2086_),
    .C(_2088_),
    .Y(_2171_)
);

NAND2X1 _3054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[6]),
    .Y(_2172_)
);

NAND3X1 _3055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[7]),
    .C(\preg[7] [15]),
    .Y(_2173_)
);

INVX1 _3056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .Y(_2174_)
);

AOI21X1 _3057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[7]),
    .C(\preg[7] [15]),
    .Y(_2175_)
);

NOR3X1 _3058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .B(_2175_),
    .C(_2174_),
    .Y(_2176_)
);

INVX1 _3059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2172_),
    .Y(_2177_)
);

INVX1 _3060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2175_),
    .Y(_2178_)
);

AOI21X1 _3061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2173_),
    .B(_2178_),
    .C(_2177_),
    .Y(_2179_)
);

OAI21X1 _3062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .B(_2179_),
    .C(_2171_),
    .Y(_2180_)
);

INVX1 _3063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .Y(_2181_)
);

NAND3X1 _3064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2177_),
    .B(_2173_),
    .C(_2178_),
    .Y(_2182_)
);

OAI21X1 _3065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2174_),
    .B(_2175_),
    .C(_2172_),
    .Y(_2183_)
);

NAND3X1 _3066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2183_),
    .C(_2181_),
    .Y(_2184_)
);

AOI21X1 _3067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2180_),
    .B(_2184_),
    .C(_2170_),
    .Y(_2185_)
);

XNOR2X1 _3068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2169_),
    .B(_2164_),
    .Y(_2186_)
);

NAND3X1 _3069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2171_),
    .B(_2182_),
    .C(_2183_),
    .Y(_2187_)
);

OAI21X1 _3070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2176_),
    .B(_2179_),
    .C(_2181_),
    .Y(_2188_)
);

AOI21X1 _3071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .B(_2188_),
    .C(_2186_),
    .Y(_2189_)
);

OAI21X1 _3072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2189_),
    .C(_2162_),
    .Y(_2190_)
);

INVX1 _3073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2094_),
    .Y(_2191_)
);

AOI21X1 _3074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2098_),
    .B(_2084_),
    .C(_2191_),
    .Y(_2192_)
);

NAND3X1 _3075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .B(_2188_),
    .C(_2186_),
    .Y(_2193_)
);

INVX1 _3076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2187_),
    .Y(_2194_)
);

AOI21X1 _3077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2182_),
    .B(_2183_),
    .C(_2171_),
    .Y(_2195_)
);

OAI21X1 _3078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2194_),
    .B(_2195_),
    .C(_2170_),
    .Y(_2196_)
);

NAND3X1 _3079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2192_),
    .B(_2193_),
    .C(_2196_),
    .Y(_2197_)
);

AOI21X1 _3080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2190_),
    .B(_2197_),
    .C(_2160_),
    .Y(_2198_)
);

NAND3X1 _3081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2064_),
    .B(_2155_),
    .C(_2152_),
    .Y(_2199_)
);

NAND3X1 _3082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2063_),
    .B(_2158_),
    .C(_2157_),
    .Y(_2200_)
);

NAND2X1 _3083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2199_),
    .B(_2200_),
    .Y(_2201_)
);

NAND3X1 _3084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2162_),
    .B(_2193_),
    .C(_2196_),
    .Y(_2202_)
);

OAI21X1 _3085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2189_),
    .C(_2192_),
    .Y(_2203_)
);

AOI21X1 _3086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2202_),
    .B(_2203_),
    .C(_2201_),
    .Y(_2204_)
);

OAI21X1 _3087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2204_),
    .C(_2139_),
    .Y(_2205_)
);

NOR3X1 _3088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2107_),
    .B(_2108_),
    .C(_2106_),
    .Y(_2206_)
);

AOI21X1 _3089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2075_),
    .B(_2109_),
    .C(_2206_),
    .Y(_2207_)
);

NAND3X1 _3090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2202_),
    .B(_2203_),
    .C(_2201_),
    .Y(_2208_)
);

NOR3X1 _3091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2185_),
    .B(_2189_),
    .C(_2192_),
    .Y(_2209_)
);

AOI21X1 _3092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2193_),
    .B(_2196_),
    .C(_2162_),
    .Y(_2210_)
);

OAI21X1 _3093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2209_),
    .B(_2210_),
    .C(_2160_),
    .Y(_2211_)
);

NAND3X1 _3094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2207_),
    .B(_2208_),
    .C(_2211_),
    .Y(_2212_)
);

AOI21X1 _3095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2212_),
    .B(_2205_),
    .C(_2072_),
    .Y(_2213_)
);

NAND3X1 _3096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2139_),
    .B(_2208_),
    .C(_2211_),
    .Y(_2214_)
);

OAI21X1 _3097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2204_),
    .C(_2207_),
    .Y(_2215_)
);

AOI21X1 _3098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2214_),
    .B(_2215_),
    .C(_2073_),
    .Y(_2216_)
);

OAI21X1 _3099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2213_),
    .B(_2216_),
    .C(_2137_),
    .Y(_2217_)
);

INVX1 _3100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2137_),
    .Y(_2218_)
);

NAND3X1 _3101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2214_),
    .C(_2215_),
    .Y(_2219_)
);

NOR3X1 _3102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2198_),
    .B(_2207_),
    .C(_2204_),
    .Y(_2220_)
);

AOI21X1 _3103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2208_),
    .B(_2211_),
    .C(_2139_),
    .Y(_2221_)
);

OAI21X1 _3104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2220_),
    .B(_2221_),
    .C(_2072_),
    .Y(_2222_)
);

NAND3X1 _3105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2219_),
    .B(_2222_),
    .C(_2218_),
    .Y(_2223_)
);

NAND2X1 _3106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2217_),
    .B(_2223_),
    .Y(_2224_)
);

XOR2X1 _3107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .B(_2135_),
    .Y(\partials[15] [15])
);

NOR3X1 _3108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2132_),
    .B(_2133_),
    .C(_2131_),
    .Y(_2225_)
);

NAND3X1 _3109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2137_),
    .B(_2219_),
    .C(_2222_),
    .Y(_2226_)
);

AOI21X1 _3110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2219_),
    .B(_2222_),
    .C(_2137_),
    .Y(_2227_)
);

AOI21X1 _3111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2125_),
    .B(_2226_),
    .C(_2227_),
    .Y(_2228_)
);

AOI21X1 _3112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2224_),
    .B(_2225_),
    .C(_2228_),
    .Y(_2229_)
);

OAI21X1 _3113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2221_),
    .B(_2072_),
    .C(_2214_),
    .Y(_2230_)
);

NAND2X1 _3114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2152_),
    .B(_2156_),
    .Y(_2231_)
);

INVX2 _3115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .Y(_2232_)
);

OAI21X1 _3116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2160_),
    .B(_2210_),
    .C(_2202_),
    .Y(_2233_)
);

NAND2X1 _3117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[2]),
    .B(aregp1_13_bF$buf0),
    .Y(_2234_)
);

OAI21X1 _3118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2062_),
    .B(_2234_),
    .C(_2145_),
    .Y(_2235_)
);

NOR2X1 _3119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_2146_),
    .Y(_2236_)
);

NAND2X1 _3120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[3]),
    .B(aregp1_13_bF$buf3),
    .Y(_2237_)
);

OR2X2 _3121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2141_),
    .B(_2237_),
    .Y(_2238_)
);

OAI21X1 _3122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_2142_),
    .C(_2141_),
    .Y(_2239_)
);

NAND3X1 _3123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2236_),
    .B(_2239_),
    .C(_2238_),
    .Y(_2240_)
);

NAND2X1 _3124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[3]),
    .B(aregp1[14]),
    .Y(_2241_)
);

OAI21X1 _3125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2241_),
    .C(_2239_),
    .Y(_2242_)
);

OAI21X1 _3126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_268_),
    .B(_2146_),
    .C(_2242_),
    .Y(_2243_)
);

NAND2X1 _3127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf1),
    .B(bregp1[5]),
    .Y(_2244_)
);

NOR2X1 _3128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2079_),
    .B(_2244_),
    .Y(_2245_)
);

AOI21X1 _3129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2164_),
    .B(_2168_),
    .C(_2245_),
    .Y(_2246_)
);

INVX1 _3130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2246_),
    .Y(_2247_)
);

NAND3X1 _3131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2243_),
    .C(_2247_),
    .Y(_2248_)
);

INVX1 _3132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .Y(_2249_)
);

AOI21X1 _3133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2239_),
    .B(_2238_),
    .C(_2236_),
    .Y(_2250_)
);

OAI21X1 _3134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2249_),
    .B(_2250_),
    .C(_2246_),
    .Y(_2251_)
);

NAND3X1 _3135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2248_),
    .C(_2251_),
    .Y(_2252_)
);

NOR2X1 _3136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2062_),
    .B(_2234_),
    .Y(_2253_)
);

NOR2X1 _3137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2253_),
    .B(_2153_),
    .Y(_2254_)
);

NAND3X1 _3138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2240_),
    .B(_2246_),
    .C(_2243_),
    .Y(_2255_)
);

OAI21X1 _3139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2249_),
    .B(_2250_),
    .C(_2247_),
    .Y(_2256_)
);

NAND3X1 _3140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2255_),
    .C(_2256_),
    .Y(_2257_)
);

NAND2X1 _3141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2257_),
    .B(_2252_),
    .Y(_2258_)
);

OAI21X1 _3142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2170_),
    .B(_2195_),
    .C(_2187_),
    .Y(_2259_)
);

NOR2X1 _3143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_1639_),
    .Y(_2260_)
);

INVX1 _3144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2260_),
    .Y(_2261_)
);

NAND2X1 _3145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf0),
    .B(bregp1[6]),
    .Y(_2262_)
);

INVX2 _3146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[6]),
    .Y(_2263_)
);

OAI21X1 _3147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2263_),
    .C(_2166_),
    .Y(_2264_)
);

OAI21X1 _3148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2244_),
    .B(_2262_),
    .C(_2264_),
    .Y(_2265_)
);

XNOR2X1 _3149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2265_),
    .B(_2261_),
    .Y(_2266_)
);

OAI21X1 _3150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2175_),
    .B(_2172_),
    .C(_2173_),
    .Y(_2267_)
);

NAND2X1 _3151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[7]),
    .Y(_2268_)
);

NAND3X1 _3152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[8]),
    .C(\preg[7] [16]),
    .Y(_2269_)
);

INVX1 _3153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .Y(_2270_)
);

AOI21X1 _3154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .B(bregp1[8]),
    .C(\preg[7] [16]),
    .Y(_2271_)
);

NOR3X1 _3155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2268_),
    .B(_2271_),
    .C(_2270_),
    .Y(_2272_)
);

INVX1 _3156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2268_),
    .Y(_2273_)
);

INVX1 _3157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .Y(_2274_)
);

AOI21X1 _3158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2269_),
    .B(_2274_),
    .C(_2273_),
    .Y(_2275_)
);

OAI21X1 _3159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2272_),
    .B(_2275_),
    .C(_2267_),
    .Y(_2276_)
);

INVX1 _3160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2267_),
    .Y(_2277_)
);

NAND3X1 _3161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2273_),
    .B(_2269_),
    .C(_2274_),
    .Y(_2278_)
);

OAI21X1 _3162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2270_),
    .B(_2271_),
    .C(_2268_),
    .Y(_2279_)
);

NAND3X1 _3163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .B(_2279_),
    .C(_2277_),
    .Y(_2280_)
);

AOI21X1 _3164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2276_),
    .B(_2280_),
    .C(_2266_),
    .Y(_2281_)
);

XNOR2X1 _3165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2265_),
    .B(_2260_),
    .Y(_2282_)
);

NAND3X1 _3166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2267_),
    .B(_2278_),
    .C(_2279_),
    .Y(_2283_)
);

OAI21X1 _3167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2272_),
    .B(_2275_),
    .C(_2277_),
    .Y(_2284_)
);

AOI21X1 _3168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2283_),
    .B(_2284_),
    .C(_2282_),
    .Y(_2285_)
);

OAI21X1 _3169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2281_),
    .B(_2285_),
    .C(_2259_),
    .Y(_2286_)
);

AOI21X1 _3170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2188_),
    .B(_2186_),
    .C(_2194_),
    .Y(_2287_)
);

NAND3X1 _3171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2283_),
    .B(_2284_),
    .C(_2282_),
    .Y(_2288_)
);

INVX1 _3172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2283_),
    .Y(_2289_)
);

AOI21X1 _3173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2278_),
    .B(_2279_),
    .C(_2267_),
    .Y(_2290_)
);

OAI21X1 _3174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2289_),
    .B(_2290_),
    .C(_2266_),
    .Y(_2291_)
);

NAND3X1 _3175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2287_),
    .B(_2288_),
    .C(_2291_),
    .Y(_2292_)
);

AOI21X1 _3176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2286_),
    .B(_2292_),
    .C(_2258_),
    .Y(_2293_)
);

NAND3X1 _3177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2254_),
    .B(_2248_),
    .C(_2251_),
    .Y(_2294_)
);

NAND3X1 _3178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2235_),
    .B(_2255_),
    .C(_2256_),
    .Y(_2295_)
);

NAND2X1 _3179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2294_),
    .B(_2295_),
    .Y(_2296_)
);

NAND3X1 _3180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2259_),
    .B(_2288_),
    .C(_2291_),
    .Y(_2297_)
);

OAI21X1 _3181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2281_),
    .B(_2285_),
    .C(_2287_),
    .Y(_2298_)
);

AOI21X1 _3182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2298_),
    .B(_2297_),
    .C(_2296_),
    .Y(_2299_)
);

OAI21X1 _3183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2299_),
    .C(_2233_),
    .Y(_2300_)
);

AOI21X1 _3184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2203_),
    .B(_2201_),
    .C(_2209_),
    .Y(_2301_)
);

NAND3X1 _3185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2297_),
    .B(_2298_),
    .C(_2296_),
    .Y(_2302_)
);

NOR3X1 _3186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2281_),
    .B(_2285_),
    .C(_2287_),
    .Y(_2303_)
);

AOI21X1 _3187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2288_),
    .B(_2291_),
    .C(_2259_),
    .Y(_2304_)
);

OAI21X1 _3188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2303_),
    .B(_2304_),
    .C(_2258_),
    .Y(_2305_)
);

NAND3X1 _3189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2305_),
    .C(_2301_),
    .Y(_2306_)
);

AOI21X1 _3190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2300_),
    .B(_2306_),
    .C(_2232_),
    .Y(_2307_)
);

NAND3X1 _3191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2305_),
    .C(_2233_),
    .Y(_2308_)
);

OAI21X1 _3192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2299_),
    .C(_2301_),
    .Y(_2309_)
);

AOI21X1 _3193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2309_),
    .B(_2308_),
    .C(_2231_),
    .Y(_2310_)
);

OAI21X1 _3194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2310_),
    .C(_2230_),
    .Y(_2311_)
);

AOI21X1 _3195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2073_),
    .B(_2215_),
    .C(_2220_),
    .Y(_2312_)
);

NAND3X1 _3196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2309_),
    .C(_2308_),
    .Y(_2313_)
);

NAND3X1 _3197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2232_),
    .B(_2300_),
    .C(_2306_),
    .Y(_2314_)
);

NAND3X1 _3198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2313_),
    .B(_2314_),
    .C(_2312_),
    .Y(_2315_)
);

NAND2X1 _3199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2315_),
    .B(_2311_),
    .Y(_2316_)
);

XNOR2X1 _3200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2316_),
    .Y(\partials[15] [16])
);

AND2X2 _3201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2223_),
    .B(_2217_),
    .Y(_2317_)
);

AND2X2 _3202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2226_),
    .B(_2125_),
    .Y(_2318_)
);

OAI22X1 _3203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2227_),
    .B(_2318_),
    .C(_2317_),
    .D(_2129_),
    .Y(_2319_)
);

NOR3X1 _3204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2307_),
    .B(_2310_),
    .C(_2312_),
    .Y(_2320_)
);

AOI21X1 _3205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2316_),
    .B(_2319_),
    .C(_2320_),
    .Y(_2321_)
);

AOI21X1 _3206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2302_),
    .B(_2305_),
    .C(_2233_),
    .Y(_2322_)
);

OAI21X1 _3207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2322_),
    .B(_2232_),
    .C(_2308_),
    .Y(_2323_)
);

NAND2X1 _3208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2248_),
    .B(_2252_),
    .Y(_2324_)
);

INVX2 _3209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .Y(_2325_)
);

OAI21X1 _3210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2258_),
    .B(_2304_),
    .C(_2297_),
    .Y(_2326_)
);

OAI21X1 _3211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2234_),
    .B(_2241_),
    .C(_2240_),
    .Y(_2327_)
);

NOR2X1 _3212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2146_),
    .Y(_2328_)
);

NAND2X1 _3213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[4]),
    .B(aregp1_13_bF$buf2),
    .Y(_2329_)
);

OR2X2 _3214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2241_),
    .B(_2329_),
    .Y(_2330_)
);

OAI21X1 _3215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_2142_),
    .C(_2241_),
    .Y(_2331_)
);

NAND3X1 _3216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2328_),
    .B(_2331_),
    .C(_2330_),
    .Y(_2332_)
);

NAND2X1 _3217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[4]),
    .B(aregp1[14]),
    .Y(_2333_)
);

OAI21X1 _3218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2237_),
    .B(_2333_),
    .C(_2331_),
    .Y(_2334_)
);

OAI21X1 _3219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2077_),
    .B(_2146_),
    .C(_2334_),
    .Y(_2335_)
);

NAND2X1 _3220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf0),
    .B(bregp1[6]),
    .Y(_2336_)
);

NOR2X1 _3221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2166_),
    .B(_2336_),
    .Y(_2337_)
);

AOI21X1 _3222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2260_),
    .B(_2264_),
    .C(_2337_),
    .Y(_2338_)
);

INVX1 _3223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2338_),
    .Y(_2339_)
);

NAND3X1 _3224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .B(_2335_),
    .C(_2339_),
    .Y(_2340_)
);

INVX1 _3225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2328_),
    .Y(_2341_)
);

NOR2X1 _3226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2341_),
    .B(_2334_),
    .Y(_2342_)
);

AOI21X1 _3227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2331_),
    .B(_2330_),
    .C(_2328_),
    .Y(_2343_)
);

OAI21X1 _3228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2342_),
    .B(_2343_),
    .C(_2338_),
    .Y(_2344_)
);

NAND3X1 _3229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2340_),
    .C(_2344_),
    .Y(_2345_)
);

INVX1 _3230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .Y(_2346_)
);

NAND3X1 _3231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2332_),
    .B(_2338_),
    .C(_2335_),
    .Y(_2347_)
);

OAI21X1 _3232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2342_),
    .B(_2343_),
    .C(_2339_),
    .Y(_2348_)
);

NAND3X1 _3233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .B(_2347_),
    .C(_2348_),
    .Y(_2349_)
);

NAND2X1 _3234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2345_),
    .B(_2349_),
    .Y(_2350_)
);

OAI21X1 _3235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2266_),
    .B(_2290_),
    .C(_2283_),
    .Y(_2351_)
);

NOR2X1 _3236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1639_),
    .B(_2167_),
    .Y(_2352_)
);

INVX1 _3237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .Y(_2353_)
);

NAND2X1 _3238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf3),
    .B(bregp1[7]),
    .Y(_2354_)
);

INVX4 _3239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[7]),
    .Y(_2355_)
);

OAI21X1 _3240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2355_),
    .C(_2262_),
    .Y(_2356_)
);

OAI21X1 _3241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2336_),
    .B(_2354_),
    .C(_2356_),
    .Y(_2357_)
);

XNOR2X1 _3242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2353_),
    .Y(_2358_)
);

OAI21X1 _3243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2271_),
    .B(_2268_),
    .C(_2269_),
    .Y(_2359_)
);

NAND2X1 _3244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[8]),
    .Y(_2360_)
);

NAND3X1 _3245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[9]),
    .C(\preg[7] [17]),
    .Y(_2361_)
);

INVX1 _3246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2361_),
    .Y(_2362_)
);

AOI21X1 _3247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[9]),
    .C(\preg[7] [17]),
    .Y(_2363_)
);

NOR3X1 _3248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .B(_2363_),
    .C(_2362_),
    .Y(_2364_)
);

INVX1 _3249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2360_),
    .Y(_2365_)
);

INVX1 _3250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .Y(_2366_)
);

AOI21X1 _3251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2361_),
    .B(_2366_),
    .C(_2365_),
    .Y(_2367_)
);

OAI21X1 _3252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2367_),
    .C(_2359_),
    .Y(_2368_)
);

INVX2 _3253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .Y(_2369_)
);

NAND3X1 _3254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2365_),
    .B(_2361_),
    .C(_2366_),
    .Y(_2370_)
);

OAI21X1 _3255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2362_),
    .B(_2363_),
    .C(_2360_),
    .Y(_2371_)
);

NAND3X1 _3256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2370_),
    .B(_2371_),
    .C(_2369_),
    .Y(_2372_)
);

AOI21X1 _3257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2368_),
    .B(_2372_),
    .C(_2358_),
    .Y(_2373_)
);

XNOR2X1 _3258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2357_),
    .B(_2352_),
    .Y(_2374_)
);

NAND3X1 _3259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2359_),
    .B(_2370_),
    .C(_2371_),
    .Y(_2375_)
);

OAI21X1 _3260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2364_),
    .B(_2367_),
    .C(_2369_),
    .Y(_2376_)
);

AOI21X1 _3261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2375_),
    .B(_2376_),
    .C(_2374_),
    .Y(_2377_)
);

OAI21X1 _3262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2377_),
    .C(_2351_),
    .Y(_2378_)
);

AOI21X1 _3263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2284_),
    .B(_2282_),
    .C(_2289_),
    .Y(_2379_)
);

NAND3X1 _3264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2375_),
    .B(_2376_),
    .C(_2374_),
    .Y(_2380_)
);

NOR3X1 _3265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2367_),
    .B(_2369_),
    .C(_2364_),
    .Y(_2381_)
);

AOI21X1 _3266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2370_),
    .B(_2371_),
    .C(_2359_),
    .Y(_2382_)
);

OAI21X1 _3267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2381_),
    .B(_2382_),
    .C(_2358_),
    .Y(_2383_)
);

NAND3X1 _3268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2380_),
    .B(_2383_),
    .C(_2379_),
    .Y(_2384_)
);

AOI21X1 _3269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .B(_2384_),
    .C(_2350_),
    .Y(_2385_)
);

NAND3X1 _3270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2346_),
    .B(_2340_),
    .C(_2344_),
    .Y(_2386_)
);

NAND3X1 _3271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2327_),
    .B(_2347_),
    .C(_2348_),
    .Y(_2387_)
);

NAND2X1 _3272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2386_),
    .B(_2387_),
    .Y(_2388_)
);

NAND3X1 _3273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2380_),
    .C(_2351_),
    .Y(_2389_)
);

OAI21X1 _3274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2377_),
    .C(_2379_),
    .Y(_2390_)
);

AOI21X1 _3275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2389_),
    .B(_2390_),
    .C(_2388_),
    .Y(_2391_)
);

OAI21X1 _3276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2391_),
    .C(_2326_),
    .Y(_2392_)
);

AOI21X1 _3277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2298_),
    .B(_2296_),
    .C(_2303_),
    .Y(_2393_)
);

NAND3X1 _3278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2389_),
    .B(_2390_),
    .C(_2388_),
    .Y(_2394_)
);

NAND3X1 _3279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2378_),
    .B(_2384_),
    .C(_2350_),
    .Y(_2395_)
);

NAND3X1 _3280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2394_),
    .B(_2395_),
    .C(_2393_),
    .Y(_2396_)
);

AOI21X1 _3281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2392_),
    .B(_2396_),
    .C(_2325_),
    .Y(_2397_)
);

NAND3X1 _3282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2394_),
    .B(_2395_),
    .C(_2326_),
    .Y(_2398_)
);

OAI21X1 _3283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2391_),
    .C(_2393_),
    .Y(_2399_)
);

AOI21X1 _3284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2399_),
    .B(_2398_),
    .C(_2324_),
    .Y(_2400_)
);

OAI21X1 _3285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2400_),
    .B(_2397_),
    .C(_2323_),
    .Y(_2401_)
);

NOR3X1 _3286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2293_),
    .B(_2299_),
    .C(_2301_),
    .Y(_2402_)
);

AOI21X1 _3287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2231_),
    .B(_2309_),
    .C(_2402_),
    .Y(_2403_)
);

NAND3X1 _3288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .B(_2399_),
    .C(_2398_),
    .Y(_2404_)
);

NOR3X1 _3289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2385_),
    .B(_2391_),
    .C(_2393_),
    .Y(_2405_)
);

AOI21X1 _3290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2394_),
    .B(_2395_),
    .C(_2326_),
    .Y(_2406_)
);

OAI21X1 _3291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2405_),
    .B(_2406_),
    .C(_2325_),
    .Y(_2407_)
);

NAND3X1 _3292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_2403_),
    .C(_2407_),
    .Y(_2408_)
);

NAND2X1 _3293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2401_),
    .B(_2408_),
    .Y(_2409_)
);

XNOR2X1 _3294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2321_),
    .B(_2409_),
    .Y(\partials[15] [17])
);

NAND3X1 _3295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2313_),
    .B(_2314_),
    .C(_2230_),
    .Y(_2410_)
);

NAND3X1 _3296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2323_),
    .B(_2404_),
    .C(_2407_),
    .Y(_2411_)
);

AOI21X1 _3297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2404_),
    .B(_2407_),
    .C(_2323_),
    .Y(_2412_)
);

AOI21X1 _3298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2410_),
    .B(_2411_),
    .C(_2412_),
    .Y(_2413_)
);

AOI22X1 _3299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2311_),
    .B(_2315_),
    .C(_2401_),
    .D(_2408_),
    .Y(_2414_)
);

AOI21X1 _3300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2414_),
    .B(_2319_),
    .C(_2413_),
    .Y(_2415_)
);

OAI21X1 _3301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2406_),
    .B(_2325_),
    .C(_2398_),
    .Y(_2416_)
);

NAND2X1 _3302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2340_),
    .B(_2345_),
    .Y(_2417_)
);

INVX2 _3303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2417_),
    .Y(_2418_)
);

AOI21X1 _3304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2383_),
    .B(_2380_),
    .C(_2351_),
    .Y(_2419_)
);

OAI21X1 _3305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2350_),
    .B(_2419_),
    .C(_2389_),
    .Y(_2420_)
);

OAI21X1 _3306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2334_),
    .B(_2341_),
    .C(_2330_),
    .Y(_2421_)
);

NOR2X1 _3307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_2146_),
    .Y(_2422_)
);

NAND2X1 _3308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[5]),
    .B(aregp1_13_bF$buf1),
    .Y(_2423_)
);

OR2X2 _3309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2333_),
    .B(_2423_),
    .Y(_2424_)
);

OAI21X1 _3310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2142_),
    .C(_2333_),
    .Y(_2425_)
);

NAND3X1 _3311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2422_),
    .B(_2425_),
    .C(_2424_),
    .Y(_2426_)
);

NAND2X1 _3312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[5]),
    .B(aregp1[14]),
    .Y(_2427_)
);

OAI21X1 _3313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2329_),
    .B(_2427_),
    .C(_2425_),
    .Y(_2428_)
);

OAI21X1 _3314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2163_),
    .B(_2146_),
    .C(_2428_),
    .Y(_2429_)
);

NAND2X1 _3315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf3),
    .B(bregp1[7]),
    .Y(_2430_)
);

NOR2X1 _3316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2262_),
    .B(_2430_),
    .Y(_2431_)
);

AOI21X1 _3317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2352_),
    .B(_2356_),
    .C(_2431_),
    .Y(_2432_)
);

INVX1 _3318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2432_),
    .Y(_2433_)
);

NAND3X1 _3319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2426_),
    .B(_2429_),
    .C(_2433_),
    .Y(_2434_)
);

INVX1 _3320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2422_),
    .Y(_2435_)
);

NOR2X1 _3321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2435_),
    .B(_2428_),
    .Y(_2436_)
);

AOI21X1 _3322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2425_),
    .B(_2424_),
    .C(_2422_),
    .Y(_2437_)
);

OAI21X1 _3323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2437_),
    .C(_2432_),
    .Y(_2438_)
);

NAND3X1 _3324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2421_),
    .B(_2434_),
    .C(_2438_),
    .Y(_2439_)
);

INVX1 _3325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2421_),
    .Y(_2440_)
);

NAND3X1 _3326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2426_),
    .B(_2432_),
    .C(_2429_),
    .Y(_2441_)
);

OAI21X1 _3327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2436_),
    .B(_2437_),
    .C(_2433_),
    .Y(_2442_)
);

NAND3X1 _3328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .B(_2441_),
    .C(_2442_),
    .Y(_2443_)
);

NAND2X1 _3329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2439_),
    .B(_2443_),
    .Y(_2444_)
);

OAI21X1 _3330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2358_),
    .B(_2382_),
    .C(_2375_),
    .Y(_2445_)
);

NOR2X1 _3331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1639_),
    .B(_2263_),
    .Y(_2446_)
);

INVX1 _3332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2446_),
    .Y(_2447_)
);

NAND2X1 _3333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf2),
    .B(bregp1[8]),
    .Y(_2448_)
);

INVX2 _3334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[8]),
    .Y(_2449_)
);

OAI21X1 _3335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2449_),
    .C(_2354_),
    .Y(_2450_)
);

OAI21X1 _3336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2430_),
    .B(_2448_),
    .C(_2450_),
    .Y(_2451_)
);

XNOR2X1 _3337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2447_),
    .Y(_2452_)
);

OAI21X1 _3338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2363_),
    .B(_2360_),
    .C(_2361_),
    .Y(_2453_)
);

NAND2X1 _3339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[9]),
    .Y(_2454_)
);

NAND3X1 _3340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[10]),
    .C(\preg[7] [18]),
    .Y(_2455_)
);

INVX1 _3341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .Y(_2456_)
);

AOI21X1 _3342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[10]),
    .C(\preg[7] [18]),
    .Y(_2457_)
);

NOR3X1 _3343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2454_),
    .B(_2457_),
    .C(_2456_),
    .Y(_2458_)
);

INVX1 _3344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2454_),
    .Y(_2459_)
);

INVX1 _3345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .Y(_2460_)
);

AOI21X1 _3346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2455_),
    .B(_2460_),
    .C(_2459_),
    .Y(_2461_)
);

OAI21X1 _3347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2458_),
    .B(_2461_),
    .C(_2453_),
    .Y(_2462_)
);

INVX2 _3348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2453_),
    .Y(_2463_)
);

NAND3X1 _3349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2459_),
    .B(_2455_),
    .C(_2460_),
    .Y(_2464_)
);

OAI21X1 _3350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2456_),
    .B(_2457_),
    .C(_2454_),
    .Y(_2465_)
);

NAND3X1 _3351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2464_),
    .B(_2465_),
    .C(_2463_),
    .Y(_2466_)
);

AOI21X1 _3352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2462_),
    .B(_2466_),
    .C(_2452_),
    .Y(_2467_)
);

XNOR2X1 _3353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2451_),
    .B(_2446_),
    .Y(_2468_)
);

NAND3X1 _3354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2453_),
    .B(_2464_),
    .C(_2465_),
    .Y(_2469_)
);

OAI21X1 _3355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2458_),
    .B(_2461_),
    .C(_2463_),
    .Y(_2470_)
);

AOI21X1 _3356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2470_),
    .C(_2468_),
    .Y(_2471_)
);

OAI21X1 _3357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2471_),
    .C(_2445_),
    .Y(_2472_)
);

AOI21X1 _3358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2376_),
    .B(_2374_),
    .C(_2381_),
    .Y(_2473_)
);

NAND3X1 _3359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2469_),
    .B(_2470_),
    .C(_2468_),
    .Y(_2474_)
);

NOR3X1 _3360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2461_),
    .B(_2463_),
    .C(_2458_),
    .Y(_2475_)
);

AOI21X1 _3361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2464_),
    .B(_2465_),
    .C(_2453_),
    .Y(_2476_)
);

OAI21X1 _3362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2475_),
    .B(_2476_),
    .C(_2452_),
    .Y(_2477_)
);

NAND3X1 _3363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2474_),
    .C(_2473_),
    .Y(_2478_)
);

AOI21X1 _3364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2472_),
    .B(_2478_),
    .C(_2444_),
    .Y(_2479_)
);

NAND3X1 _3365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2440_),
    .B(_2434_),
    .C(_2438_),
    .Y(_2480_)
);

NAND3X1 _3366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2421_),
    .B(_2441_),
    .C(_2442_),
    .Y(_2481_)
);

NAND2X1 _3367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2480_),
    .B(_2481_),
    .Y(_2482_)
);

NAND3X1 _3368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2474_),
    .C(_2445_),
    .Y(_2483_)
);

OAI21X1 _3369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2471_),
    .C(_2473_),
    .Y(_2484_)
);

AOI21X1 _3370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2484_),
    .C(_2482_),
    .Y(_2485_)
);

OAI21X1 _3371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2485_),
    .C(_2420_),
    .Y(_2486_)
);

NOR3X1 _3372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2373_),
    .B(_2377_),
    .C(_2379_),
    .Y(_2487_)
);

AOI21X1 _3373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2390_),
    .B(_2388_),
    .C(_2487_),
    .Y(_2488_)
);

NAND3X1 _3374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2483_),
    .B(_2484_),
    .C(_2482_),
    .Y(_2489_)
);

NOR3X1 _3375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2467_),
    .B(_2471_),
    .C(_2473_),
    .Y(_2490_)
);

AOI21X1 _3376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2477_),
    .B(_2474_),
    .C(_2445_),
    .Y(_2491_)
);

OAI21X1 _3377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2490_),
    .B(_2491_),
    .C(_2444_),
    .Y(_2492_)
);

NAND3X1 _3378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .B(_2488_),
    .C(_2492_),
    .Y(_2493_)
);

AOI21X1 _3379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2486_),
    .B(_2493_),
    .C(_2418_),
    .Y(_2494_)
);

NAND3X1 _3380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .B(_2420_),
    .C(_2492_),
    .Y(_2495_)
);

OAI21X1 _3381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2485_),
    .C(_2488_),
    .Y(_2496_)
);

AOI21X1 _3382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2496_),
    .B(_2495_),
    .C(_2417_),
    .Y(_2497_)
);

OAI21X1 _3383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2494_),
    .B(_2497_),
    .C(_2416_),
    .Y(_2498_)
);

AOI21X1 _3384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2324_),
    .B(_2399_),
    .C(_2405_),
    .Y(_2499_)
);

NAND3X1 _3385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2417_),
    .B(_2496_),
    .C(_2495_),
    .Y(_2500_)
);

NOR3X1 _3386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2479_),
    .B(_2485_),
    .C(_2488_),
    .Y(_2501_)
);

AOI21X1 _3387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2489_),
    .B(_2492_),
    .C(_2420_),
    .Y(_2502_)
);

OAI21X1 _3388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2501_),
    .B(_2502_),
    .C(_2418_),
    .Y(_2503_)
);

NAND3X1 _3389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2500_),
    .B(_2499_),
    .C(_2503_),
    .Y(_2504_)
);

NAND2X1 _3390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2498_),
    .B(_2504_),
    .Y(_2505_)
);

XNOR2X1 _3391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2505_),
    .Y(\partials[15] [18])
);

NAND3X1 _3392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2500_),
    .B(_2416_),
    .C(_2503_),
    .Y(_2506_)
);

INVX1 _3393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2505_),
    .Y(_2507_)
);

OAI21X1 _3394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2415_),
    .B(_2507_),
    .C(_2506_),
    .Y(_2508_)
);

OAI21X1 _3395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2502_),
    .B(_2418_),
    .C(_2495_),
    .Y(_2509_)
);

NAND2X1 _3396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2434_),
    .B(_2439_),
    .Y(_2510_)
);

OAI21X1 _3397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2444_),
    .B(_2491_),
    .C(_2483_),
    .Y(_2511_)
);

OAI21X1 _3398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2428_),
    .B(_2435_),
    .C(_2424_),
    .Y(_2512_)
);

INVX1 _3399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2512_),
    .Y(_2513_)
);

NOR2X1 _3400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_2146_),
    .Y(_2514_)
);

INVX1 _3401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2427_),
    .Y(_2515_)
);

NAND2X1 _3402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf0),
    .B(bregp1[6]),
    .Y(_2516_)
);

INVX1 _3403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .Y(_2517_)
);

NAND2X1 _3404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2515_),
    .B(_2517_),
    .Y(_2518_)
);

OAI21X1 _3405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2263_),
    .C(_2427_),
    .Y(_2519_)
);

NAND3X1 _3406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .B(_2519_),
    .C(_2518_),
    .Y(_2520_)
);

NAND2X1 _3407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[6]),
    .B(aregp1[14]),
    .Y(_2521_)
);

OAI21X1 _3408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2423_),
    .B(_2521_),
    .C(_2519_),
    .Y(_2522_)
);

OAI21X1 _3409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2080_),
    .B(_2146_),
    .C(_2522_),
    .Y(_2523_)
);

NAND2X1 _3410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf2),
    .B(bregp1[8]),
    .Y(_2524_)
);

NOR2X1 _3411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2354_),
    .B(_2524_),
    .Y(_2525_)
);

AOI21X1 _3412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2446_),
    .B(_2450_),
    .C(_2525_),
    .Y(_2526_)
);

INVX1 _3413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2526_),
    .Y(_2527_)
);

NAND3X1 _3414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2520_),
    .B(_2523_),
    .C(_2527_),
    .Y(_2528_)
);

INVX1 _3415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2514_),
    .Y(_2529_)
);

NOR2X1 _3416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2529_),
    .B(_2522_),
    .Y(_2530_)
);

AOI21X1 _3417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2519_),
    .B(_2518_),
    .C(_2514_),
    .Y(_2531_)
);

OAI21X1 _3418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2531_),
    .C(_2526_),
    .Y(_2532_)
);

NAND3X1 _3419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2528_),
    .C(_2532_),
    .Y(_2533_)
);

NAND3X1 _3420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2526_),
    .B(_2520_),
    .C(_2523_),
    .Y(_2534_)
);

OAI21X1 _3421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2530_),
    .B(_2531_),
    .C(_2527_),
    .Y(_2535_)
);

NAND3X1 _3422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2512_),
    .B(_2534_),
    .C(_2535_),
    .Y(_2536_)
);

NAND2X1 _3423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2533_),
    .B(_2536_),
    .Y(_2537_)
);

OAI21X1 _3424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2452_),
    .B(_2476_),
    .C(_2469_),
    .Y(_2538_)
);

NOR2X1 _3425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1639_),
    .B(_2355_),
    .Y(_2539_)
);

NAND2X1 _3426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf1),
    .B(bregp1[9]),
    .Y(_2540_)
);

INVX1 _3427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[9]),
    .Y(_2541_)
);

OAI21X1 _3428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2541_),
    .C(_2448_),
    .Y(_2542_)
);

OAI21X1 _3429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2524_),
    .B(_2540_),
    .C(_2542_),
    .Y(_2543_)
);

XNOR2X1 _3430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_2539_),
    .Y(_2544_)
);

OAI21X1 _3431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2457_),
    .B(_2454_),
    .C(_2455_),
    .Y(_2545_)
);

NAND2X1 _3432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[10]),
    .Y(_2546_)
);

INVX1 _3433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .Y(_2547_)
);

NAND3X1 _3434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .B(bregp1[11]),
    .C(\preg[7] [19]),
    .Y(_2548_)
);

AOI21X1 _3435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[11]),
    .C(\preg[7] [19]),
    .Y(_2549_)
);

INVX1 _3436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2549_),
    .Y(_2550_)
);

NAND3X1 _3437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2547_),
    .B(_2548_),
    .C(_2550_),
    .Y(_2551_)
);

INVX1 _3438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2548_),
    .Y(_2552_)
);

OAI21X1 _3439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2552_),
    .B(_2549_),
    .C(_2546_),
    .Y(_2553_)
);

NAND3X1 _3440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .B(_2551_),
    .C(_2553_),
    .Y(_2554_)
);

INVX2 _3441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2545_),
    .Y(_2555_)
);

NOR3X1 _3442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2546_),
    .B(_2549_),
    .C(_2552_),
    .Y(_2556_)
);

AOI21X1 _3443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2548_),
    .B(_2550_),
    .C(_2547_),
    .Y(_2557_)
);

OAI21X1 _3444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2556_),
    .B(_2557_),
    .C(_2555_),
    .Y(_2558_)
);

NAND3X1 _3445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2558_),
    .C(_2544_),
    .Y(_2559_)
);

INVX1 _3446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2539_),
    .Y(_2560_)
);

XNOR2X1 _3447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2543_),
    .B(_2560_),
    .Y(_2561_)
);

NOR3X1 _3448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2557_),
    .B(_2555_),
    .C(_2556_),
    .Y(_2562_)
);

AOI21X1 _3449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_2553_),
    .C(_2545_),
    .Y(_2563_)
);

OAI21X1 _3450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2562_),
    .B(_2563_),
    .C(_2561_),
    .Y(_2564_)
);

NAND3X1 _3451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2559_),
    .C(_2538_),
    .Y(_2565_)
);

AOI21X1 _3452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2470_),
    .B(_2468_),
    .C(_2475_),
    .Y(_2566_)
);

OAI21X1 _3453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2556_),
    .B(_2557_),
    .C(_2545_),
    .Y(_2567_)
);

NAND3X1 _3454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2551_),
    .B(_2553_),
    .C(_2555_),
    .Y(_2568_)
);

AOI21X1 _3455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2567_),
    .B(_2568_),
    .C(_2561_),
    .Y(_2569_)
);

AOI21X1 _3456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2554_),
    .B(_2558_),
    .C(_2544_),
    .Y(_2570_)
);

OAI21X1 _3457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2569_),
    .B(_2570_),
    .C(_2566_),
    .Y(_2571_)
);

NAND3X1 _3458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2565_),
    .B(_2571_),
    .C(_2537_),
    .Y(_2572_)
);

NAND3X1 _3459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2512_),
    .B(_2528_),
    .C(_2532_),
    .Y(_2573_)
);

NAND3X1 _3460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2513_),
    .B(_2534_),
    .C(_2535_),
    .Y(_2574_)
);

NAND2X1 _3461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2573_),
    .B(_2574_),
    .Y(_2575_)
);

NOR3X1 _3462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2569_),
    .B(_2570_),
    .C(_2566_),
    .Y(_2576_)
);

AOI21X1 _3463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2559_),
    .C(_2538_),
    .Y(_2577_)
);

OAI21X1 _3464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2576_),
    .B(_2577_),
    .C(_2575_),
    .Y(_2578_)
);

NAND3X1 _3465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2572_),
    .B(_2511_),
    .C(_2578_),
    .Y(_2579_)
);

AOI21X1 _3466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2484_),
    .B(_2482_),
    .C(_2490_),
    .Y(_2580_)
);

OAI21X1 _3467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2569_),
    .B(_2570_),
    .C(_2538_),
    .Y(_2581_)
);

NAND3X1 _3468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2564_),
    .B(_2559_),
    .C(_2566_),
    .Y(_2582_)
);

AOI21X1 _3469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2581_),
    .B(_2582_),
    .C(_2575_),
    .Y(_2583_)
);

AOI21X1 _3470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2565_),
    .B(_2571_),
    .C(_2537_),
    .Y(_2584_)
);

OAI21X1 _3471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2580_),
    .Y(_2585_)
);

NAND3X1 _3472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2585_),
    .C(_2579_),
    .Y(_2586_)
);

INVX2 _3473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .Y(_2587_)
);

NOR3X1 _3474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2580_),
    .Y(_2588_)
);

AOI21X1 _3475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2572_),
    .B(_2578_),
    .C(_2511_),
    .Y(_2589_)
);

OAI21X1 _3476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2588_),
    .B(_2589_),
    .C(_2587_),
    .Y(_2590_)
);

NAND3X1 _3477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2509_),
    .C(_2590_),
    .Y(_2591_)
);

AOI21X1 _3478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2417_),
    .B(_2496_),
    .C(_2501_),
    .Y(_2592_)
);

OAI21X1 _3479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2583_),
    .B(_2584_),
    .C(_2511_),
    .Y(_2593_)
);

NAND3X1 _3480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2572_),
    .B(_2580_),
    .C(_2578_),
    .Y(_2594_)
);

AOI21X1 _3481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2593_),
    .B(_2594_),
    .C(_2587_),
    .Y(_2595_)
);

AOI21X1 _3482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2585_),
    .B(_2579_),
    .C(_2510_),
    .Y(_2596_)
);

OAI21X1 _3483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .B(_2596_),
    .C(_2592_),
    .Y(_2597_)
);

NAND2X1 _3484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2591_),
    .Y(_2598_)
);

XNOR2X1 _3485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2508_),
    .B(_2598_),
    .Y(\partials[15] [19])
);

OAI21X1 _3486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .B(_2596_),
    .C(_2509_),
    .Y(_2599_)
);

NAND3X1 _3487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2592_),
    .B(_2586_),
    .C(_2590_),
    .Y(_2600_)
);

AOI22X1 _3488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2600_),
    .B(_2599_),
    .C(_2498_),
    .D(_2504_),
    .Y(_2601_)
);

NAND2X1 _3489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2591_),
    .B(_2506_),
    .Y(_2602_)
);

AOI22X1 _3490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2602_),
    .C(_2413_),
    .D(_2601_),
    .Y(_2603_)
);

NAND2X1 _3491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2601_),
    .B(_2414_),
    .Y(_2604_)
);

OAI21X1 _3492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2229_),
    .B(_2604_),
    .C(_2603_),
    .Y(_2605_)
);

AOI21X1 _3493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2510_),
    .B(_2585_),
    .C(_2588_),
    .Y(_2606_)
);

NAND2X1 _3494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2528_),
    .B(_2573_),
    .Y(_2607_)
);

INVX2 _3495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .Y(_2608_)
);

OAI21X1 _3496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2575_),
    .B(_2577_),
    .C(_2565_),
    .Y(_2609_)
);

OAI21X1 _3497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2522_),
    .B(_2529_),
    .C(_2518_),
    .Y(_2610_)
);

NOR2X1 _3498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2146_),
    .Y(_2611_)
);

AND2X2 _3499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[7]),
    .Y(_2612_)
);

NAND2X1 _3500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2612_),
    .B(_2517_),
    .Y(_2613_)
);

OAI21X1 _3501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2355_),
    .C(_2521_),
    .Y(_2614_)
);

NAND3X1 _3502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .B(_2614_),
    .C(_2613_),
    .Y(_2615_)
);

NAND2X1 _3503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[7]),
    .Y(_2616_)
);

OAI21X1 _3504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2516_),
    .B(_2616_),
    .C(_2614_),
    .Y(_2617_)
);

OAI21X1 _3505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2167_),
    .B(_2146_),
    .C(_2617_),
    .Y(_2618_)
);

NAND2X1 _3506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf1),
    .B(bregp1[9]),
    .Y(_2619_)
);

NOR2X1 _3507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2448_),
    .B(_2619_),
    .Y(_2620_)
);

AOI21X1 _3508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2539_),
    .B(_2542_),
    .C(_2620_),
    .Y(_2621_)
);

INVX1 _3509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .Y(_2622_)
);

NAND3X1 _3510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2615_),
    .B(_2618_),
    .C(_2622_),
    .Y(_2623_)
);

INVX1 _3511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2611_),
    .Y(_2624_)
);

NOR2X1 _3512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2624_),
    .B(_2617_),
    .Y(_2625_)
);

AOI21X1 _3513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2614_),
    .B(_2613_),
    .C(_2611_),
    .Y(_2626_)
);

OAI21X1 _3514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2625_),
    .B(_2626_),
    .C(_2621_),
    .Y(_2627_)
);

NAND3X1 _3515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2623_),
    .C(_2627_),
    .Y(_2628_)
);

INVX1 _3516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .Y(_2629_)
);

NAND3X1 _3517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2621_),
    .B(_2615_),
    .C(_2618_),
    .Y(_2630_)
);

OAI21X1 _3518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2625_),
    .B(_2626_),
    .C(_2622_),
    .Y(_2631_)
);

NAND3X1 _3519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2629_),
    .B(_2630_),
    .C(_2631_),
    .Y(_2632_)
);

NAND2X1 _3520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2628_),
    .B(_2632_),
    .Y(_2633_)
);

OAI21X1 _3521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2561_),
    .B(_2563_),
    .C(_2554_),
    .Y(_2634_)
);

NAND2X1 _3522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[8]),
    .Y(_2635_)
);

NAND2X1 _3523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf0),
    .B(bregp1[10]),
    .Y(_2636_)
);

INVX1 _3524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[10]),
    .Y(_2637_)
);

OAI21X1 _3525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_2637_),
    .C(_2540_),
    .Y(_2638_)
);

OAI21X1 _3526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2636_),
    .C(_2638_),
    .Y(_2639_)
);

XNOR2X1 _3527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2635_),
    .Y(_2640_)
);

OAI21X1 _3528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2549_),
    .B(_2546_),
    .C(_2548_),
    .Y(_2641_)
);

NAND2X1 _3529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[11]),
    .Y(_2642_)
);

NAND3X1 _3530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[12]),
    .C(\preg[7] [20]),
    .Y(_2643_)
);

INVX1 _3531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2643_),
    .Y(_2644_)
);

AOI21X1 _3532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[12]),
    .C(\preg[7] [20]),
    .Y(_2645_)
);

NOR3X1 _3533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2642_),
    .B(_2645_),
    .C(_2644_),
    .Y(_2646_)
);

INVX1 _3534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2642_),
    .Y(_2647_)
);

INVX1 _3535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2645_),
    .Y(_2648_)
);

AOI21X1 _3536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2643_),
    .B(_2648_),
    .C(_2647_),
    .Y(_2649_)
);

OAI21X1 _3537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2646_),
    .B(_2649_),
    .C(_2641_),
    .Y(_2650_)
);

INVX2 _3538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2641_),
    .Y(_2651_)
);

NAND3X1 _3539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2647_),
    .B(_2643_),
    .C(_2648_),
    .Y(_2652_)
);

OAI21X1 _3540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2644_),
    .B(_2645_),
    .C(_2642_),
    .Y(_2653_)
);

NAND3X1 _3541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2653_),
    .C(_2651_),
    .Y(_2654_)
);

AOI21X1 _3542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2650_),
    .B(_2654_),
    .C(_2640_),
    .Y(_2655_)
);

INVX2 _3543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2635_),
    .Y(_2656_)
);

XNOR2X1 _3544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2639_),
    .B(_2656_),
    .Y(_2657_)
);

NAND3X1 _3545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2641_),
    .B(_2652_),
    .C(_2653_),
    .Y(_2658_)
);

OAI21X1 _3546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2646_),
    .B(_2649_),
    .C(_2651_),
    .Y(_2659_)
);

AOI21X1 _3547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2659_),
    .C(_2657_),
    .Y(_2660_)
);

OAI21X1 _3548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2660_),
    .C(_2634_),
    .Y(_2661_)
);

AOI21X1 _3549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2558_),
    .B(_2544_),
    .C(_2562_),
    .Y(_2662_)
);

NAND3X1 _3550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2658_),
    .B(_2659_),
    .C(_2657_),
    .Y(_2663_)
);

NOR3X1 _3551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2649_),
    .B(_2651_),
    .C(_2646_),
    .Y(_2664_)
);

AOI21X1 _3552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2652_),
    .B(_2653_),
    .C(_2641_),
    .Y(_2665_)
);

OAI21X1 _3553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2664_),
    .B(_2665_),
    .C(_2640_),
    .Y(_2666_)
);

NAND3X1 _3554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .B(_2663_),
    .C(_2662_),
    .Y(_2667_)
);

AOI21X1 _3555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2667_),
    .C(_2633_),
    .Y(_2668_)
);

NAND3X1 _3556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2629_),
    .B(_2623_),
    .C(_2627_),
    .Y(_2669_)
);

NAND3X1 _3557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2610_),
    .B(_2630_),
    .C(_2631_),
    .Y(_2670_)
);

NAND2X1 _3558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2669_),
    .B(_2670_),
    .Y(_2671_)
);

NAND3X1 _3559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .B(_2663_),
    .C(_2634_),
    .Y(_2672_)
);

OAI21X1 _3560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2660_),
    .C(_2662_),
    .Y(_2673_)
);

AOI21X1 _3561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .B(_2673_),
    .C(_2671_),
    .Y(_2674_)
);

OAI21X1 _3562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2668_),
    .B(_2674_),
    .C(_2609_),
    .Y(_2675_)
);

AOI21X1 _3563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2571_),
    .B(_2537_),
    .C(_2576_),
    .Y(_2676_)
);

NAND3X1 _3564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2672_),
    .B(_2673_),
    .C(_2671_),
    .Y(_2677_)
);

NAND3X1 _3565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2661_),
    .B(_2667_),
    .C(_2633_),
    .Y(_2678_)
);

NAND3X1 _3566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2678_),
    .C(_2676_),
    .Y(_2679_)
);

AOI21X1 _3567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2679_),
    .B(_2675_),
    .C(_2608_),
    .Y(_2680_)
);

NAND3X1 _3568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2678_),
    .C(_2609_),
    .Y(_2681_)
);

OAI21X1 _3569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2668_),
    .B(_2674_),
    .C(_2676_),
    .Y(_2682_)
);

AOI21X1 _3570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2681_),
    .B(_2682_),
    .C(_2607_),
    .Y(_2683_)
);

OAI21X1 _3571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .B(_2683_),
    .C(_2606_),
    .Y(_2684_)
);

OAI21X1 _3572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2589_),
    .B(_2587_),
    .C(_2579_),
    .Y(_2685_)
);

NAND3X1 _3573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2681_),
    .C(_2682_),
    .Y(_2686_)
);

NAND3X1 _3574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2608_),
    .B(_2679_),
    .C(_2675_),
    .Y(_2687_)
);

NAND3X1 _3575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2686_),
    .B(_2687_),
    .C(_2685_),
    .Y(_2688_)
);

NAND2X1 _3576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2688_),
    .Y(_2689_)
);

XNOR2X1 _3577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2605_),
    .B(_2689_),
    .Y(\partials[15] [20])
);

NOR3X1 _3578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2680_),
    .B(_2683_),
    .C(_2606_),
    .Y(_2690_)
);

AOI21X1 _3579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2684_),
    .B(_2605_),
    .C(_2690_),
    .Y(_2691_)
);

NOR3X1 _3580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2668_),
    .B(_2674_),
    .C(_2676_),
    .Y(_2692_)
);

AOI21X1 _3581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2607_),
    .B(_2682_),
    .C(_2692_),
    .Y(_2693_)
);

NAND2X1 _3582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2623_),
    .B(_2628_),
    .Y(_2694_)
);

INVX2 _3583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .Y(_2695_)
);

AOI21X1 _3584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2666_),
    .B(_2663_),
    .C(_2634_),
    .Y(_2696_)
);

OAI21X1 _3585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2633_),
    .B(_2696_),
    .C(_2672_),
    .Y(_2697_)
);

OAI21X1 _3586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2617_),
    .B(_2624_),
    .C(_2613_),
    .Y(_2698_)
);

NOR2X1 _3587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2263_),
    .B(_2146_),
    .Y(_2699_)
);

AND2X2 _3588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf3),
    .B(bregp1[8]),
    .Y(_2700_)
);

NAND2X1 _3589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2612_),
    .B(_2700_),
    .Y(_2701_)
);

NAND2X1 _3590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf2),
    .B(bregp1[8]),
    .Y(_2702_)
);

OAI21X1 _3591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2355_),
    .C(_2702_),
    .Y(_2703_)
);

NAND3X1 _3592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2699_),
    .B(_2703_),
    .C(_2701_),
    .Y(_2704_)
);

INVX1 _3593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2699_),
    .Y(_2705_)
);

OAI21X1 _3594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2355_),
    .C(_2700_),
    .Y(_2706_)
);

OAI21X1 _3595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_2449_),
    .C(_2612_),
    .Y(_2707_)
);

NAND3X1 _3596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .B(_2707_),
    .C(_2705_),
    .Y(_2708_)
);

NAND2X1 _3597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf0),
    .B(bregp1[10]),
    .Y(_2709_)
);

NOR2X1 _3598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_2709_),
    .Y(_2710_)
);

AOI21X1 _3599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2656_),
    .B(_2638_),
    .C(_2710_),
    .Y(_2711_)
);

NAND3X1 _3600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2711_),
    .B(_2704_),
    .C(_2708_),
    .Y(_2712_)
);

AOI21X1 _3601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2706_),
    .B(_2707_),
    .C(_2705_),
    .Y(_2713_)
);

AOI21X1 _3602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2703_),
    .B(_2701_),
    .C(_2699_),
    .Y(_2714_)
);

AND2X2 _3603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2540_),
    .B(_2709_),
    .Y(_2715_)
);

OAI22X1 _3604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2619_),
    .B(_2636_),
    .C(_2715_),
    .D(_2635_),
    .Y(_2716_)
);

OAI21X1 _3605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2713_),
    .B(_2714_),
    .C(_2716_),
    .Y(_2717_)
);

AOI21X1 _3606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2717_),
    .C(_2698_),
    .Y(_2718_)
);

INVX1 _3607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2698_),
    .Y(_2719_)
);

NAND3X1 _3608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2704_),
    .B(_2716_),
    .C(_2708_),
    .Y(_2720_)
);

OAI21X1 _3609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2713_),
    .B(_2714_),
    .C(_2711_),
    .Y(_2721_)
);

AOI21X1 _3610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .B(_2721_),
    .C(_2719_),
    .Y(_2722_)
);

NOR2X1 _3611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2718_),
    .B(_2722_),
    .Y(_2723_)
);

OAI21X1 _3612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2640_),
    .B(_2665_),
    .C(_2658_),
    .Y(_2724_)
);

NAND2X1 _3613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[9]),
    .Y(_2725_)
);

INVX1 _3614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2725_),
    .Y(_2726_)
);

NAND2X1 _3615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf3),
    .B(bregp1[11]),
    .Y(_2727_)
);

OR2X2 _3616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2727_),
    .Y(_2728_)
);

OAI21X1 _3617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_2637_),
    .C(_2727_),
    .Y(_2729_)
);

NAND3X1 _3618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2726_),
    .B(_2729_),
    .C(_2728_),
    .Y(_2730_)
);

NOR2X1 _3619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2727_),
    .Y(_2731_)
);

AND2X2 _3620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2636_),
    .B(_2727_),
    .Y(_2732_)
);

OAI21X1 _3621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2732_),
    .B(_2731_),
    .C(_2725_),
    .Y(_2733_)
);

NAND2X1 _3622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2733_),
    .B(_2730_),
    .Y(_2734_)
);

OAI21X1 _3623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2645_),
    .B(_2642_),
    .C(_2643_),
    .Y(_2735_)
);

NAND2X1 _3624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[12]),
    .Y(_2736_)
);

NAND3X1 _3625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[13]),
    .C(\preg[7] [21]),
    .Y(_2737_)
);

INVX1 _3626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .Y(_2738_)
);

AOI21X1 _3627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf4),
    .B(bregp1[13]),
    .C(\preg[7] [21]),
    .Y(_2739_)
);

NOR3X1 _3628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .B(_2739_),
    .C(_2738_),
    .Y(_2740_)
);

INVX1 _3629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2736_),
    .Y(_2741_)
);

INVX1 _3630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .Y(_2742_)
);

AOI21X1 _3631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2737_),
    .B(_2742_),
    .C(_2741_),
    .Y(_2743_)
);

OAI21X1 _3632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2740_),
    .B(_2743_),
    .C(_2735_),
    .Y(_0_)
);

INVX2 _3633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2735_),
    .Y(_1_)
);

NAND3X1 _3634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2741_),
    .B(_2737_),
    .C(_2742_),
    .Y(_2_)
);

OAI21X1 _3635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2738_),
    .B(_2739_),
    .C(_2736_),
    .Y(_3_)
);

NAND3X1 _3636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_3_),
    .C(_1_),
    .Y(_4_)
);

AOI21X1 _3637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_4_),
    .B(_0_),
    .C(_2734_),
    .Y(_5_)
);

AND2X2 _3638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2730_),
    .B(_2733_),
    .Y(_6_)
);

NAND3X1 _3639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2735_),
    .B(_2_),
    .C(_3_),
    .Y(_7_)
);

OAI21X1 _3640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2740_),
    .B(_2743_),
    .C(_1_),
    .Y(_8_)
);

AOI21X1 _3641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_8_),
    .C(_6_),
    .Y(_9_)
);

OAI21X1 _3642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_5_),
    .C(_2724_),
    .Y(_10_)
);

AOI21X1 _3643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2659_),
    .B(_2657_),
    .C(_2664_),
    .Y(_11_)
);

NAND3X1 _3644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_7_),
    .B(_8_),
    .C(_6_),
    .Y(_12_)
);

NOR3X1 _3645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2743_),
    .B(_1_),
    .C(_2740_),
    .Y(_13_)
);

AOI21X1 _3646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2_),
    .B(_3_),
    .C(_2735_),
    .Y(_14_)
);

OAI21X1 _3647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_13_),
    .B(_14_),
    .C(_2734_),
    .Y(_15_)
);

NAND3X1 _3648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_15_),
    .C(_11_),
    .Y(_16_)
);

AOI21X1 _3649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(_16_),
    .C(_2723_),
    .Y(_17_)
);

AOI21X1 _3650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2712_),
    .B(_2717_),
    .C(_2719_),
    .Y(_18_)
);

AOI21X1 _3651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .B(_2721_),
    .C(_2698_),
    .Y(_19_)
);

NOR2X1 _3652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_19_),
    .B(_18_),
    .Y(_20_)
);

NAND3X1 _3653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_15_),
    .C(_2724_),
    .Y(_21_)
);

OAI21X1 _3654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_5_),
    .C(_11_),
    .Y(_22_)
);

AOI21X1 _3655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_22_),
    .B(_21_),
    .C(_20_),
    .Y(_23_)
);

OAI21X1 _3656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_23_),
    .C(_2697_),
    .Y(_24_)
);

NOR3X1 _3657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2655_),
    .B(_2660_),
    .C(_2662_),
    .Y(_25_)
);

AOI21X1 _3658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2673_),
    .B(_2671_),
    .C(_25_),
    .Y(_26_)
);

NAND3X1 _3659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_22_),
    .B(_21_),
    .C(_20_),
    .Y(_27_)
);

NAND3X1 _3660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_10_),
    .B(_16_),
    .C(_2723_),
    .Y(_28_)
);

NAND3X1 _3661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_28_),
    .C(_26_),
    .Y(_29_)
);

AOI21X1 _3662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_24_),
    .B(_29_),
    .C(_2695_),
    .Y(_30_)
);

NAND3X1 _3663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_28_),
    .C(_2697_),
    .Y(_31_)
);

OAI21X1 _3664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_23_),
    .C(_26_),
    .Y(_32_)
);

AOI21X1 _3665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_32_),
    .B(_31_),
    .C(_2694_),
    .Y(_33_)
);

NOR3X1 _3666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_33_),
    .C(_2693_),
    .Y(_34_)
);

AOI21X1 _3667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2677_),
    .B(_2678_),
    .C(_2609_),
    .Y(_35_)
);

OAI21X1 _3668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_35_),
    .B(_2608_),
    .C(_2681_),
    .Y(_36_)
);

NAND3X1 _3669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .B(_32_),
    .C(_31_),
    .Y(_37_)
);

NOR3X1 _3670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_17_),
    .B(_23_),
    .C(_26_),
    .Y(_38_)
);

AOI21X1 _3671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_27_),
    .B(_28_),
    .C(_2697_),
    .Y(_39_)
);

OAI21X1 _3672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_38_),
    .B(_39_),
    .C(_2695_),
    .Y(_40_)
);

AOI21X1 _3673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_37_),
    .B(_40_),
    .C(_36_),
    .Y(_41_)
);

NOR2X1 _3674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_34_),
    .Y(_42_)
);

XNOR2X1 _3675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2691_),
    .B(_42_),
    .Y(\partials[15] [21])
);

OAI21X1 _3676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_30_),
    .B(_33_),
    .C(_2693_),
    .Y(_43_)
);

AOI21X1 _3677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_2690_),
    .C(_34_),
    .Y(_44_)
);

NAND3X1 _3678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_36_),
    .B(_37_),
    .C(_40_),
    .Y(_45_)
);

NAND2X1 _3679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_43_),
    .B(_45_),
    .Y(_46_)
);

NOR2X1 _3680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_46_),
    .Y(_47_)
);

NAND2X1 _3681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_47_),
    .B(_2605_),
    .Y(_48_)
);

OAI21X1 _3682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_39_),
    .B(_2695_),
    .C(_31_),
    .Y(_49_)
);

INVX1 _3683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2720_),
    .Y(_50_)
);

NOR2X1 _3684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_50_),
    .B(_18_),
    .Y(_51_)
);

AOI21X1 _3685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_12_),
    .B(_15_),
    .C(_2724_),
    .Y(_52_)
);

OAI21X1 _3686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2723_),
    .B(_52_),
    .C(_21_),
    .Y(_53_)
);

OAI21X1 _3687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2616_),
    .B(_2702_),
    .C(_2704_),
    .Y(_54_)
);

NOR2X1 _3688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2355_),
    .B(_2146_),
    .Y(_55_)
);

NAND2X1 _3689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[9]),
    .Y(_56_)
);

INVX2 _3690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_56_),
    .Y(_57_)
);

NAND2X1 _3691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2700_),
    .B(_57_),
    .Y(_58_)
);

NAND2X1 _3692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf1),
    .B(bregp1[9]),
    .Y(_59_)
);

OAI21X1 _3693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2449_),
    .C(_59_),
    .Y(_60_)
);

NAND3X1 _3694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .B(_60_),
    .C(_58_),
    .Y(_61_)
);

INVX1 _3695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_55_),
    .Y(_62_)
);

INVX1 _3696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .Y(_63_)
);

OAI21X1 _3697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2449_),
    .C(_63_),
    .Y(_64_)
);

NAND3X1 _3698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[8]),
    .C(_59_),
    .Y(_65_)
);

NAND3X1 _3699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_65_),
    .B(_62_),
    .C(_64_),
    .Y(_66_)
);

AOI21X1 _3700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2726_),
    .B(_2729_),
    .C(_2731_),
    .Y(_67_)
);

INVX1 _3701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .Y(_68_)
);

NAND3X1 _3702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_66_),
    .C(_68_),
    .Y(_69_)
);

AOI21X1 _3703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_65_),
    .B(_64_),
    .C(_62_),
    .Y(_70_)
);

AOI21X1 _3704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_60_),
    .B(_58_),
    .C(_55_),
    .Y(_71_)
);

OAI21X1 _3705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_71_),
    .C(_67_),
    .Y(_72_)
);

NAND3X1 _3706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_72_),
    .C(_69_),
    .Y(_73_)
);

INVX1 _3707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .Y(_74_)
);

NAND3X1 _3708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_67_),
    .B(_61_),
    .C(_66_),
    .Y(_75_)
);

OAI21X1 _3709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_70_),
    .B(_71_),
    .C(_68_),
    .Y(_76_)
);

NAND3X1 _3710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_75_),
    .B(_74_),
    .C(_76_),
    .Y(_77_)
);

NAND2X1 _3711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_77_),
    .B(_73_),
    .Y(_78_)
);

OAI21X1 _3712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_14_),
    .B(_2734_),
    .C(_7_),
    .Y(_79_)
);

NAND2X1 _3713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[10]),
    .Y(_80_)
);

NAND2X1 _3714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf3),
    .B(bregp1[11]),
    .Y(_81_)
);

NAND2X1 _3715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf2),
    .B(bregp1[12]),
    .Y(_82_)
);

OR2X2 _3716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_82_),
    .Y(_83_)
);

INVX1 _3717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[12]),
    .Y(_84_)
);

OAI21X1 _3718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_84_),
    .C(_81_),
    .Y(_85_)
);

NAND3X1 _3719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .B(_85_),
    .C(_83_),
    .Y(_86_)
);

INVX1 _3720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_80_),
    .Y(_87_)
);

NAND2X1 _3721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf2),
    .B(bregp1[12]),
    .Y(_88_)
);

NOR2X1 _3722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2727_),
    .B(_88_),
    .Y(_89_)
);

AND2X2 _3723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_81_),
    .B(_82_),
    .Y(_90_)
);

OAI21X1 _3724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_90_),
    .B(_89_),
    .C(_87_),
    .Y(_91_)
);

AND2X2 _3725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_86_),
    .B(_91_),
    .Y(_92_)
);

OAI21X1 _3726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2739_),
    .B(_2736_),
    .C(_2737_),
    .Y(_93_)
);

NAND2X1 _3727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[13]),
    .Y(_94_)
);

NAND3X1 _3728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf3),
    .B(bregp1[14]),
    .C(\preg[7] [22]),
    .Y(_95_)
);

INVX1 _3729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .Y(_96_)
);

AOI21X1 _3730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf2),
    .B(bregp1[14]),
    .C(\preg[7] [22]),
    .Y(_97_)
);

NOR3X1 _3731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .B(_97_),
    .C(_96_),
    .Y(_98_)
);

INVX1 _3732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_94_),
    .Y(_99_)
);

INVX1 _3733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .Y(_100_)
);

AOI21X1 _3734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_95_),
    .B(_100_),
    .C(_99_),
    .Y(_101_)
);

OAI21X1 _3735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_101_),
    .C(_93_),
    .Y(_102_)
);

INVX2 _3736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .Y(_103_)
);

NAND3X1 _3737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_99_),
    .B(_95_),
    .C(_100_),
    .Y(_104_)
);

OAI21X1 _3738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_96_),
    .B(_97_),
    .C(_94_),
    .Y(_105_)
);

NAND3X1 _3739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_105_),
    .C(_103_),
    .Y(_106_)
);

AOI21X1 _3740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_102_),
    .B(_106_),
    .C(_92_),
    .Y(_107_)
);

NAND2X1 _3741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_91_),
    .B(_86_),
    .Y(_108_)
);

NAND3X1 _3742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_93_),
    .B(_104_),
    .C(_105_),
    .Y(_109_)
);

OAI21X1 _3743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_98_),
    .B(_101_),
    .C(_103_),
    .Y(_110_)
);

AOI21X1 _3744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_109_),
    .B(_110_),
    .C(_108_),
    .Y(_111_)
);

OAI21X1 _3745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_111_),
    .C(_79_),
    .Y(_112_)
);

AOI21X1 _3746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_8_),
    .B(_6_),
    .C(_13_),
    .Y(_113_)
);

NAND3X1 _3747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_109_),
    .C(_110_),
    .Y(_114_)
);

NOR3X1 _3748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_101_),
    .B(_103_),
    .C(_98_),
    .Y(_115_)
);

AOI21X1 _3749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_104_),
    .B(_105_),
    .C(_93_),
    .Y(_116_)
);

OAI21X1 _3750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_115_),
    .B(_116_),
    .C(_92_),
    .Y(_117_)
);

NAND3X1 _3751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(_113_),
    .C(_117_),
    .Y(_118_)
);

AOI21X1 _3752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_112_),
    .B(_118_),
    .C(_78_),
    .Y(_119_)
);

NAND3X1 _3753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_74_),
    .B(_69_),
    .C(_72_),
    .Y(_120_)
);

NAND3X1 _3754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_54_),
    .B(_75_),
    .C(_76_),
    .Y(_121_)
);

NAND2X1 _3755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_121_),
    .B(_120_),
    .Y(_122_)
);

NAND3X1 _3756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_79_),
    .B(_114_),
    .C(_117_),
    .Y(_123_)
);

OAI21X1 _3757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_111_),
    .C(_113_),
    .Y(_124_)
);

AOI21X1 _3758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_125_)
);

OAI21X1 _3759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_125_),
    .C(_53_),
    .Y(_126_)
);

NOR3X1 _3760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_9_),
    .B(_5_),
    .C(_11_),
    .Y(_127_)
);

AOI21X1 _3761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_20_),
    .B(_22_),
    .C(_127_),
    .Y(_128_)
);

NAND3X1 _3762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_123_),
    .B(_124_),
    .C(_122_),
    .Y(_130_)
);

NOR3X1 _3763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_107_),
    .B(_111_),
    .C(_113_),
    .Y(_131_)
);

AOI21X1 _3764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_114_),
    .B(_117_),
    .C(_79_),
    .Y(_132_)
);

OAI21X1 _3765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_131_),
    .B(_132_),
    .C(_78_),
    .Y(_133_)
);

NAND3X1 _3766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_128_),
    .C(_133_),
    .Y(_134_)
);

AOI21X1 _3767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_126_),
    .B(_134_),
    .C(_51_),
    .Y(_135_)
);

INVX2 _3768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .Y(_136_)
);

NAND3X1 _3769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_53_),
    .C(_133_),
    .Y(_137_)
);

OAI21X1 _3770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_125_),
    .C(_128_),
    .Y(_138_)
);

AOI21X1 _3771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_138_),
    .B(_137_),
    .C(_136_),
    .Y(_139_)
);

OAI21X1 _3772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_135_),
    .B(_139_),
    .C(_49_),
    .Y(_141_)
);

AOI21X1 _3773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2694_),
    .B(_32_),
    .C(_38_),
    .Y(_142_)
);

NAND3X1 _3774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_138_),
    .C(_137_),
    .Y(_143_)
);

NAND3X1 _3775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_51_),
    .B(_126_),
    .C(_134_),
    .Y(_144_)
);

NAND3X1 _3776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_143_),
    .B(_144_),
    .C(_142_),
    .Y(_145_)
);

AOI22X1 _3777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_145_),
    .C(_48_),
    .D(_44_),
    .Y(_146_)
);

NAND2X1 _3778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_48_),
    .Y(_147_)
);

NAND2X1 _3779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_141_),
    .B(_145_),
    .Y(_148_)
);

NOR2X1 _3780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_147_),
    .Y(_149_)
);

NOR2X1 _3781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_149_),
    .Y(\partials[15] [22])
);

NAND3X1 _3782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_143_),
    .B(_144_),
    .C(_49_),
    .Y(_150_)
);

NAND2X1 _3783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_148_),
    .B(_147_),
    .Y(_151_)
);

AOI21X1 _3784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_130_),
    .B(_133_),
    .C(_53_),
    .Y(_152_)
);

OAI21X1 _3785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_152_),
    .B(_51_),
    .C(_137_),
    .Y(_153_)
);

NAND2X1 _3786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_69_),
    .B(_73_),
    .Y(_154_)
);

INVX1 _3787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .Y(_155_)
);

OAI21X1 _3788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_78_),
    .B(_132_),
    .C(_123_),
    .Y(_156_)
);

AND2X2 _3789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_61_),
    .B(_58_),
    .Y(_157_)
);

NAND2X1 _3790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .B(bregp1[8]),
    .Y(_158_)
);

AOI22X1 _3791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf0),
    .B(bregp1[10]),
    .C(aregp1[14]),
    .D(bregp1[9]),
    .Y(_159_)
);

NAND2X1 _3792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[10]),
    .Y(_161_)
);

NOR2X1 _3793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_161_),
    .Y(_162_)
);

OAI21X1 _3794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_159_),
    .C(_158_),
    .Y(_163_)
);

INVX1 _3795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .Y(_164_)
);

INVX1 _3796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_159_),
    .Y(_165_)
);

OR2X2 _3797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_59_),
    .B(_161_),
    .Y(_166_)
);

NAND3X1 _3798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_164_),
    .B(_165_),
    .C(_166_),
    .Y(_167_)
);

OAI21X1 _3799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_90_),
    .B(_80_),
    .C(_83_),
    .Y(_168_)
);

NAND3X1 _3800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_163_),
    .B(_168_),
    .C(_167_),
    .Y(_169_)
);

AOI21X1 _3801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_165_),
    .B(_166_),
    .C(_164_),
    .Y(_170_)
);

NOR3X1 _3802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_158_),
    .B(_159_),
    .C(_162_),
    .Y(_172_)
);

AOI21X1 _3803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_87_),
    .B(_85_),
    .C(_89_),
    .Y(_173_)
);

OAI21X1 _3804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_172_),
    .C(_173_),
    .Y(_174_)
);

NAND3X1 _3805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_174_),
    .C(_157_),
    .Y(_175_)
);

OAI21X1 _3806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2702_),
    .B(_56_),
    .C(_61_),
    .Y(_176_)
);

NAND3X1 _3807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_173_),
    .B(_163_),
    .C(_167_),
    .Y(_177_)
);

OAI21X1 _3808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_170_),
    .B(_172_),
    .C(_168_),
    .Y(_178_)
);

NAND3X1 _3809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_177_),
    .B(_176_),
    .C(_178_),
    .Y(_179_)
);

AND2X2 _3810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_175_),
    .B(_179_),
    .Y(_180_)
);

OAI21X1 _3811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_92_),
    .B(_116_),
    .C(_109_),
    .Y(_181_)
);

NAND2X1 _3812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[11]),
    .Y(_183_)
);

NAND2X1 _3813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf1),
    .B(bregp1[13]),
    .Y(_184_)
);

AOI21X1 _3814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf1),
    .B(bregp1[12]),
    .C(_184_),
    .Y(_185_)
);

AOI21X1 _3815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf0),
    .B(bregp1[13]),
    .C(_88_),
    .Y(_186_)
);

OAI21X1 _3816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_186_),
    .C(_183_),
    .Y(_187_)
);

INVX1 _3817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_183_),
    .Y(_188_)
);

NOR2X1 _3818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_184_),
    .Y(_189_)
);

AND2X2 _3819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_184_),
    .Y(_190_)
);

OAI21X1 _3820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_190_),
    .B(_189_),
    .C(_188_),
    .Y(_191_)
);

AND2X2 _3821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_191_),
    .B(_187_),
    .Y(_192_)
);

OAI21X1 _3822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_97_),
    .B(_94_),
    .C(_95_),
    .Y(_194_)
);

NAND2X1 _3823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[14]),
    .Y(_195_)
);

NAND3X1 _3824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf1),
    .B(bregp1[15]),
    .C(\preg[7] [23]),
    .Y(_196_)
);

INVX2 _3825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .Y(_197_)
);

AOI21X1 _3826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_8_bF$buf0),
    .B(bregp1[15]),
    .C(\preg[7] [23]),
    .Y(_198_)
);

NOR3X1 _3827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_198_),
    .C(_197_),
    .Y(_199_)
);

INVX2 _3828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .Y(_200_)
);

INVX1 _3829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .Y(_201_)
);

AOI21X1 _3830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_196_),
    .B(_201_),
    .C(_200_),
    .Y(_202_)
);

OAI21X1 _3831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_202_),
    .C(_194_),
    .Y(_203_)
);

INVX1 _3832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .Y(_205_)
);

NAND3X1 _3833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_196_),
    .C(_201_),
    .Y(_206_)
);

OAI21X1 _3834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_197_),
    .B(_198_),
    .C(_195_),
    .Y(_207_)
);

NAND3X1 _3835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_206_),
    .B(_207_),
    .C(_205_),
    .Y(_208_)
);

AOI21X1 _3836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_208_),
    .B(_203_),
    .C(_192_),
    .Y(_209_)
);

NAND2X1 _3837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_187_),
    .B(_191_),
    .Y(_210_)
);

NAND3X1 _3838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_194_),
    .B(_206_),
    .C(_207_),
    .Y(_211_)
);

OAI21X1 _3839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_202_),
    .C(_205_),
    .Y(_212_)
);

AOI21X1 _3840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_212_),
    .C(_210_),
    .Y(_213_)
);

OAI21X1 _3841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_213_),
    .C(_181_),
    .Y(_214_)
);

AOI21X1 _3842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_108_),
    .B(_110_),
    .C(_115_),
    .Y(_216_)
);

NAND3X1 _3843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_210_),
    .B(_211_),
    .C(_212_),
    .Y(_217_)
);

NAND3X1 _3844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_203_),
    .B(_208_),
    .C(_192_),
    .Y(_218_)
);

NAND3X1 _3845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_218_),
    .C(_216_),
    .Y(_219_)
);

AOI21X1 _3846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_219_),
    .C(_180_),
    .Y(_220_)
);

NAND2X1 _3847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_179_),
    .B(_175_),
    .Y(_221_)
);

NAND3X1 _3848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_217_),
    .B(_218_),
    .C(_181_),
    .Y(_222_)
);

OAI21X1 _3849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_209_),
    .B(_213_),
    .C(_216_),
    .Y(_223_)
);

AOI21X1 _3850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_223_),
    .B(_222_),
    .C(_221_),
    .Y(_224_)
);

OAI21X1 _3851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_224_),
    .C(_156_),
    .Y(_225_)
);

AOI21X1 _3852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_124_),
    .B(_122_),
    .C(_131_),
    .Y(_226_)
);

NAND3X1 _3853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_221_),
    .B(_222_),
    .C(_223_),
    .Y(_227_)
);

NAND3X1 _3854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_214_),
    .B(_219_),
    .C(_180_),
    .Y(_228_)
);

NAND3X1 _3855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_226_),
    .C(_228_),
    .Y(_229_)
);

AOI21X1 _3856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_229_),
    .B(_225_),
    .C(_155_),
    .Y(_230_)
);

NAND3X1 _3857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_227_),
    .B(_156_),
    .C(_228_),
    .Y(_231_)
);

OAI21X1 _3858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_220_),
    .B(_224_),
    .C(_226_),
    .Y(_232_)
);

AOI21X1 _3859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_232_),
    .C(_154_),
    .Y(_233_)
);

OAI21X1 _3860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_233_),
    .C(_153_),
    .Y(_234_)
);

NOR3X1 _3861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_119_),
    .B(_125_),
    .C(_128_),
    .Y(_235_)
);

AOI21X1 _3862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_136_),
    .B(_138_),
    .C(_235_),
    .Y(_237_)
);

NAND3X1 _3863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_154_),
    .B(_231_),
    .C(_232_),
    .Y(_238_)
);

NAND3X1 _3864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_155_),
    .B(_229_),
    .C(_225_),
    .Y(_239_)
);

NAND3X1 _3865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_239_),
    .C(_237_),
    .Y(_240_)
);

NAND2X1 _3866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_240_),
    .B(_234_),
    .Y(_241_)
);

NAND3X1 _3867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .B(_241_),
    .C(_151_),
    .Y(_242_)
);

INVX1 _3868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_150_),
    .Y(_243_)
);

INVX1 _3869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_241_),
    .Y(_244_)
);

OAI21X1 _3870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_146_),
    .B(_243_),
    .C(_244_),
    .Y(_245_)
);

NAND2X1 _3871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_245_),
    .B(_242_),
    .Y(\partials[15] [23])
);

AND2X2 _3872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2688_),
    .B(_2684_),
    .Y(_247_)
);

AOI22X1 _3873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_234_),
    .B(_240_),
    .C(_141_),
    .D(_145_),
    .Y(_248_)
);

NAND3X1 _3874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_247_),
    .C(_42_),
    .Y(_249_)
);

NOR3X1 _3875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_249_),
    .B(_2604_),
    .C(_2229_),
    .Y(_250_)
);

OAI21X1 _3876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_41_),
    .B(_2688_),
    .C(_45_),
    .Y(_251_)
);

NOR2X1 _3877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_233_),
    .Y(_252_)
);

OAI21X1 _3878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_235_),
    .B(_135_),
    .C(_252_),
    .Y(_253_)
);

AOI21X1 _3879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_239_),
    .C(_153_),
    .Y(_254_)
);

OAI21X1 _3880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_254_),
    .B(_150_),
    .C(_253_),
    .Y(_255_)
);

AOI21X1 _3881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_248_),
    .B(_251_),
    .C(_255_),
    .Y(_256_)
);

OAI21X1 _3882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2603_),
    .B(_249_),
    .C(_256_),
    .Y(_258_)
);

NOR2X1 _3883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_258_),
    .B(_250_),
    .Y(_259_)
);

NAND2X1 _3884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_231_),
    .B(_238_),
    .Y(_260_)
);

NAND3X1 _3885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_176_),
    .C(_174_),
    .Y(_261_)
);

NAND2X1 _3886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_169_),
    .B(_261_),
    .Y(_262_)
);

NAND2X1 _3887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_222_),
    .B(_227_),
    .Y(_263_)
);

NOR2X1 _3888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_162_),
    .B(_172_),
    .Y(_264_)
);

NAND2X1 _3889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .B(bregp1[10]),
    .Y(_265_)
);

INVX2 _3890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_265_),
    .Y(_266_)
);

AOI22X1 _3891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[10]),
    .C(aregp1[15]),
    .D(bregp1[9]),
    .Y(_267_)
);

AOI21X1 _3892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_266_),
    .B(_57_),
    .C(_267_),
    .Y(_269_)
);

OAI21X1 _3893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_185_),
    .B(_186_),
    .C(_188_),
    .Y(_270_)
);

OAI21X1 _3894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_184_),
    .C(_270_),
    .Y(_271_)
);

XNOR2X1 _3895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_271_),
    .B(_269_),
    .Y(_272_)
);

OR2X2 _3896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_264_),
    .Y(_273_)
);

NAND2X1 _3897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_264_),
    .B(_272_),
    .Y(_274_)
);

AND2X2 _3898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_273_),
    .B(_274_),
    .Y(_275_)
);

NAND2X1 _3899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_217_),
    .Y(_276_)
);

NAND2X1 _3900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf3),
    .B(bregp1[11]),
    .Y(_277_)
);

NAND2X1 _3901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[13]),
    .Y(_278_)
);

NOR2X1 _3902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_278_),
    .Y(_280_)
);

AOI22X1 _3903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf0),
    .B(bregp1[13]),
    .C(aregp1[12]),
    .D(bregp1[12]),
    .Y(_281_)
);

OAI21X1 _3904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_280_),
    .B(_281_),
    .C(_277_),
    .Y(_282_)
);

NOR2X1 _3905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_281_),
    .B(_280_),
    .Y(_283_)
);

NAND3X1 _3906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf2),
    .B(bregp1[11]),
    .C(_283_),
    .Y(_284_)
);

NAND2X1 _3907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_282_),
    .B(_284_),
    .Y(_285_)
);

OAI21X1 _3908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_198_),
    .B(_195_),
    .C(_196_),
    .Y(_286_)
);

NAND2X1 _3909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_10_bF$buf3),
    .B(bregp1[15]),
    .Y(_287_)
);

INVX1 _3910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .Y(_288_)
);

AOI22X1 _3911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[9]),
    .B(bregp1[15]),
    .C(aregp1_10_bF$buf2),
    .D(bregp1[14]),
    .Y(_289_)
);

AOI21X1 _3912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_200_),
    .B(_288_),
    .C(_289_),
    .Y(_291_)
);

XNOR2X1 _3913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_291_),
    .B(_286_),
    .Y(_292_)
);

XOR2X1 _3914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_292_),
    .Y(_293_)
);

NAND2X1 _3915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_293_),
    .Y(_294_)
);

XNOR2X1 _3916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_292_),
    .Y(_295_)
);

NAND3X1 _3917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_211_),
    .B(_217_),
    .C(_295_),
    .Y(_296_)
);

NAND3X1 _3918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_296_),
    .C(_275_),
    .Y(_297_)
);

NAND2X1 _3919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_274_),
    .B(_273_),
    .Y(_298_)
);

INVX1 _3920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .Y(_299_)
);

NOR2X1 _3921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_276_),
    .B(_293_),
    .Y(_300_)
);

OAI21X1 _3922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_299_),
    .B(_300_),
    .C(_298_),
    .Y(_302_)
);

NAND3X1 _3923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .B(_297_),
    .C(_302_),
    .Y(_303_)
);

INVX2 _3924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_263_),
    .Y(_304_)
);

NAND2X1 _3925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_296_),
    .Y(_305_)
);

NOR2X1 _3926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_305_),
    .Y(_306_)
);

AOI21X1 _3927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_294_),
    .B(_296_),
    .C(_275_),
    .Y(_307_)
);

OAI21X1 _3928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_307_),
    .C(_304_),
    .Y(_308_)
);

NAND3X1 _3929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .B(_303_),
    .C(_308_),
    .Y(_309_)
);

INVX2 _3930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_262_),
    .Y(_310_)
);

NOR3X1 _3931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_304_),
    .B(_307_),
    .C(_306_),
    .Y(_311_)
);

AOI21X1 _3932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_302_),
    .C(_263_),
    .Y(_313_)
);

OAI21X1 _3933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_311_),
    .B(_313_),
    .C(_310_),
    .Y(_314_)
);

NAND3X1 _3934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .B(_309_),
    .C(_314_),
    .Y(_315_)
);

INVX1 _3935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_260_),
    .Y(_316_)
);

OAI21X1 _3936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_306_),
    .B(_307_),
    .C(_263_),
    .Y(_317_)
);

NAND3X1 _3937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_297_),
    .B(_304_),
    .C(_302_),
    .Y(_318_)
);

AOI21X1 _3938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_318_),
    .B(_317_),
    .C(_310_),
    .Y(_319_)
);

AOI21X1 _3939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_303_),
    .B(_308_),
    .C(_262_),
    .Y(_320_)
);

OAI21X1 _3940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_319_),
    .B(_320_),
    .C(_316_),
    .Y(_321_)
);

AND2X2 _3941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_315_),
    .B(_321_),
    .Y(_322_)
);

XNOR2X1 _3942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_322_),
    .Y(\partials[15] [24])
);

NAND2X1 _3943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_321_),
    .B(_315_),
    .Y(_324_)
);

OAI21X1 _3944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_324_),
    .C(_315_),
    .Y(_325_)
);

OAI21X1 _3945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_313_),
    .B(_310_),
    .C(_303_),
    .Y(_326_)
);

INVX1 _3946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .Y(_327_)
);

NAND2X1 _3947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_269_),
    .B(_271_),
    .Y(_328_)
);

OAI21X1 _3948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_272_),
    .B(_264_),
    .C(_328_),
    .Y(_329_)
);

AOI21X1 _3949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_296_),
    .B(_275_),
    .C(_299_),
    .Y(_330_)
);

OAI21X1 _3950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_199_),
    .B(_197_),
    .C(_291_),
    .Y(_331_)
);

OAI21X1 _3951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_285_),
    .B(_292_),
    .C(_331_),
    .Y(_332_)
);

NAND2X1 _3952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[11]),
    .Y(_333_)
);

NAND2X1 _3953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf1),
    .B(bregp1[12]),
    .Y(_334_)
);

NOR2X1 _3954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_334_),
    .Y(_335_)
);

AOI22X1 _3955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[13]),
    .C(aregp1_13_bF$buf0),
    .D(bregp1[12]),
    .Y(_336_)
);

OAI21X1 _3956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_335_),
    .B(_336_),
    .C(_333_),
    .Y(_337_)
);

INVX1 _3957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_333_),
    .Y(_338_)
);

NOR2X1 _3958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_336_),
    .B(_335_),
    .Y(_339_)
);

NAND2X1 _3959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_338_),
    .B(_339_),
    .Y(_340_)
);

NAND2X1 _3960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_337_),
    .B(_340_),
    .Y(_341_)
);

NAND2X1 _3961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_11_bF$buf3),
    .B(bregp1[14]),
    .Y(_342_)
);

NOR2X1 _3962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_342_),
    .Y(_345_)
);

AND2X2 _3963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_342_),
    .Y(_346_)
);

OAI22X1 _3964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_195_),
    .B(_287_),
    .C(_346_),
    .D(_345_),
    .Y(_347_)
);

NAND3X1 _3965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_342_),
    .B(_200_),
    .C(_288_),
    .Y(_348_)
);

NAND2X1 _3966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .B(_347_),
    .Y(_349_)
);

XOR2X1 _3967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_349_),
    .Y(_350_)
);

OR2X2 _3968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_350_),
    .B(_332_),
    .Y(_351_)
);

NAND2X1 _3969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_350_),
    .Y(_352_)
);

OAI21X1 _3970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_88_),
    .B(_278_),
    .C(_284_),
    .Y(_353_)
);

OAI21X1 _3971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_2541_),
    .C(_266_),
    .Y(_354_)
);

XNOR2X1 _3972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_354_),
    .Y(_355_)
);

AOI21X1 _3973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_351_),
    .C(_355_),
    .Y(_356_)
);

NOR2X1 _3974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_332_),
    .B(_350_),
    .Y(_357_)
);

INVX2 _3975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .Y(_358_)
);

INVX2 _3976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .Y(_359_)
);

NOR3X1 _3977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_357_),
    .B(_359_),
    .C(_358_),
    .Y(_360_)
);

OAI21X1 _3978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_356_),
    .C(_330_),
    .Y(_361_)
);

OAI21X1 _3979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_298_),
    .B(_300_),
    .C(_294_),
    .Y(_362_)
);

OAI21X1 _3980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_358_),
    .B(_357_),
    .C(_359_),
    .Y(_363_)
);

NAND3X1 _3981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_352_),
    .B(_355_),
    .C(_351_),
    .Y(_364_)
);

NAND3X1 _3982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_362_),
    .B(_364_),
    .C(_363_),
    .Y(_366_)
);

AOI21X1 _3983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_366_),
    .B(_361_),
    .C(_329_),
    .Y(_367_)
);

INVX2 _3984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .Y(_368_)
);

AOI21X1 _3985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_364_),
    .B(_363_),
    .C(_362_),
    .Y(_369_)
);

NOR3X1 _3986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_360_),
    .B(_356_),
    .C(_330_),
    .Y(_370_)
);

NOR3X1 _3987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_368_),
    .B(_369_),
    .C(_370_),
    .Y(_371_)
);

OAI21X1 _3988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_371_),
    .B(_367_),
    .C(_327_),
    .Y(_372_)
);

OAI21X1 _3989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_369_),
    .C(_368_),
    .Y(_373_)
);

NAND3X1 _3990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_366_),
    .C(_361_),
    .Y(_374_)
);

NAND3X1 _3991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_326_),
    .B(_374_),
    .C(_373_),
    .Y(_375_)
);

NAND2X1 _3992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_372_),
    .Y(_377_)
);

XNOR2X1 _3993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_325_),
    .B(_377_),
    .Y(\partials[15] [25])
);

NOR2X1 _3994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_324_),
    .B(_377_),
    .Y(_378_)
);

OAI21X1 _3995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_258_),
    .C(_378_),
    .Y(_379_)
);

NAND2X1 _3996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_375_),
    .B(_315_),
    .Y(_380_)
);

NAND2X1 _3997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_380_),
    .Y(_381_)
);

AOI21X1 _3998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_329_),
    .B(_361_),
    .C(_370_),
    .Y(_382_)
);

OAI21X1 _3999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_357_),
    .B(_359_),
    .C(_352_),
    .Y(_383_)
);

OAI21X1 _4000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_278_),
    .B(_334_),
    .C(_340_),
    .Y(_384_)
);

INVX1 _4001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_348_),
    .Y(_385_)
);

NOR2X1 _4002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_349_),
    .B(_341_),
    .Y(_387_)
);

NAND2X1 _4003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .B(bregp1[11]),
    .Y(_388_)
);

NAND2X1 _4004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf3),
    .B(bregp1[13]),
    .Y(_389_)
);

NAND2X1 _4005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[14]),
    .B(bregp1[12]),
    .Y(_390_)
);

AND2X2 _4006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .Y(_391_)
);

NOR2X1 _4007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .Y(_392_)
);

OAI21X1 _4008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_391_),
    .B(_392_),
    .C(_388_),
    .Y(_393_)
);

INVX1 _4009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_388_),
    .Y(_394_)
);

NOR2X1 _4010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_392_),
    .B(_391_),
    .Y(_395_)
);

NAND2X1 _4011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_394_),
    .B(_395_),
    .Y(_396_)
);

NAND2X1 _4012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_393_),
    .B(_396_),
    .Y(_398_)
);

NAND2X1 _4013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[15]),
    .Y(_399_)
);

NOR2X1 _4014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_342_),
    .B(_399_),
    .Y(_400_)
);

INVX2 _4015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[15]),
    .Y(_401_)
);

NOR2X1 _4016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_652_),
    .B(_401_),
    .Y(_402_)
);

NAND2X1 _4017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[12]),
    .B(bregp1[14]),
    .Y(_403_)
);

INVX1 _4018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .Y(_404_)
);

NOR2X1 _4019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_402_),
    .Y(_405_)
);

OAI22X1 _4020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_287_),
    .B(_342_),
    .C(_405_),
    .D(_400_),
    .Y(_406_)
);

INVX1 _4021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[14]),
    .Y(_407_)
);

NOR2X1 _4022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_365_),
    .B(_407_),
    .Y(_409_)
);

NAND3X1 _4023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_403_),
    .B(_409_),
    .C(_402_),
    .Y(_410_)
);

NAND2X1 _4024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_410_),
    .B(_406_),
    .Y(_411_)
);

XOR2X1 _4025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_411_),
    .Y(_412_)
);

OAI21X1 _4026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_387_),
    .C(_412_),
    .Y(_413_)
);

OAI21X1 _4027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_341_),
    .B(_349_),
    .C(_348_),
    .Y(_414_)
);

INVX1 _4028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .Y(_415_)
);

NAND2X1 _4029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_411_),
    .B(_398_),
    .Y(_416_)
);

OR2X2 _4030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_411_),
    .Y(_417_)
);

NAND2X1 _4031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_416_),
    .B(_417_),
    .Y(_418_)
);

NAND2X1 _4032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_418_),
    .Y(_420_)
);

NAND3X1 _4033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_413_),
    .C(_420_),
    .Y(_421_)
);

INVX2 _4034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .Y(_422_)
);

NOR2X1 _4035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_418_),
    .Y(_423_)
);

NOR2X1 _4036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_414_),
    .B(_412_),
    .Y(_424_)
);

OAI21X1 _4037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_423_),
    .B(_424_),
    .C(_422_),
    .Y(_425_)
);

NAND3X1 _4038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_383_),
    .B(_421_),
    .C(_425_),
    .Y(_426_)
);

AOI21X1 _4039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_355_),
    .B(_351_),
    .C(_358_),
    .Y(_427_)
);

OAI21X1 _4040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_385_),
    .B(_387_),
    .C(_418_),
    .Y(_428_)
);

NAND2X1 _4041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_415_),
    .B(_412_),
    .Y(_429_)
);

AOI21X1 _4042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_429_),
    .B(_428_),
    .C(_422_),
    .Y(_431_)
);

AOI21X1 _4043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_413_),
    .B(_420_),
    .C(_384_),
    .Y(_432_)
);

OAI21X1 _4044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_432_),
    .C(_427_),
    .Y(_433_)
);

OAI21X1 _4045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_353_),
    .B(_57_),
    .C(_266_),
    .Y(_434_)
);

INVX1 _4046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .Y(_435_)
);

NAND3X1 _4047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_435_),
    .B(_433_),
    .C(_426_),
    .Y(_436_)
);

OAI21X1 _4048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_431_),
    .B(_432_),
    .C(_383_),
    .Y(_437_)
);

NAND3X1 _4049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_427_),
    .B(_421_),
    .C(_425_),
    .Y(_438_)
);

NAND3X1 _4050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_434_),
    .B(_437_),
    .C(_438_),
    .Y(_439_)
);

AOI21X1 _4051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_436_),
    .B(_439_),
    .C(_382_),
    .Y(_440_)
);

OAI21X1 _4052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_369_),
    .B(_368_),
    .C(_366_),
    .Y(_442_)
);

AOI21X1 _4053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_437_),
    .B(_438_),
    .C(_434_),
    .Y(_443_)
);

AOI21X1 _4054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_433_),
    .B(_426_),
    .C(_435_),
    .Y(_444_)
);

NOR3X1 _4055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_444_),
    .C(_442_),
    .Y(_445_)
);

NOR2X1 _4056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_440_),
    .B(_445_),
    .Y(_446_)
);

AOI21X1 _4057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_379_),
    .C(_446_),
    .Y(_447_)
);

AND2X2 _4058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_372_),
    .B(_375_),
    .Y(_448_)
);

NAND2X1 _4059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_448_),
    .Y(_449_)
);

OAI21X1 _4060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_449_),
    .C(_381_),
    .Y(_450_)
);

INVX1 _4061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_446_),
    .Y(_451_)
);

NOR2X1 _4062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_451_),
    .B(_450_),
    .Y(_453_)
);

NOR2X1 _4063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_447_),
    .B(_453_),
    .Y(\partials[15] [26])
);

NOR2X1 _4064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_444_),
    .B(_443_),
    .Y(_454_)
);

OAI21X1 _4065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_370_),
    .B(_371_),
    .C(_454_),
    .Y(_455_)
);

AND2X2 _4066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2414_),
    .B(_2601_),
    .Y(_456_)
);

AOI21X1 _4067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_143_),
    .B(_144_),
    .C(_142_),
    .Y(_457_)
);

NOR3X1 _4068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_49_),
    .B(_139_),
    .C(_135_),
    .Y(_458_)
);

AOI21X1 _4069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_238_),
    .B(_239_),
    .C(_237_),
    .Y(_459_)
);

NOR3X1 _4070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_230_),
    .B(_233_),
    .C(_153_),
    .Y(_460_)
);

OAI22X1 _4071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_460_),
    .B(_459_),
    .C(_457_),
    .D(_458_),
    .Y(_461_)
);

NOR3X1 _4072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2689_),
    .B(_46_),
    .C(_461_),
    .Y(_463_)
);

NAND3X1 _4073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_456_),
    .B(_463_),
    .C(_2319_),
    .Y(_464_)
);

NOR3X1 _4074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2400_),
    .B(_2397_),
    .C(_2403_),
    .Y(_465_)
);

OAI21X1 _4075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2400_),
    .B(_2397_),
    .C(_2403_),
    .Y(_466_)
);

OAI21X1 _4076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2320_),
    .B(_465_),
    .C(_466_),
    .Y(_467_)
);

AOI21X1 _4077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2500_),
    .B(_2503_),
    .C(_2499_),
    .Y(_468_)
);

NOR3X1 _4078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2494_),
    .B(_2497_),
    .C(_2416_),
    .Y(_469_)
);

AOI21X1 _4079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2586_),
    .B(_2590_),
    .C(_2592_),
    .Y(_470_)
);

NOR3X1 _4080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2595_),
    .B(_2596_),
    .C(_2509_),
    .Y(_471_)
);

OAI22X1 _4081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_469_),
    .B(_468_),
    .C(_470_),
    .D(_471_),
    .Y(_472_)
);

NAND2X1 _4082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2597_),
    .B(_2602_),
    .Y(_474_)
);

OAI21X1 _4083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_467_),
    .B(_472_),
    .C(_474_),
    .Y(_475_)
);

AOI21X1 _4084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_153_),
    .B(_252_),
    .C(_243_),
    .Y(_476_)
);

OAI22X1 _4085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_44_),
    .B(_461_),
    .C(_476_),
    .D(_254_),
    .Y(_477_)
);

AOI21X1 _4086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_463_),
    .B(_475_),
    .C(_477_),
    .Y(_478_)
);

AOI21X1 _4087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_478_),
    .C(_449_),
    .Y(_479_)
);

OAI21X1 _4088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_377_),
    .B(_315_),
    .C(_375_),
    .Y(_480_)
);

OAI21X1 _4089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_479_),
    .B(_480_),
    .C(_451_),
    .Y(_481_)
);

AOI21X1 _4090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_421_),
    .B(_425_),
    .C(_383_),
    .Y(_482_)
);

OAI21X1 _4091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_482_),
    .B(_434_),
    .C(_426_),
    .Y(_483_)
);

AOI21X1 _4092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_384_),
    .B(_420_),
    .C(_423_),
    .Y(_484_)
);

OAI21X1 _4093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_389_),
    .B(_390_),
    .C(_396_),
    .Y(_485_)
);

OAI21X1 _4094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_398_),
    .B(_411_),
    .C(_410_),
    .Y(_486_)
);

INVX2 _4095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(bregp1[13]),
    .Y(_487_)
);

NOR2X1 _4096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2146_),
    .B(_487_),
    .Y(_488_)
);

INVX2 _4097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_488_),
    .Y(_489_)
);

OAI22X1 _4098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_487_),
    .C(_2146_),
    .D(_84_),
    .Y(_490_)
);

OAI21X1 _4099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_390_),
    .C(_490_),
    .Y(_491_)
);

NAND2X1 _4100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1_13_bF$buf2),
    .B(bregp1[14]),
    .Y(_492_)
);

XOR2X1 _4101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_399_),
    .B(_492_),
    .Y(_493_)
);

XOR2X1 _4102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_493_),
    .B(_400_),
    .Y(_495_)
);

XNOR2X1 _4103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_495_),
    .B(_491_),
    .Y(_496_)
);

OR2X2 _4104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_486_),
    .Y(_497_)
);

NAND2X1 _4105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .B(_496_),
    .Y(_498_)
);

AOI21X1 _4106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_498_),
    .B(_497_),
    .C(_485_),
    .Y(_499_)
);

INVX2 _4107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .Y(_500_)
);

NOR2X1 _4108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_486_),
    .B(_496_),
    .Y(_501_)
);

AND2X2 _4109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_496_),
    .B(_486_),
    .Y(_502_)
);

NOR3X1 _4110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_500_),
    .C(_502_),
    .Y(_503_)
);

OAI21X1 _4111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_503_),
    .B(_499_),
    .C(_484_),
    .Y(_504_)
);

OAI21X1 _4112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_424_),
    .B(_422_),
    .C(_413_),
    .Y(_507_)
);

OAI21X1 _4113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_502_),
    .B(_501_),
    .C(_500_),
    .Y(_508_)
);

NAND3X1 _4114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_485_),
    .B(_498_),
    .C(_497_),
    .Y(_509_)
);

NAND3X1 _4115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_508_),
    .B(_509_),
    .C(_507_),
    .Y(_510_)
);

NAND2X1 _4116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_510_),
    .Y(_511_)
);

XNOR2X1 _4117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_483_),
    .B(_511_),
    .Y(_512_)
);

NAND3X1 _4118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .B(_512_),
    .C(_481_),
    .Y(_513_)
);

INVX1 _4119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_455_),
    .Y(_514_)
);

NAND3X1 _4120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_426_),
    .B(_511_),
    .C(_436_),
    .Y(_515_)
);

NAND3X1 _4121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_504_),
    .B(_510_),
    .C(_483_),
    .Y(_516_)
);

NAND2X1 _4122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_516_),
    .Y(_517_)
);

OAI21X1 _4123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_447_),
    .B(_514_),
    .C(_517_),
    .Y(_518_)
);

NAND2X1 _4124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_518_),
    .B(_513_),
    .Y(\partials[15] [27])
);

OAI21X1 _4125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_445_),
    .B(_440_),
    .C(_512_),
    .Y(_519_)
);

NOR3X1 _4126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_519_),
    .B(_324_),
    .C(_377_),
    .Y(_520_)
);

OAI21X1 _4127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_250_),
    .B(_258_),
    .C(_520_),
    .Y(_521_)
);

OAI21X1 _4128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_443_),
    .B(_444_),
    .C(_442_),
    .Y(_522_)
);

NAND2X1 _4129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_382_),
    .B(_454_),
    .Y(_523_)
);

AOI21X1 _4130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_522_),
    .B(_523_),
    .C(_517_),
    .Y(_524_)
);

NAND2X1 _4131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_516_),
    .B(_455_),
    .Y(_525_)
);

AOI22X1 _4132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_525_),
    .C(_480_),
    .D(_524_),
    .Y(_528_)
);

INVX1 _4133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_510_),
    .Y(_529_)
);

OAI21X1 _4134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_501_),
    .B(_500_),
    .C(_498_),
    .Y(_530_)
);

OR2X2 _4135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_489_),
    .B(_390_),
    .Y(_531_)
);

INVX2 _4136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_531_),
    .Y(_532_)
);

NOR2X1 _4137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_493_),
    .Y(_533_)
);

NAND2X1 _4138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_400_),
    .B(_493_),
    .Y(_534_)
);

OAI21X1 _4139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_533_),
    .B(_491_),
    .C(_534_),
    .Y(_535_)
);

INVX1 _4140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_492_),
    .Y(_536_)
);

NOR2X1 _4141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_401_),
    .Y(_537_)
);

NAND2X1 _4142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_536_),
    .B(_537_),
    .Y(_539_)
);

INVX1 _4143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_539_),
    .Y(_540_)
);

NOR2X1 _4144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2142_),
    .B(_401_),
    .Y(_541_)
);

NOR2X1 _4145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2065_),
    .B(_407_),
    .Y(_542_)
);

NOR2X1 _4146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_541_),
    .B(_542_),
    .Y(_543_)
);

OAI22X1 _4147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_399_),
    .B(_492_),
    .C(_540_),
    .D(_543_),
    .Y(_544_)
);

INVX1 _4148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .Y(_545_)
);

NAND3X1 _4149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_404_),
    .B(_541_),
    .C(_545_),
    .Y(_546_)
);

NAND2X1 _4150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_546_),
    .B(_544_),
    .Y(_547_)
);

OAI21X1 _4151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2146_),
    .B(_487_),
    .C(_547_),
    .Y(_548_)
);

OR2X2 _4152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_489_),
    .Y(_550_)
);

NAND2X1 _4153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_548_),
    .B(_550_),
    .Y(_551_)
);

XNOR2X1 _4154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_551_),
    .B(_535_),
    .Y(_552_)
);

XNOR2X1 _4155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_552_),
    .B(_532_),
    .Y(_553_)
);

XNOR2X1 _4156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_553_),
    .B(_530_),
    .Y(_554_)
);

NOR2X1 _4157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_554_),
    .Y(_555_)
);

NAND2X1 _4158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_529_),
    .B(_554_),
    .Y(_556_)
);

INVX2 _4159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .Y(_557_)
);

OR2X2 _4160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_557_),
    .B(_555_),
    .Y(_558_)
);

AOI21X1 _4161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_521_),
    .C(_558_),
    .Y(_559_)
);

NAND3X1 _4162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_322_),
    .B(_524_),
    .C(_448_),
    .Y(_561_)
);

OAI21X1 _4163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_259_),
    .B(_561_),
    .C(_528_),
    .Y(_562_)
);

NOR2X1 _4164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_555_),
    .B(_557_),
    .Y(_563_)
);

NOR2X1 _4165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_563_),
    .B(_562_),
    .Y(_564_)
);

NOR2X1 _4166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_564_),
    .Y(\partials[15] [28])
);

AOI21X1 _4167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_464_),
    .B(_478_),
    .C(_561_),
    .Y(_565_)
);

NAND2X1 _4168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_515_),
    .B(_525_),
    .Y(_566_)
);

OAI21X1 _4169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_381_),
    .B(_519_),
    .C(_566_),
    .Y(_567_)
);

OAI21X1 _4170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_567_),
    .C(_563_),
    .Y(_568_)
);

INVX1 _4171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_530_),
    .Y(_569_)
);

OR2X2 _4172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_553_),
    .B(_569_),
    .Y(_571_)
);

NAND3X1 _4173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_535_),
    .B(_548_),
    .C(_550_),
    .Y(_572_)
);

NAND2X1 _4174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_532_),
    .B(_552_),
    .Y(_573_)
);

NAND2X1 _4175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_572_),
    .B(_573_),
    .Y(_574_)
);

OAI21X1 _4176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_547_),
    .B(_489_),
    .C(_546_),
    .Y(_575_)
);

NAND2X1 _4177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .B(bregp1[15]),
    .Y(_576_)
);

NOR2X1 _4178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_576_),
    .B(_545_),
    .Y(_577_)
);

AOI21X1 _4179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(aregp1[15]),
    .B(bregp1[14]),
    .C(_537_),
    .Y(_578_)
);

OAI21X1 _4180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_578_),
    .C(_539_),
    .Y(_579_)
);

NOR2X1 _4181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_578_),
    .Y(_580_)
);

NAND2X1 _4182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_540_),
    .B(_580_),
    .Y(_582_)
);

AND2X2 _4183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_582_),
    .B(_579_),
    .Y(_583_)
);

XOR2X1 _4184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_583_),
    .B(_575_),
    .Y(_584_)
);

XOR2X1 _4185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_574_),
    .B(_584_),
    .Y(_585_)
);

XNOR2X1 _4186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .B(_571_),
    .Y(_586_)
);

NAND3X1 _4187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_556_),
    .B(_586_),
    .C(_568_),
    .Y(_587_)
);

INVX2 _4188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .Y(_588_)
);

OAI21X1 _4189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_559_),
    .B(_557_),
    .C(_588_),
    .Y(_589_)
);

NAND2X1 _4190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_589_),
    .B(_587_),
    .Y(\partials[15] [29])
);

NOR2X1 _4191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_558_),
    .Y(_590_)
);

OAI21X1 _4192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_565_),
    .B(_567_),
    .C(_590_),
    .Y(_592_)
);

INVX1 _4193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_585_),
    .Y(_593_)
);

OR2X2 _4194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_593_),
    .B(_571_),
    .Y(_594_)
);

OAI21X1 _4195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_588_),
    .B(_556_),
    .C(_594_),
    .Y(_595_)
);

INVX1 _4196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_595_),
    .Y(_596_)
);

OAI21X1 _4197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_542_),
    .B(_576_),
    .C(_582_),
    .Y(_597_)
);

NAND2X1 _4198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_575_),
    .B(_583_),
    .Y(_598_)
);

NAND2X1 _4199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_584_),
    .B(_574_),
    .Y(_599_)
);

NAND2X1 _4200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_598_),
    .B(_599_),
    .Y(_600_)
);

AND2X2 _4201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_600_),
    .B(_597_),
    .Y(_601_)
);

NOR2X1 _4202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_597_),
    .B(_600_),
    .Y(_603_)
);

NOR2X1 _4203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_603_),
    .B(_601_),
    .Y(_604_)
);

NAND3X1 _4204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_596_),
    .B(_604_),
    .C(_592_),
    .Y(_605_)
);

NAND2X1 _4205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_586_),
    .B(_563_),
    .Y(_606_)
);

AOI21X1 _4206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_528_),
    .B(_521_),
    .C(_606_),
    .Y(_607_)
);

INVX1 _4207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_604_),
    .Y(_608_)
);

OAI21X1 _4208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_595_),
    .C(_608_),
    .Y(_609_)
);

NAND2X1 _4209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_609_),
    .B(_605_),
    .Y(\partials[15] [30])
);

OAI21X1 _4210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_607_),
    .B(_595_),
    .C(_604_),
    .Y(_610_)
);

NOR2X1 _4211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_577_),
    .B(_601_),
    .Y(_611_)
);

NAND2X1 _4212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_611_),
    .B(_610_),
    .Y(\partials[15] [31])
);

INVX4 _4213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .Y(_613_)
);

NOR2X1 _4214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_613_),
    .Y(_614_)
);

NAND2X1 _4215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[1]),
    .Y(_615_)
);

INVX2 _4216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .Y(_616_)
);

NAND2X1 _4217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_616_),
    .B(_614_),
    .Y(_617_)
);

INVX2 _4218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .Y(_618_)
);

NOR2X1 _4219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_616_),
    .B(_614_),
    .Y(_619_)
);

NOR2X1 _4220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_619_),
    .B(_618_),
    .Y(\partials[7] [1])
);

NAND2X1 _4221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[2]),
    .Y(_620_)
);

NAND2X1 _4222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[2]),
    .Y(_622_)
);

INVX2 _4223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .Y(_623_)
);

NAND2X1 _4224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[2]),
    .Y(_624_)
);

OAI21X1 _4225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_613_),
    .C(_624_),
    .Y(_625_)
);

OAI21X1 _4226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_622_),
    .C(_625_),
    .Y(_626_)
);

OR2X2 _4227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_626_),
    .B(_620_),
    .Y(_627_)
);

INVX4 _4228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .Y(_628_)
);

OAI21X1 _4229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_628_),
    .C(_626_),
    .Y(_629_)
);

NAND2X1 _4230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_629_),
    .B(_627_),
    .Y(_630_)
);

XNOR2X1 _4231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_630_),
    .B(_618_),
    .Y(\partials[7] [2])
);

NOR2X1 _4232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_617_),
    .B(_630_),
    .Y(_631_)
);

INVX1 _4233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .Y(_632_)
);

NOR2X1 _4234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_628_),
    .Y(_633_)
);

INVX2 _4235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .Y(_634_)
);

OAI21X1 _4236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_615_),
    .B(_622_),
    .C(_627_),
    .Y(_635_)
);

INVX4 _4237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .Y(_636_)
);

NOR2X1 _4238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_636_),
    .Y(_637_)
);

NAND2X1 _4239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg[3]),
    .Y(_638_)
);

INVX1 _4240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .Y(_639_)
);

OAI21X1 _4241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_639_),
    .C(_622_),
    .Y(_640_)
);

OAI21X1 _4242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_638_),
    .C(_640_),
    .Y(_642_)
);

XNOR2X1 _4243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_637_),
    .Y(_643_)
);

NAND2X1 _4244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_635_),
    .Y(_644_)
);

INVX1 _4245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_622_),
    .Y(_645_)
);

NOR2X1 _4246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_620_),
    .B(_626_),
    .Y(_646_)
);

AOI21X1 _4247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_616_),
    .B(_645_),
    .C(_646_),
    .Y(_647_)
);

INVX1 _4248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .Y(_648_)
);

XNOR2X1 _4249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_642_),
    .B(_648_),
    .Y(_649_)
);

NAND2X1 _4250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_647_),
    .Y(_650_)
);

NAND3X1 _4251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_634_),
    .B(_650_),
    .C(_644_),
    .Y(_651_)
);

NOR2X1 _4252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_649_),
    .B(_647_),
    .Y(_653_)
);

NOR2X1 _4253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_643_),
    .B(_635_),
    .Y(_654_)
);

OAI21X1 _4254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_653_),
    .C(_633_),
    .Y(_655_)
);

AOI21X1 _4255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_651_),
    .B(_655_),
    .C(_632_),
    .Y(_656_)
);

NAND3X1 _4256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_650_),
    .C(_644_),
    .Y(_657_)
);

OAI21X1 _4257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_653_),
    .C(_634_),
    .Y(_658_)
);

AOI21X1 _4258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_657_),
    .B(_658_),
    .C(_631_),
    .Y(_659_)
);

NOR2X1 _4259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_656_),
    .B(_659_),
    .Y(\partials[7] [3])
);

NAND3X1 _4260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_631_),
    .B(_657_),
    .C(_658_),
    .Y(_660_)
);

OAI21X1 _4261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_654_),
    .B(_634_),
    .C(_644_),
    .Y(_661_)
);

NAND2X1 _4262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg[3]),
    .Y(_663_)
);

NOR2X1 _4263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_634_),
    .Y(_664_)
);

AOI22X1 _4264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg[3]),
    .C(breg[2]),
    .D(areg[2]),
    .Y(_665_)
);

OR2X2 _4265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_665_),
    .Y(_666_)
);

NOR2X1 _4266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_624_),
    .B(_638_),
    .Y(_667_)
);

AOI21X1 _4267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_637_),
    .B(_640_),
    .C(_667_),
    .Y(_668_)
);

NAND2X1 _4268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_4_bF$buf3),
    .Y(_669_)
);

INVX2 _4269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .Y(_670_)
);

NAND2X1 _4270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[4]),
    .Y(_671_)
);

OR2X2 _4271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_671_),
    .Y(_672_)
);

INVX2 _4272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .Y(_674_)
);

OAI21X1 _4273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_674_),
    .C(_638_),
    .Y(_675_)
);

NAND3X1 _4274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_675_),
    .C(_672_),
    .Y(_676_)
);

NOR2X1 _4275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_671_),
    .Y(_677_)
);

AND2X2 _4276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_638_),
    .B(_671_),
    .Y(_678_)
);

OAI21X1 _4277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_677_),
    .C(_669_),
    .Y(_679_)
);

NAND2X1 _4278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_679_),
    .B(_676_),
    .Y(_680_)
);

NOR2X1 _4279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .B(_680_),
    .Y(_681_)
);

INVX1 _4280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_668_),
    .Y(_682_)
);

AOI21X1 _4281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_676_),
    .B(_679_),
    .C(_682_),
    .Y(_683_)
);

NOR3X1 _4282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_666_),
    .B(_683_),
    .C(_681_),
    .Y(_685_)
);

NOR2X1 _4283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_665_),
    .B(_664_),
    .Y(_686_)
);

NOR3X1 _4284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_669_),
    .B(_677_),
    .C(_678_),
    .Y(_687_)
);

AOI21X1 _4285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_675_),
    .B(_672_),
    .C(_670_),
    .Y(_688_)
);

NOR2X1 _4286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_688_),
    .B(_687_),
    .Y(_689_)
);

NAND2X1 _4287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_682_),
    .B(_689_),
    .Y(_690_)
);

OAI21X1 _4288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_687_),
    .B(_688_),
    .C(_668_),
    .Y(_691_)
);

AOI21X1 _4289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_691_),
    .B(_690_),
    .C(_686_),
    .Y(_692_)
);

OAI21X1 _4290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .B(_692_),
    .C(_661_),
    .Y(_693_)
);

AOI21X1 _4291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_633_),
    .B(_650_),
    .C(_653_),
    .Y(_694_)
);

INVX1 _4292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .Y(_696_)
);

INVX1 _4293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_692_),
    .Y(_697_)
);

NAND3X1 _4294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_694_),
    .B(_697_),
    .C(_696_),
    .Y(_698_)
);

AOI21X1 _4295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_693_),
    .B(_698_),
    .C(_660_),
    .Y(_699_)
);

NAND3X1 _4296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_696_),
    .B(_697_),
    .C(_661_),
    .Y(_700_)
);

OAI21X1 _4297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .B(_692_),
    .C(_694_),
    .Y(_701_)
);

AOI21X1 _4298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_700_),
    .C(_656_),
    .Y(_702_)
);

NOR2X1 _4299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_702_),
    .Y(\partials[7] [4])
);

NAND3X1 _4300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_701_),
    .B(_656_),
    .C(_700_),
    .Y(_703_)
);

OAI21X1 _4301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_683_),
    .B(_666_),
    .C(_690_),
    .Y(_704_)
);

NOR2X1 _4302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_639_),
    .Y(_706_)
);

NAND2X1 _4303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg[5]),
    .Y(_707_)
);

XOR2X1 _4304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_707_),
    .Y(_708_)
);

XOR2X1 _4305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_706_),
    .Y(_709_)
);

OAI21X1 _4306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_678_),
    .B(_669_),
    .C(_672_),
    .Y(_710_)
);

NAND2X1 _4307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_4_bF$buf2),
    .Y(_711_)
);

INVX2 _4308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .Y(_712_)
);

AND2X2 _4309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg[4]),
    .Y(_713_)
);

AND2X2 _4310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg[5]),
    .Y(_714_)
);

NAND2X1 _4311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_713_),
    .B(_714_),
    .Y(_715_)
);

INVX2 _4312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .Y(_717_)
);

OAI22X1 _4313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_717_),
    .C(_613_),
    .D(_674_),
    .Y(_718_)
);

NAND3X1 _4314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_718_),
    .C(_715_),
    .Y(_719_)
);

NAND2X1 _4315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg[5]),
    .Y(_720_)
);

NOR2X1 _4316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_671_),
    .B(_720_),
    .Y(_721_)
);

NOR2X1 _4317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_713_),
    .B(_714_),
    .Y(_722_)
);

OAI21X1 _4318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_721_),
    .C(_711_),
    .Y(_723_)
);

NAND3X1 _4319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_710_),
    .B(_719_),
    .C(_723_),
    .Y(_724_)
);

AOI21X1 _4320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_670_),
    .B(_675_),
    .C(_677_),
    .Y(_725_)
);

NOR3X1 _4321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_711_),
    .B(_721_),
    .C(_722_),
    .Y(_726_)
);

AOI21X1 _4322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_718_),
    .B(_715_),
    .C(_712_),
    .Y(_728_)
);

OAI21X1 _4323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_728_),
    .C(_725_),
    .Y(_729_)
);

NAND3X1 _4324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_729_),
    .C(_709_),
    .Y(_730_)
);

XNOR2X1 _4325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_708_),
    .B(_706_),
    .Y(_731_)
);

NOR3X1 _4326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_728_),
    .B(_725_),
    .C(_726_),
    .Y(_732_)
);

AOI21X1 _4327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_719_),
    .B(_723_),
    .C(_710_),
    .Y(_733_)
);

OAI21X1 _4328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_732_),
    .B(_733_),
    .C(_731_),
    .Y(_734_)
);

NAND3X1 _4329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_734_),
    .C(_704_),
    .Y(_735_)
);

AOI21X1 _4330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_686_),
    .B(_691_),
    .C(_681_),
    .Y(_736_)
);

OAI21X1 _4331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_726_),
    .B(_728_),
    .C(_710_),
    .Y(_737_)
);

NAND3X1 _4332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_725_),
    .B(_719_),
    .C(_723_),
    .Y(_739_)
);

AOI21X1 _4333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_739_),
    .B(_737_),
    .C(_731_),
    .Y(_740_)
);

AOI21X1 _4334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_724_),
    .B(_729_),
    .C(_709_),
    .Y(_741_)
);

OAI21X1 _4335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_741_),
    .C(_736_),
    .Y(_742_)
);

NAND3X1 _4336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_742_),
    .C(_735_),
    .Y(_743_)
);

INVX2 _4337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .Y(_744_)
);

OAI21X1 _4338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_741_),
    .B(_740_),
    .C(_704_),
    .Y(_745_)
);

NAND3X1 _4339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_734_),
    .C(_736_),
    .Y(_746_)
);

NAND3X1 _4340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_745_),
    .C(_746_),
    .Y(_747_)
);

NAND3X1 _4341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_743_),
    .B(_700_),
    .C(_747_),
    .Y(_748_)
);

NOR3X1 _4342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_685_),
    .B(_692_),
    .C(_694_),
    .Y(_749_)
);

NAND3X1 _4343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_744_),
    .B(_742_),
    .C(_735_),
    .Y(_750_)
);

NAND3X1 _4344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_745_),
    .C(_746_),
    .Y(_751_)
);

NAND3X1 _4345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(_750_),
    .C(_751_),
    .Y(_752_)
);

AOI21X1 _4346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_752_),
    .B(_748_),
    .C(_703_),
    .Y(_753_)
);

NAND3X1 _4347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_749_),
    .B(_743_),
    .C(_747_),
    .Y(_754_)
);

NAND3X1 _4348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_700_),
    .C(_751_),
    .Y(_755_)
);

AOI21X1 _4349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_755_),
    .C(_699_),
    .Y(_756_)
);

NOR2X1 _4350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_756_),
    .Y(\partials[7] [5])
);

AOI21X1 _4351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_750_),
    .B(_751_),
    .C(_700_),
    .Y(_757_)
);

AOI21X1 _4352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_730_),
    .B(_734_),
    .C(_704_),
    .Y(_760_)
);

OAI21X1 _4353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_760_),
    .B(_744_),
    .C(_735_),
    .Y(_761_)
);

NOR2X1 _4354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_674_),
    .Y(_762_)
);

NAND2X1 _4355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_706_),
    .B(_708_),
    .Y(_763_)
);

OAI21X1 _4356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_663_),
    .B(_707_),
    .C(_763_),
    .Y(_764_)
);

XOR2X1 _4357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .B(_762_),
    .Y(_765_)
);

OAI21X1 _4358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_731_),
    .B(_733_),
    .C(_724_),
    .Y(_766_)
);

NAND2X1 _4359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .B(areg[3]),
    .Y(_767_)
);

INVX1 _4360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_767_),
    .Y(_768_)
);

NAND2X1 _4361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_6_bF$buf3),
    .Y(_769_)
);

NAND2X1 _4362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg[5]),
    .Y(_771_)
);

OR2X2 _4363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_771_),
    .Y(_772_)
);

INVX4 _4364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .Y(_773_)
);

OAI21X1 _4365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_140_),
    .B(_773_),
    .C(_771_),
    .Y(_774_)
);

NAND3X1 _4366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_768_),
    .B(_774_),
    .C(_772_),
    .Y(_775_)
);

NAND2X1 _4367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_6_bF$buf1),
    .Y(_776_)
);

NOR2X1 _4368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_707_),
    .B(_776_),
    .Y(_777_)
);

AND2X2 _4369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_769_),
    .B(_771_),
    .Y(_778_)
);

OAI21X1 _4370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_777_),
    .C(_767_),
    .Y(_779_)
);

AND2X2 _4371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_775_),
    .B(_779_),
    .Y(_780_)
);

OAI21X1 _4372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_722_),
    .B(_711_),
    .C(_715_),
    .Y(_782_)
);

NAND2X1 _4373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_4_bF$buf1),
    .Y(_783_)
);

INVX2 _4374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .Y(_784_)
);

NAND2X1 _4375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .B(breg[6]),
    .Y(_785_)
);

OR2X2 _4376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .B(_785_),
    .Y(_786_)
);

AOI22X1 _4377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[6]),
    .C(areg_1_bF$buf4),
    .D(breg[5]),
    .Y(_787_)
);

INVX2 _4378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_787_),
    .Y(_788_)
);

NAND3X1 _4379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_788_),
    .C(_786_),
    .Y(_789_)
);

NOR2X1 _4380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_720_),
    .B(_785_),
    .Y(_790_)
);

OAI21X1 _4381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_790_),
    .B(_787_),
    .C(_783_),
    .Y(_791_)
);

NAND3X1 _4382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_789_),
    .B(_791_),
    .C(_782_),
    .Y(_793_)
);

AOI21X1 _4383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_712_),
    .B(_718_),
    .C(_721_),
    .Y(_794_)
);

NOR3X1 _4384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_787_),
    .C(_790_),
    .Y(_795_)
);

AOI21X1 _4385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_788_),
    .B(_786_),
    .C(_784_),
    .Y(_796_)
);

OAI21X1 _4386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_795_),
    .C(_794_),
    .Y(_797_)
);

NAND3X1 _4387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_793_),
    .C(_797_),
    .Y(_798_)
);

NAND2X1 _4388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_779_),
    .B(_775_),
    .Y(_799_)
);

OAI21X1 _4389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_796_),
    .B(_795_),
    .C(_782_),
    .Y(_800_)
);

NAND3X1 _4390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_794_),
    .B(_791_),
    .C(_789_),
    .Y(_801_)
);

NAND3X1 _4391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_799_),
    .B(_801_),
    .C(_800_),
    .Y(_802_)
);

NAND3X1 _4392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_802_),
    .C(_766_),
    .Y(_804_)
);

AOI21X1 _4393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_729_),
    .B(_709_),
    .C(_732_),
    .Y(_805_)
);

AOI21X1 _4394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_801_),
    .B(_800_),
    .C(_799_),
    .Y(_806_)
);

AOI21X1 _4395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_793_),
    .B(_797_),
    .C(_780_),
    .Y(_807_)
);

OAI21X1 _4396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_807_),
    .B(_806_),
    .C(_805_),
    .Y(_808_)
);

NAND3X1 _4397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_808_),
    .C(_804_),
    .Y(_809_)
);

XNOR2X1 _4398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_764_),
    .B(_762_),
    .Y(_810_)
);

NOR3X1 _4399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_806_),
    .B(_807_),
    .C(_805_),
    .Y(_811_)
);

AOI21X1 _4400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_802_),
    .C(_766_),
    .Y(_812_)
);

OAI21X1 _4401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_811_),
    .B(_812_),
    .C(_810_),
    .Y(_813_)
);

NAND3X1 _4402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_813_),
    .C(_761_),
    .Y(_815_)
);

NOR3X1 _4403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_740_),
    .B(_741_),
    .C(_736_),
    .Y(_816_)
);

AOI21X1 _4404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_664_),
    .B(_742_),
    .C(_816_),
    .Y(_817_)
);

OAI21X1 _4405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_807_),
    .B(_806_),
    .C(_766_),
    .Y(_818_)
);

NAND3X1 _4406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_798_),
    .B(_802_),
    .C(_805_),
    .Y(_819_)
);

AOI21X1 _4407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_818_),
    .B(_819_),
    .C(_810_),
    .Y(_820_)
);

AOI21X1 _4408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_808_),
    .B(_804_),
    .C(_765_),
    .Y(_821_)
);

OAI21X1 _4409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(_821_),
    .C(_817_),
    .Y(_822_)
);

NAND3X1 _4410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_815_),
    .B(_822_),
    .C(_757_),
    .Y(_823_)
);

OAI21X1 _4411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_820_),
    .B(_821_),
    .C(_761_),
    .Y(_824_)
);

NAND3X1 _4412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_809_),
    .B(_813_),
    .C(_817_),
    .Y(_826_)
);

NAND3X1 _4413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_754_),
    .B(_824_),
    .C(_826_),
    .Y(_827_)
);

NAND2X1 _4414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_823_),
    .B(_827_),
    .Y(_828_)
);

XNOR2X1 _4415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_828_),
    .B(_753_),
    .Y(\partials[7] [6])
);

NAND3X1 _4416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_699_),
    .B(_754_),
    .C(_755_),
    .Y(_829_)
);

AOI21X1 _4417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_815_),
    .B(_822_),
    .C(_757_),
    .Y(_830_)
);

OAI21X1 _4418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_830_),
    .B(_829_),
    .C(_823_),
    .Y(_831_)
);

NAND2X1 _4419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_762_),
    .B(_764_),
    .Y(_832_)
);

OAI21X1 _4420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_812_),
    .B(_810_),
    .C(_804_),
    .Y(_833_)
);

NOR2X1 _4421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_717_),
    .Y(_834_)
);

INVX1 _4422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_834_),
    .Y(_836_)
);

NOR2X1 _4423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_674_),
    .Y(_837_)
);

INVX1 _4424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_837_),
    .Y(_838_)
);

OAI21X1 _4425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_778_),
    .B(_767_),
    .C(_772_),
    .Y(_839_)
);

AND2X2 _4426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_838_),
    .Y(_840_)
);

NOR2X1 _4427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_838_),
    .B(_839_),
    .Y(_841_)
);

OAI21X1 _4428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_840_),
    .B(_841_),
    .C(_836_),
    .Y(_842_)
);

AND2X2 _4429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_839_),
    .B(_837_),
    .Y(_843_)
);

NOR2X1 _4430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_837_),
    .B(_839_),
    .Y(_844_)
);

OAI21X1 _4431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_844_),
    .C(_834_),
    .Y(_845_)
);

NAND2X1 _4432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_845_),
    .Y(_847_)
);

AOI21X1 _4433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_791_),
    .B(_789_),
    .C(_782_),
    .Y(_848_)
);

OAI21X1 _4434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_848_),
    .B(_799_),
    .C(_793_),
    .Y(_849_)
);

NAND2X1 _4435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[0]),
    .B(areg_7_bF$buf3),
    .Y(_850_)
);

INVX1 _4436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_850_),
    .Y(_851_)
);

NAND2X1 _4437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg[5]),
    .Y(_852_)
);

OR2X2 _4438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_776_),
    .Y(_853_)
);

OAI21X1 _4439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_623_),
    .B(_773_),
    .C(_852_),
    .Y(_854_)
);

NAND3X1 _4440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_851_),
    .B(_854_),
    .C(_853_),
    .Y(_855_)
);

NOR2X1 _4441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_776_),
    .Y(_856_)
);

AND2X2 _4442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_776_),
    .Y(_858_)
);

OAI21X1 _4443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_856_),
    .C(_850_),
    .Y(_859_)
);

AND2X2 _4444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_855_),
    .B(_859_),
    .Y(_860_)
);

OAI21X1 _4445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_783_),
    .B(_787_),
    .C(_786_),
    .Y(_861_)
);

NAND2X1 _4446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .B(areg_4_bF$buf0),
    .Y(_862_)
);

INVX2 _4447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .Y(_863_)
);

AND2X2 _4448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[6]),
    .Y(_864_)
);

AND2X2 _4449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[7]),
    .Y(_865_)
);

NAND2X1 _4450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_864_),
    .B(_865_),
    .Y(_866_)
);

AOI22X1 _4451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[7]),
    .C(areg_1_bF$buf2),
    .D(breg[6]),
    .Y(_867_)
);

INVX2 _4452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_867_),
    .Y(_869_)
);

NAND3X1 _4453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_869_),
    .C(_866_),
    .Y(_870_)
);

NAND2X1 _4454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg[6]),
    .Y(_871_)
);

NAND2X1 _4455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg[7]),
    .Y(_872_)
);

NOR2X1 _4456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_871_),
    .B(_872_),
    .Y(_873_)
);

OAI21X1 _4457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_873_),
    .B(_867_),
    .C(_862_),
    .Y(_874_)
);

NAND3X1 _4458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_861_),
    .C(_870_),
    .Y(_875_)
);

AOI21X1 _4459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_784_),
    .B(_788_),
    .C(_790_),
    .Y(_876_)
);

NAND3X1 _4460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .B(breg[7]),
    .C(_871_),
    .Y(_877_)
);

NAND3X1 _4461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg[6]),
    .C(_872_),
    .Y(_878_)
);

AOI21X1 _4462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_877_),
    .B(_878_),
    .C(_862_),
    .Y(_880_)
);

AOI21X1 _4463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_869_),
    .B(_866_),
    .C(_863_),
    .Y(_881_)
);

OAI21X1 _4464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_880_),
    .C(_876_),
    .Y(_882_)
);

NAND3X1 _4465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_882_),
    .C(_860_),
    .Y(_883_)
);

NAND2X1 _4466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_859_),
    .B(_855_),
    .Y(_884_)
);

OAI21X1 _4467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_881_),
    .B(_880_),
    .C(_861_),
    .Y(_885_)
);

NAND3X1 _4468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_876_),
    .C(_870_),
    .Y(_886_)
);

NAND3X1 _4469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_884_),
    .B(_886_),
    .C(_885_),
    .Y(_887_)
);

NAND3X1 _4470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_883_),
    .C(_849_),
    .Y(_888_)
);

NOR3X1 _4471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_795_),
    .B(_794_),
    .C(_796_),
    .Y(_889_)
);

AOI21X1 _4472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_780_),
    .B(_797_),
    .C(_889_),
    .Y(_891_)
);

AOI21X1 _4473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_886_),
    .B(_885_),
    .C(_884_),
    .Y(_892_)
);

AOI21X1 _4474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_875_),
    .B(_882_),
    .C(_860_),
    .Y(_893_)
);

OAI21X1 _4475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_893_),
    .C(_891_),
    .Y(_894_)
);

NAND3X1 _4476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_888_),
    .C(_894_),
    .Y(_895_)
);

AND2X2 _4477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_842_),
    .B(_845_),
    .Y(_896_)
);

OAI21X1 _4478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_893_),
    .C(_849_),
    .Y(_897_)
);

NAND3X1 _4479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_883_),
    .B(_887_),
    .C(_891_),
    .Y(_898_)
);

NAND3X1 _4480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_897_),
    .C(_898_),
    .Y(_899_)
);

NAND3X1 _4481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_899_),
    .C(_833_),
    .Y(_900_)
);

AOI21X1 _4482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_765_),
    .B(_808_),
    .C(_811_),
    .Y(_902_)
);

AOI21X1 _4483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_897_),
    .B(_898_),
    .C(_896_),
    .Y(_903_)
);

AOI21X1 _4484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_888_),
    .B(_894_),
    .C(_847_),
    .Y(_904_)
);

OAI21X1 _4485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_903_),
    .B(_904_),
    .C(_902_),
    .Y(_905_)
);

NAND3X1 _4486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .B(_900_),
    .C(_905_),
    .Y(_906_)
);

INVX2 _4487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_832_),
    .Y(_907_)
);

NOR3X1 _4488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_903_),
    .B(_904_),
    .C(_902_),
    .Y(_908_)
);

AOI21X1 _4489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_895_),
    .B(_899_),
    .C(_833_),
    .Y(_909_)
);

OAI21X1 _4490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_909_),
    .C(_907_),
    .Y(_910_)
);

NAND3X1 _4491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_815_),
    .B(_906_),
    .C(_910_),
    .Y(_911_)
);

INVX1 _4492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_815_),
    .Y(_913_)
);

NAND3X1 _4493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_900_),
    .C(_905_),
    .Y(_914_)
);

OAI21X1 _4494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_908_),
    .B(_909_),
    .C(_832_),
    .Y(_915_)
);

NAND3X1 _4495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_913_),
    .B(_914_),
    .C(_915_),
    .Y(_916_)
);

AOI21X1 _4496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_916_),
    .B(_911_),
    .C(_831_),
    .Y(_917_)
);

AOI21X1 _4497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_831_),
    .B(_911_),
    .C(_917_),
    .Y(\partials[7] [7])
);

AOI21X1 _4498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_907_),
    .B(_905_),
    .C(_908_),
    .Y(_918_)
);

NOR2X1 _4499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_841_),
    .B(_840_),
    .Y(_919_)
);

NOR2X1 _4500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_836_),
    .B(_919_),
    .Y(_920_)
);

NOR2X1 _4501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_843_),
    .B(_920_),
    .Y(_921_)
);

INVX2 _4502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_921_),
    .Y(_923_)
);

AOI21X1 _4503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_887_),
    .B(_883_),
    .C(_849_),
    .Y(_924_)
);

OAI21X1 _4504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_896_),
    .B(_924_),
    .C(_888_),
    .Y(_925_)
);

INVX2 _4505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .Y(_926_)
);

NOR2X1 _4506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_926_),
    .Y(_927_)
);

INVX1 _4507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_927_),
    .Y(_928_)
);

NOR2X1 _4508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_717_),
    .Y(_929_)
);

INVX1 _4509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_929_),
    .Y(_930_)
);

OAI21X1 _4510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_858_),
    .B(_850_),
    .C(_853_),
    .Y(_931_)
);

AND2X2 _4511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_930_),
    .Y(_932_)
);

NOR2X1 _4512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_930_),
    .B(_931_),
    .Y(_934_)
);

OAI21X1 _4513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_932_),
    .B(_934_),
    .C(_928_),
    .Y(_935_)
);

AND2X2 _4514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_931_),
    .B(_929_),
    .Y(_936_)
);

NOR2X1 _4515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_929_),
    .B(_931_),
    .Y(_937_)
);

OAI21X1 _4516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(_937_),
    .C(_927_),
    .Y(_938_)
);

NAND2X1 _4517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(_938_),
    .Y(_939_)
);

AOI21X1 _4518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_874_),
    .B(_870_),
    .C(_861_),
    .Y(_940_)
);

OAI21X1 _4519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_940_),
    .B(_884_),
    .C(_875_),
    .Y(_941_)
);

NAND2X1 _4520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[1]),
    .B(areg_7_bF$buf2),
    .Y(_942_)
);

INVX1 _4521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .Y(_943_)
);

NAND2X1 _4522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .B(areg_6_bF$buf0),
    .Y(_945_)
);

OR2X2 _4523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_945_),
    .Y(_946_)
);

AOI22X1 _4524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_6_bF$buf3),
    .C(breg[3]),
    .D(areg[5]),
    .Y(_947_)
);

INVX1 _4525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_947_),
    .Y(_948_)
);

NAND3X1 _4526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_943_),
    .B(_948_),
    .C(_946_),
    .Y(_949_)
);

NOR2X1 _4527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_852_),
    .B(_945_),
    .Y(_950_)
);

OAI21X1 _4528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_950_),
    .B(_947_),
    .C(_942_),
    .Y(_951_)
);

AND2X2 _4529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_949_),
    .B(_951_),
    .Y(_952_)
);

OAI21X1 _4530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_862_),
    .B(_867_),
    .C(_866_),
    .Y(_953_)
);

NAND2X1 _4531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .B(areg_4_bF$buf3),
    .Y(_954_)
);

INVX2 _4532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_954_),
    .Y(_956_)
);

AND2X2 _4533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[8]),
    .Y(_957_)
);

NAND2X1 _4534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_865_),
    .B(_957_),
    .Y(_958_)
);

AOI22X1 _4535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[8]),
    .C(areg_1_bF$buf4),
    .D(breg[7]),
    .Y(_959_)
);

INVX2 _4536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_959_),
    .Y(_960_)
);

NAND3X1 _4537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(_960_),
    .C(_958_),
    .Y(_961_)
);

NAND2X1 _4538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[7]),
    .Y(_962_)
);

NAND2X1 _4539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[8]),
    .Y(_963_)
);

NOR2X1 _4540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_962_),
    .B(_963_),
    .Y(_964_)
);

OAI21X1 _4541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_964_),
    .B(_959_),
    .C(_954_),
    .Y(_965_)
);

NAND3X1 _4542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_953_),
    .B(_965_),
    .C(_961_),
    .Y(_966_)
);

AOI21X1 _4543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_863_),
    .B(_869_),
    .C(_873_),
    .Y(_967_)
);

NAND3X1 _4544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg[8]),
    .C(_962_),
    .Y(_968_)
);

NAND3X1 _4545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg[7]),
    .C(_963_),
    .Y(_969_)
);

AOI21X1 _4546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_968_),
    .B(_969_),
    .C(_954_),
    .Y(_970_)
);

AOI21X1 _4547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_960_),
    .B(_958_),
    .C(_956_),
    .Y(_971_)
);

OAI21X1 _4548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_970_),
    .C(_967_),
    .Y(_972_)
);

NAND3X1 _4549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_966_),
    .B(_972_),
    .C(_952_),
    .Y(_973_)
);

NAND2X1 _4550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_951_),
    .B(_949_),
    .Y(_974_)
);

OAI21X1 _4551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_971_),
    .B(_970_),
    .C(_953_),
    .Y(_975_)
);

NAND3X1 _4552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_967_),
    .C(_961_),
    .Y(_977_)
);

NAND3X1 _4553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_974_),
    .B(_977_),
    .C(_975_),
    .Y(_978_)
);

NAND3X1 _4554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_941_),
    .B(_978_),
    .C(_973_),
    .Y(_979_)
);

NOR3X1 _4555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_876_),
    .B(_880_),
    .C(_881_),
    .Y(_980_)
);

AOI21X1 _4556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_882_),
    .B(_860_),
    .C(_980_),
    .Y(_981_)
);

AOI21X1 _4557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_977_),
    .B(_975_),
    .C(_974_),
    .Y(_982_)
);

AOI21X1 _4558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_966_),
    .B(_972_),
    .C(_952_),
    .Y(_983_)
);

OAI21X1 _4559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .B(_983_),
    .C(_981_),
    .Y(_984_)
);

NAND3X1 _4560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_939_),
    .B(_979_),
    .C(_984_),
    .Y(_985_)
);

AND2X2 _4561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_935_),
    .B(_938_),
    .Y(_986_)
);

OAI21X1 _4562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .B(_983_),
    .C(_941_),
    .Y(_989_)
);

NAND3X1 _4563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_978_),
    .B(_973_),
    .C(_981_),
    .Y(_990_)
);

NAND3X1 _4564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_990_),
    .B(_986_),
    .C(_989_),
    .Y(_991_)
);

NAND3X1 _4565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .B(_991_),
    .C(_925_),
    .Y(_992_)
);

NOR3X1 _4566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_892_),
    .B(_893_),
    .C(_891_),
    .Y(_993_)
);

AOI21X1 _4567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_847_),
    .B(_894_),
    .C(_993_),
    .Y(_994_)
);

AOI21X1 _4568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_990_),
    .B(_989_),
    .C(_986_),
    .Y(_995_)
);

AOI21X1 _4569_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_979_),
    .B(_984_),
    .C(_939_),
    .Y(_996_)
);

OAI21X1 _4570_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(_996_),
    .C(_994_),
    .Y(_997_)
);

NAND3X1 _4571_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_992_),
    .C(_997_),
    .Y(_998_)
);

NOR3X1 _4572_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(_996_),
    .C(_994_),
    .Y(_999_)
);

AOI21X1 _4573_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .B(_991_),
    .C(_925_),
    .Y(_1000_)
);

OAI21X1 _4574_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_999_),
    .B(_1000_),
    .C(_921_),
    .Y(_1001_)
);

AOI21X1 _4575_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_1001_),
    .C(_918_),
    .Y(_1002_)
);

OAI21X1 _4576_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_909_),
    .B(_832_),
    .C(_900_),
    .Y(_1003_)
);

OAI21X1 _4577_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_995_),
    .B(_996_),
    .C(_925_),
    .Y(_1004_)
);

NAND3X1 _4578_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_985_),
    .B(_991_),
    .C(_994_),
    .Y(_1005_)
);

AOI21X1 _4579_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1005_),
    .B(_1004_),
    .C(_921_),
    .Y(_1006_)
);

AOI21X1 _4580_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_992_),
    .B(_997_),
    .C(_923_),
    .Y(_1007_)
);

NOR3X1 _4581_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1006_),
    .B(_1003_),
    .C(_1007_),
    .Y(_1008_)
);

NOR2X1 _4582_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1002_),
    .B(_1008_),
    .Y(_1010_)
);

AOI21X1 _4583_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_824_),
    .B(_826_),
    .C(_754_),
    .Y(_1011_)
);

AOI21X1 _4584_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_753_),
    .B(_827_),
    .C(_1011_),
    .Y(_1012_)
);

AOI21X1 _4585_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_914_),
    .B(_915_),
    .C(_913_),
    .Y(_1013_)
);

OAI21X1 _4586_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1012_),
    .B(_1013_),
    .C(_916_),
    .Y(_1014_)
);

XNOR2X1 _4587_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1014_),
    .B(_1010_),
    .Y(\partials[7] [8])
);

NAND3X1 _4588_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1003_),
    .B(_998_),
    .C(_1001_),
    .Y(_1015_)
);

AOI21X1 _4589_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_906_),
    .B(_910_),
    .C(_815_),
    .Y(_1016_)
);

AOI21X1 _4590_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_911_),
    .B(_831_),
    .C(_1016_),
    .Y(_1017_)
);

OAI21X1 _4591_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1017_),
    .B(_1010_),
    .C(_1015_),
    .Y(_1018_)
);

OAI21X1 _4592_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1000_),
    .B(_921_),
    .C(_992_),
    .Y(_1020_)
);

NOR2X1 _4593_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_934_),
    .B(_932_),
    .Y(_1021_)
);

NOR2X1 _4594_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_928_),
    .B(_1021_),
    .Y(_1022_)
);

NOR2X1 _4595_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_936_),
    .B(_1022_),
    .Y(_1023_)
);

INVX2 _4596_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1023_),
    .Y(_1024_)
);

AOI21X1 _4597_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_978_),
    .B(_973_),
    .C(_941_),
    .Y(_1025_)
);

OAI21X1 _4598_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_986_),
    .B(_1025_),
    .C(_979_),
    .Y(_1026_)
);

INVX1 _4599_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .Y(_1027_)
);

NOR2X1 _4600_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1027_),
    .Y(_1028_)
);

INVX1 _4601_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1028_),
    .Y(_1029_)
);

NOR2X1 _4602_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_926_),
    .Y(_1031_)
);

INVX1 _4603_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .Y(_1032_)
);

OAI21X1 _4604_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_942_),
    .B(_947_),
    .C(_946_),
    .Y(_1033_)
);

AND2X2 _4605_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(_1032_),
    .Y(_1034_)
);

NOR2X1 _4606_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1032_),
    .B(_1033_),
    .Y(_1035_)
);

OAI21X1 _4607_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1034_),
    .B(_1035_),
    .C(_1029_),
    .Y(_1036_)
);

AND2X2 _4608_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1033_),
    .B(_1031_),
    .Y(_1037_)
);

NOR2X1 _4609_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1031_),
    .B(_1033_),
    .Y(_1038_)
);

OAI21X1 _4610_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(_1038_),
    .C(_1028_),
    .Y(_1039_)
);

NAND2X1 _4611_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1039_),
    .Y(_1040_)
);

AOI21X1 _4612_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_965_),
    .B(_961_),
    .C(_953_),
    .Y(_1042_)
);

OAI21X1 _4613_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1042_),
    .B(_974_),
    .C(_966_),
    .Y(_1043_)
);

NAND2X1 _4614_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[2]),
    .B(areg_7_bF$buf1),
    .Y(_1044_)
);

INVX1 _4615_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1044_),
    .Y(_1045_)
);

NAND2X1 _4616_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .B(areg[5]),
    .Y(_1046_)
);

OR2X2 _4617_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_1046_),
    .Y(_1047_)
);

INVX4 _4618_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .Y(_1048_)
);

OAI21X1 _4619_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_674_),
    .B(_1048_),
    .C(_945_),
    .Y(_1049_)
);

NAND3X1 _4620_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1045_),
    .B(_1049_),
    .C(_1047_),
    .Y(_1050_)
);

NOR2X1 _4621_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_1046_),
    .Y(_1051_)
);

AND2X2 _4622_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_945_),
    .B(_1046_),
    .Y(_1053_)
);

OAI21X1 _4623_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1051_),
    .C(_1044_),
    .Y(_1054_)
);

AND2X2 _4624_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1050_),
    .B(_1054_),
    .Y(_1055_)
);

OAI21X1 _4625_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_954_),
    .B(_959_),
    .C(_958_),
    .Y(_1056_)
);

NAND2X1 _4626_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg[5]),
    .Y(_1057_)
);

INVX2 _4627_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1057_),
    .Y(_1058_)
);

AND2X2 _4628_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg[8]),
    .Y(_1059_)
);

AND2X2 _4629_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .B(breg[9]),
    .Y(_1060_)
);

NAND2X1 _4630_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1059_),
    .B(_1060_),
    .Y(_1061_)
);

INVX2 _4631_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[9]),
    .Y(_1062_)
);

NAND2X1 _4632_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg[8]),
    .Y(_1064_)
);

OAI21X1 _4633_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1062_),
    .C(_1064_),
    .Y(_1065_)
);

NAND3X1 _4634_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(_1065_),
    .C(_1061_),
    .Y(_1066_)
);

NAND2X1 _4635_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[9]),
    .Y(_1067_)
);

NOR2X1 _4636_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1067_),
    .Y(_1068_)
);

AND2X2 _4637_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1067_),
    .Y(_1069_)
);

OAI21X1 _4638_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .B(_1068_),
    .C(_1057_),
    .Y(_1070_)
);

NAND3X1 _4639_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1056_),
    .B(_1066_),
    .C(_1070_),
    .Y(_1071_)
);

AOI21X1 _4640_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_956_),
    .B(_960_),
    .C(_964_),
    .Y(_1072_)
);

NAND2X1 _4641_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1064_),
    .B(_1060_),
    .Y(_1073_)
);

NAND2X1 _4642_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1067_),
    .B(_1059_),
    .Y(_1075_)
);

AOI21X1 _4643_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1073_),
    .B(_1075_),
    .C(_1057_),
    .Y(_1076_)
);

AOI21X1 _4644_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1065_),
    .B(_1061_),
    .C(_1058_),
    .Y(_1077_)
);

OAI21X1 _4645_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1077_),
    .B(_1076_),
    .C(_1072_),
    .Y(_1078_)
);

NAND3X1 _4646_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1071_),
    .B(_1078_),
    .C(_1055_),
    .Y(_1079_)
);

NAND2X1 _4647_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1054_),
    .B(_1050_),
    .Y(_1080_)
);

OAI21X1 _4648_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1077_),
    .B(_1076_),
    .C(_1056_),
    .Y(_1081_)
);

NAND3X1 _4649_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1072_),
    .B(_1066_),
    .C(_1070_),
    .Y(_1082_)
);

NAND3X1 _4650_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1080_),
    .B(_1082_),
    .C(_1081_),
    .Y(_1083_)
);

NAND3X1 _4651_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1043_),
    .B(_1083_),
    .C(_1079_),
    .Y(_1084_)
);

NOR3X1 _4652_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_967_),
    .B(_970_),
    .C(_971_),
    .Y(_1086_)
);

AOI21X1 _4653_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_952_),
    .B(_972_),
    .C(_1086_),
    .Y(_1087_)
);

AOI21X1 _4654_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1082_),
    .B(_1081_),
    .C(_1080_),
    .Y(_1088_)
);

AOI21X1 _4655_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1071_),
    .B(_1078_),
    .C(_1055_),
    .Y(_1089_)
);

OAI21X1 _4656_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_1089_),
    .C(_1087_),
    .Y(_1090_)
);

NAND3X1 _4657_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_1084_),
    .C(_1090_),
    .Y(_1091_)
);

AND2X2 _4658_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1036_),
    .B(_1039_),
    .Y(_1092_)
);

OAI21X1 _4659_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_1089_),
    .C(_1043_),
    .Y(_1093_)
);

NAND3X1 _4660_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_1079_),
    .C(_1087_),
    .Y(_1094_)
);

NAND3X1 _4661_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1092_),
    .B(_1094_),
    .C(_1093_),
    .Y(_1095_)
);

NAND3X1 _4662_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1091_),
    .B(_1095_),
    .C(_1026_),
    .Y(_1097_)
);

NOR3X1 _4663_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_982_),
    .B(_983_),
    .C(_981_),
    .Y(_1098_)
);

AOI21X1 _4664_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_939_),
    .B(_984_),
    .C(_1098_),
    .Y(_1099_)
);

AOI21X1 _4665_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1094_),
    .B(_1093_),
    .C(_1092_),
    .Y(_1100_)
);

AOI21X1 _4666_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1084_),
    .B(_1090_),
    .C(_1040_),
    .Y(_1101_)
);

OAI21X1 _4667_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .B(_1101_),
    .C(_1099_),
    .Y(_1102_)
);

NAND3X1 _4668_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1097_),
    .C(_1102_),
    .Y(_1103_)
);

NOR3X1 _4669_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .B(_1101_),
    .C(_1099_),
    .Y(_1104_)
);

AOI21X1 _4670_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1091_),
    .B(_1095_),
    .C(_1026_),
    .Y(_1105_)
);

OAI21X1 _4671_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1104_),
    .B(_1105_),
    .C(_1023_),
    .Y(_1106_)
);

NAND3X1 _4672_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1020_),
    .B(_1103_),
    .C(_1106_),
    .Y(_1108_)
);

AOI21X1 _4673_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_923_),
    .B(_997_),
    .C(_999_),
    .Y(_1109_)
);

OAI21X1 _4674_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1100_),
    .B(_1101_),
    .C(_1026_),
    .Y(_1110_)
);

NAND3X1 _4675_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1091_),
    .B(_1095_),
    .C(_1099_),
    .Y(_1111_)
);

AOI21X1 _4676_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1111_),
    .B(_1110_),
    .C(_1023_),
    .Y(_1112_)
);

AOI21X1 _4677_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1097_),
    .B(_1102_),
    .C(_1024_),
    .Y(_1113_)
);

OAI21X1 _4678_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_1113_),
    .C(_1109_),
    .Y(_1114_)
);

NAND2X1 _4679_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1114_),
    .B(_1108_),
    .Y(_1115_)
);

XNOR2X1 _4680_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1018_),
    .B(_1115_),
    .Y(\partials[7] [9])
);

AOI21X1 _4681_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1103_),
    .B(_1106_),
    .C(_1020_),
    .Y(_1116_)
);

AOI21X1 _4682_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1015_),
    .B(_1108_),
    .C(_1116_),
    .Y(_1118_)
);

OAI21X1 _4683_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1006_),
    .B(_1007_),
    .C(_1003_),
    .Y(_1119_)
);

NAND3X1 _4684_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_998_),
    .B(_1001_),
    .C(_918_),
    .Y(_1120_)
);

OAI21X1 _4685_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_1113_),
    .C(_1020_),
    .Y(_1121_)
);

NAND3X1 _4686_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1109_),
    .B(_1103_),
    .C(_1106_),
    .Y(_1122_)
);

AOI22X1 _4687_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1122_),
    .B(_1121_),
    .C(_1119_),
    .D(_1120_),
    .Y(_1123_)
);

AOI21X1 _4688_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(_1014_),
    .C(_1118_),
    .Y(_1124_)
);

OAI21X1 _4689_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1105_),
    .B(_1023_),
    .C(_1097_),
    .Y(_1125_)
);

NOR2X1 _4690_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1035_),
    .B(_1034_),
    .Y(_1126_)
);

NOR2X1 _4691_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1029_),
    .B(_1126_),
    .Y(_1127_)
);

NOR2X1 _4692_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1037_),
    .B(_1127_),
    .Y(_1129_)
);

AOI21X1 _4693_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1083_),
    .B(_1079_),
    .C(_1043_),
    .Y(_1130_)
);

OAI21X1 _4694_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1130_),
    .B(_1092_),
    .C(_1084_),
    .Y(_1131_)
);

INVX1 _4695_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[8]),
    .Y(_1132_)
);

NOR2X1 _4696_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1132_),
    .Y(_1133_)
);

INVX1 _4697_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1133_),
    .Y(_1134_)
);

NOR2X1 _4698_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_1027_),
    .Y(_1135_)
);

INVX1 _4699_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .Y(_1136_)
);

OAI21X1 _4700_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1053_),
    .B(_1044_),
    .C(_1047_),
    .Y(_1137_)
);

AND2X2 _4701_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1136_),
    .Y(_1138_)
);

NOR2X1 _4702_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1136_),
    .B(_1137_),
    .Y(_1140_)
);

OAI21X1 _4703_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1138_),
    .B(_1140_),
    .C(_1134_),
    .Y(_1141_)
);

AND2X2 _4704_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1137_),
    .B(_1135_),
    .Y(_1142_)
);

NOR2X1 _4705_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1135_),
    .B(_1137_),
    .Y(_1143_)
);

OAI21X1 _4706_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1143_),
    .C(_1133_),
    .Y(_1144_)
);

AND2X2 _4707_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1144_),
    .Y(_1145_)
);

AOI21X1 _4708_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1066_),
    .B(_1070_),
    .C(_1056_),
    .Y(_1146_)
);

OAI21X1 _4709_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1146_),
    .B(_1080_),
    .C(_1071_),
    .Y(_1147_)
);

NAND2X1 _4710_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[3]),
    .B(areg_7_bF$buf0),
    .Y(_1148_)
);

NAND2X1 _4711_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .B(areg[5]),
    .Y(_1149_)
);

AOI21X1 _4712_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .B(areg_6_bF$buf2),
    .C(_1149_),
    .Y(_1151_)
);

NAND2X1 _4713_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .B(areg_6_bF$buf1),
    .Y(_1152_)
);

AOI21X1 _4714_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .B(areg[5]),
    .C(_1152_),
    .Y(_1153_)
);

OAI21X1 _4715_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1151_),
    .B(_1153_),
    .C(_1148_),
    .Y(_1154_)
);

INVX1 _4716_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1148_),
    .Y(_1155_)
);

NOR2X1 _4717_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1149_),
    .Y(_1156_)
);

AND2X2 _4718_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1152_),
    .B(_1149_),
    .Y(_1157_)
);

OAI21X1 _4719_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1157_),
    .B(_1156_),
    .C(_1155_),
    .Y(_1158_)
);

AND2X2 _4720_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1158_),
    .B(_1154_),
    .Y(_1159_)
);

OAI21X1 _4721_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1069_),
    .B(_1057_),
    .C(_1061_),
    .Y(_1160_)
);

NAND2X1 _4722_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg[6]),
    .Y(_1162_)
);

AND2X2 _4723_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[10]),
    .Y(_1163_)
);

OAI21X1 _4724_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_1062_),
    .C(_1163_),
    .Y(_1164_)
);

INVX4 _4725_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[10]),
    .Y(_1165_)
);

AND2X2 _4726_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg[9]),
    .Y(_1166_)
);

OAI21X1 _4727_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1165_),
    .C(_1166_),
    .Y(_1167_)
);

AOI21X1 _4728_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1164_),
    .B(_1167_),
    .C(_1162_),
    .Y(_1168_)
);

INVX2 _4729_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1162_),
    .Y(_1169_)
);

NAND2X1 _4730_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1163_),
    .Y(_1170_)
);

NAND2X1 _4731_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[9]),
    .Y(_1171_)
);

OAI21X1 _4732_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1165_),
    .C(_1171_),
    .Y(_1173_)
);

AOI21X1 _4733_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1173_),
    .B(_1170_),
    .C(_1169_),
    .Y(_1174_)
);

OAI21X1 _4734_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1174_),
    .C(_1160_),
    .Y(_1175_)
);

AOI21X1 _4735_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1058_),
    .B(_1065_),
    .C(_1068_),
    .Y(_1176_)
);

NAND3X1 _4736_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(_1173_),
    .C(_1170_),
    .Y(_1177_)
);

NAND2X1 _4737_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[10]),
    .Y(_1178_)
);

NOR2X1 _4738_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1171_),
    .B(_1178_),
    .Y(_1179_)
);

NOR2X1 _4739_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1166_),
    .B(_1163_),
    .Y(_1180_)
);

OAI21X1 _4740_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1180_),
    .B(_1179_),
    .C(_1162_),
    .Y(_1181_)
);

NAND3X1 _4741_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1176_),
    .B(_1177_),
    .C(_1181_),
    .Y(_1182_)
);

AOI21X1 _4742_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1175_),
    .B(_1182_),
    .C(_1159_),
    .Y(_1184_)
);

NAND2X1 _4743_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1154_),
    .B(_1158_),
    .Y(_1185_)
);

NAND3X1 _4744_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1177_),
    .B(_1160_),
    .C(_1181_),
    .Y(_1186_)
);

OAI21X1 _4745_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1168_),
    .B(_1174_),
    .C(_1176_),
    .Y(_1187_)
);

AOI21X1 _4746_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1187_),
    .B(_1186_),
    .C(_1185_),
    .Y(_1188_)
);

OAI21X1 _4747_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(_1188_),
    .C(_1147_),
    .Y(_1189_)
);

NOR3X1 _4748_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1076_),
    .B(_1072_),
    .C(_1077_),
    .Y(_1190_)
);

AOI21X1 _4749_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1055_),
    .B(_1078_),
    .C(_1190_),
    .Y(_1191_)
);

NAND3X1 _4750_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1187_),
    .C(_1186_),
    .Y(_1192_)
);

NAND3X1 _4751_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1159_),
    .B(_1175_),
    .C(_1182_),
    .Y(_1193_)
);

NAND3X1 _4752_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1193_),
    .B(_1192_),
    .C(_1191_),
    .Y(_1195_)
);

AOI21X1 _4753_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1195_),
    .B(_1189_),
    .C(_1145_),
    .Y(_1196_)
);

NAND2X1 _4754_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1141_),
    .B(_1144_),
    .Y(_1197_)
);

NAND3X1 _4755_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1147_),
    .B(_1192_),
    .C(_1193_),
    .Y(_1198_)
);

OAI21X1 _4756_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(_1188_),
    .C(_1191_),
    .Y(_1199_)
);

AOI21X1 _4757_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1198_),
    .B(_1199_),
    .C(_1197_),
    .Y(_1200_)
);

OAI21X1 _4758_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1200_),
    .C(_1131_),
    .Y(_1201_)
);

NOR3X1 _4759_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1088_),
    .B(_1089_),
    .C(_1087_),
    .Y(_1202_)
);

AOI21X1 _4760_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1040_),
    .B(_1090_),
    .C(_1202_),
    .Y(_1203_)
);

NAND3X1 _4761_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1198_),
    .B(_1197_),
    .C(_1199_),
    .Y(_1204_)
);

NAND3X1 _4762_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1195_),
    .B(_1145_),
    .C(_1189_),
    .Y(_1206_)
);

NAND3X1 _4763_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1204_),
    .B(_1206_),
    .C(_1203_),
    .Y(_1207_)
);

AOI21X1 _4764_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1207_),
    .B(_1201_),
    .C(_1129_),
    .Y(_1208_)
);

INVX2 _4765_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1129_),
    .Y(_1209_)
);

NAND3X1 _4766_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1131_),
    .B(_1204_),
    .C(_1206_),
    .Y(_1210_)
);

OAI21X1 _4767_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1200_),
    .C(_1203_),
    .Y(_1211_)
);

AOI21X1 _4768_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1210_),
    .B(_1211_),
    .C(_1209_),
    .Y(_1212_)
);

OAI21X1 _4769_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1212_),
    .C(_1125_),
    .Y(_1213_)
);

AOI21X1 _4770_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1024_),
    .B(_1102_),
    .C(_1104_),
    .Y(_1214_)
);

NAND3X1 _4771_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1209_),
    .B(_1210_),
    .C(_1211_),
    .Y(_1215_)
);

NOR3X1 _4772_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1196_),
    .B(_1200_),
    .C(_1203_),
    .Y(_1217_)
);

AOI21X1 _4773_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1204_),
    .B(_1206_),
    .C(_1131_),
    .Y(_1218_)
);

OAI21X1 _4774_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1217_),
    .B(_1218_),
    .C(_1129_),
    .Y(_1219_)
);

NAND3X1 _4775_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1214_),
    .B(_1215_),
    .C(_1219_),
    .Y(_1220_)
);

NAND2X1 _4776_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1213_),
    .B(_1220_),
    .Y(_1221_)
);

XNOR2X1 _4777_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1221_),
    .Y(\partials[7] [10])
);

NAND3X1 _4778_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1125_),
    .B(_1215_),
    .C(_1219_),
    .Y(_1222_)
);

INVX1 _4779_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1221_),
    .Y(_1223_)
);

OAI21X1 _4780_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1124_),
    .B(_1223_),
    .C(_1222_),
    .Y(_1224_)
);

OAI21X1 _4781_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1218_),
    .B(_1129_),
    .C(_1210_),
    .Y(_1225_)
);

NOR2X1 _4782_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1140_),
    .B(_1138_),
    .Y(_1227_)
);

NOR2X1 _4783_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1134_),
    .B(_1227_),
    .Y(_1228_)
);

NOR2X1 _4784_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1142_),
    .B(_1228_),
    .Y(_1229_)
);

INVX1 _4785_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1229_),
    .Y(_1230_)
);

AOI21X1 _4786_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1193_),
    .B(_1192_),
    .C(_1147_),
    .Y(_1231_)
);

OAI21X1 _4787_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1145_),
    .B(_1231_),
    .C(_1198_),
    .Y(_1232_)
);

NOR2X1 _4788_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1062_),
    .Y(_1233_)
);

INVX1 _4789_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1233_),
    .Y(_1234_)
);

NAND2X1 _4790_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[8]),
    .Y(_1235_)
);

NAND2X1 _4791_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .B(areg_6_bF$buf0),
    .Y(_1236_)
);

OAI22X1 _4792_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1046_),
    .B(_1236_),
    .C(_1157_),
    .D(_1148_),
    .Y(_1238_)
);

AND2X2 _4793_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .B(_1235_),
    .Y(_1239_)
);

NOR2X1 _4794_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1235_),
    .B(_1238_),
    .Y(_1240_)
);

OAI21X1 _4795_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .B(_1240_),
    .C(_1234_),
    .Y(_1241_)
);

INVX1 _4796_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1235_),
    .Y(_1242_)
);

AND2X2 _4797_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1238_),
    .B(_1242_),
    .Y(_1243_)
);

NOR2X1 _4798_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1242_),
    .B(_1238_),
    .Y(_1244_)
);

OAI21X1 _4799_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(_1244_),
    .C(_1233_),
    .Y(_1245_)
);

NAND2X1 _4800_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1245_),
    .Y(_1246_)
);

AOI21X1 _4801_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1177_),
    .B(_1181_),
    .C(_1160_),
    .Y(_1247_)
);

OAI21X1 _4802_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1247_),
    .B(_1159_),
    .C(_1186_),
    .Y(_1249_)
);

NAND2X1 _4803_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[4]),
    .B(areg_7_bF$buf3),
    .Y(_1250_)
);

NAND2X1 _4804_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_6_bF$buf3),
    .Y(_1251_)
);

OAI21X1 _4805_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_926_),
    .C(_1236_),
    .Y(_1252_)
);

OAI21X1 _4806_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1251_),
    .C(_1252_),
    .Y(_1253_)
);

XOR2X1 _4807_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .B(_1250_),
    .Y(_1254_)
);

OAI21X1 _4808_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1180_),
    .B(_1162_),
    .C(_1170_),
    .Y(_1255_)
);

NAND2X1 _4809_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg[7]),
    .Y(_1256_)
);

INVX2 _4810_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1256_),
    .Y(_1257_)
);

AND2X2 _4811_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg[10]),
    .Y(_1258_)
);

AND2X2 _4812_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg[11]),
    .Y(_1260_)
);

NAND2X1 _4813_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1258_),
    .B(_1260_),
    .Y(_1261_)
);

NAND2X1 _4814_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .B(breg[11]),
    .Y(_1262_)
);

OAI21X1 _4815_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_1165_),
    .C(_1262_),
    .Y(_1263_)
);

NAND3X1 _4816_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_1263_),
    .C(_1261_),
    .Y(_1264_)
);

NAND2X1 _4817_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg[11]),
    .Y(_1265_)
);

NOR2X1 _4818_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1178_),
    .B(_1265_),
    .Y(_1266_)
);

NOR2X1 _4819_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1258_),
    .B(_1260_),
    .Y(_1267_)
);

OAI21X1 _4820_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1267_),
    .B(_1266_),
    .C(_1256_),
    .Y(_1268_)
);

NAND3X1 _4821_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1264_),
    .B(_1255_),
    .C(_1268_),
    .Y(_1269_)
);

AOI21X1 _4822_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1169_),
    .B(_1173_),
    .C(_1179_),
    .Y(_1271_)
);

OAI21X1 _4823_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_1165_),
    .C(_1260_),
    .Y(_1272_)
);

INVX2 _4824_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[11]),
    .Y(_1273_)
);

OAI21X1 _4825_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1273_),
    .C(_1258_),
    .Y(_1274_)
);

AOI21X1 _4826_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1272_),
    .B(_1274_),
    .C(_1256_),
    .Y(_1275_)
);

AOI21X1 _4827_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1263_),
    .B(_1261_),
    .C(_1257_),
    .Y(_1276_)
);

OAI21X1 _4828_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(_1276_),
    .C(_1271_),
    .Y(_1277_)
);

NAND3X1 _4829_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(_1269_),
    .C(_1254_),
    .Y(_1278_)
);

XNOR2X1 _4830_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1253_),
    .B(_1250_),
    .Y(_1279_)
);

NOR3X1 _4831_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1276_),
    .B(_1271_),
    .C(_1275_),
    .Y(_1280_)
);

AOI21X1 _4832_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1264_),
    .B(_1268_),
    .C(_1255_),
    .Y(_1282_)
);

OAI21X1 _4833_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1280_),
    .B(_1282_),
    .C(_1279_),
    .Y(_1283_)
);

NAND3X1 _4834_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1249_),
    .B(_1278_),
    .C(_1283_),
    .Y(_1284_)
);

NOR3X1 _4835_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1174_),
    .B(_1176_),
    .C(_1168_),
    .Y(_1285_)
);

AOI21X1 _4836_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1185_),
    .B(_1187_),
    .C(_1285_),
    .Y(_1286_)
);

OAI21X1 _4837_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1275_),
    .B(_1276_),
    .C(_1255_),
    .Y(_1287_)
);

NAND3X1 _4838_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1271_),
    .B(_1264_),
    .C(_1268_),
    .Y(_1288_)
);

AOI21X1 _4839_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1287_),
    .B(_1288_),
    .C(_1279_),
    .Y(_1289_)
);

AOI21X1 _4840_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(_1269_),
    .C(_1254_),
    .Y(_1290_)
);

OAI21X1 _4841_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1289_),
    .C(_1286_),
    .Y(_1291_)
);

NAND3X1 _4842_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1246_),
    .B(_1291_),
    .C(_1284_),
    .Y(_1293_)
);

AND2X2 _4843_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1241_),
    .B(_1245_),
    .Y(_1294_)
);

OAI21X1 _4844_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1289_),
    .C(_1249_),
    .Y(_1295_)
);

NAND3X1 _4845_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1286_),
    .B(_1278_),
    .C(_1283_),
    .Y(_1296_)
);

NAND3X1 _4846_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1294_),
    .B(_1295_),
    .C(_1296_),
    .Y(_1297_)
);

NAND3X1 _4847_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1232_),
    .B(_1293_),
    .C(_1297_),
    .Y(_1298_)
);

NOR3X1 _4848_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1184_),
    .B(_1188_),
    .C(_1191_),
    .Y(_1299_)
);

AOI21X1 _4849_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1197_),
    .B(_1199_),
    .C(_1299_),
    .Y(_1300_)
);

AOI21X1 _4850_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1295_),
    .B(_1296_),
    .C(_1294_),
    .Y(_1301_)
);

AOI21X1 _4851_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1291_),
    .B(_1284_),
    .C(_1246_),
    .Y(_1302_)
);

OAI21X1 _4852_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1301_),
    .B(_1302_),
    .C(_1300_),
    .Y(_1304_)
);

NAND3X1 _4853_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1230_),
    .B(_1298_),
    .C(_1304_),
    .Y(_1305_)
);

NOR3X1 _4854_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1301_),
    .B(_1302_),
    .C(_1300_),
    .Y(_1306_)
);

AOI21X1 _4855_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1297_),
    .C(_1232_),
    .Y(_1307_)
);

OAI21X1 _4856_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1306_),
    .B(_1307_),
    .C(_1229_),
    .Y(_1308_)
);

NAND3X1 _4857_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1225_),
    .B(_1305_),
    .C(_1308_),
    .Y(_1309_)
);

AOI21X1 _4858_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1209_),
    .B(_1211_),
    .C(_1217_),
    .Y(_1310_)
);

OAI21X1 _4859_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1301_),
    .B(_1302_),
    .C(_1232_),
    .Y(_1311_)
);

NAND3X1 _4860_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1293_),
    .B(_1297_),
    .C(_1300_),
    .Y(_1312_)
);

AOI21X1 _4861_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1312_),
    .B(_1311_),
    .C(_1229_),
    .Y(_1313_)
);

AOI21X1 _4862_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1298_),
    .B(_1304_),
    .C(_1230_),
    .Y(_1315_)
);

OAI21X1 _4863_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1315_),
    .C(_1310_),
    .Y(_1316_)
);

NAND2X1 _4864_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1309_),
    .Y(_1317_)
);

XNOR2X1 _4865_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1224_),
    .B(_1317_),
    .Y(\partials[7] [11])
);

OAI21X1 _4866_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1315_),
    .C(_1225_),
    .Y(_1318_)
);

NAND3X1 _4867_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1310_),
    .B(_1305_),
    .C(_1308_),
    .Y(_1319_)
);

AOI22X1 _4868_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1220_),
    .B(_1213_),
    .C(_1319_),
    .D(_1318_),
    .Y(_1320_)
);

NAND3X1 _4869_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1123_),
    .B(_1320_),
    .C(_1014_),
    .Y(_1321_)
);

NAND2X1 _4870_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1222_),
    .B(_1309_),
    .Y(_1322_)
);

AOI22X1 _4871_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1322_),
    .C(_1320_),
    .D(_1118_),
    .Y(_1323_)
);

NAND2X1 _4872_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .B(_1323_),
    .Y(_1325_)
);

OAI21X1 _4873_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1307_),
    .B(_1229_),
    .C(_1298_),
    .Y(_1326_)
);

INVX2 _4874_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .Y(_1327_)
);

OAI21X1 _4875_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1239_),
    .B(_1240_),
    .C(_1233_),
    .Y(_1328_)
);

INVX1 _4876_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1328_),
    .Y(_1329_)
);

NOR2X1 _4877_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1243_),
    .B(_1329_),
    .Y(_1330_)
);

AOI21X1 _4878_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1278_),
    .B(_1283_),
    .C(_1249_),
    .Y(_1331_)
);

OAI21X1 _4879_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1331_),
    .B(_1294_),
    .C(_1284_),
    .Y(_1332_)
);

NOR2X1 _4880_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1165_),
    .Y(_1333_)
);

NAND2X1 _4881_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[9]),
    .Y(_1334_)
);

OAI22X1 _4882_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1149_),
    .B(_1251_),
    .C(_1253_),
    .D(_1250_),
    .Y(_1336_)
);

AND2X2 _4883_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1336_),
    .B(_1334_),
    .Y(_1337_)
);

NOR2X1 _4884_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .B(_1336_),
    .Y(_1338_)
);

OAI21X1 _4885_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(_1338_),
    .C(_1333_),
    .Y(_1339_)
);

INVX1 _4886_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1333_),
    .Y(_1340_)
);

INVX1 _4887_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1334_),
    .Y(_1341_)
);

AND2X2 _4888_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1336_),
    .B(_1341_),
    .Y(_1342_)
);

NOR2X1 _4889_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1341_),
    .B(_1336_),
    .Y(_1343_)
);

OAI21X1 _4890_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1343_),
    .C(_1340_),
    .Y(_1344_)
);

NAND2X1 _4891_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1339_),
    .B(_1344_),
    .Y(_1345_)
);

OAI21X1 _4892_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1279_),
    .B(_1282_),
    .C(_1269_),
    .Y(_1347_)
);

NAND2X1 _4893_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[5]),
    .B(areg_7_bF$buf2),
    .Y(_1348_)
);

NAND2X1 _4894_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[7]),
    .Y(_1349_)
);

NOR2X1 _4895_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(_1349_),
    .Y(_1350_)
);

AND2X2 _4896_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1251_),
    .B(_1349_),
    .Y(_1351_)
);

NOR2X1 _4897_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .B(_1351_),
    .Y(_1352_)
);

XOR2X1 _4898_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1348_),
    .Y(_1353_)
);

AOI21X1 _4899_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1257_),
    .B(_1263_),
    .C(_1266_),
    .Y(_1354_)
);

INVX2 _4900_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .Y(_1355_)
);

NAND2X1 _4901_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg[8]),
    .Y(_1356_)
);

NAND2X1 _4902_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg[12]),
    .Y(_1358_)
);

NOR2X1 _4903_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1262_),
    .B(_1358_),
    .Y(_1359_)
);

AOI22X1 _4904_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[12]),
    .C(areg_1_bF$buf4),
    .D(breg[11]),
    .Y(_1360_)
);

NOR3X1 _4905_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .B(_1360_),
    .C(_1359_),
    .Y(_1361_)
);

INVX2 _4906_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1356_),
    .Y(_1362_)
);

AND2X2 _4907_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[12]),
    .Y(_1363_)
);

NAND2X1 _4908_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1260_),
    .B(_1363_),
    .Y(_1364_)
);

INVX2 _4909_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .Y(_1365_)
);

AOI21X1 _4910_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1365_),
    .B(_1364_),
    .C(_1362_),
    .Y(_1366_)
);

OAI21X1 _4911_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1366_),
    .C(_1355_),
    .Y(_1367_)
);

NAND3X1 _4912_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1365_),
    .C(_1364_),
    .Y(_1369_)
);

OAI21X1 _4913_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1359_),
    .B(_1360_),
    .C(_1356_),
    .Y(_1370_)
);

NAND3X1 _4914_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1354_),
    .B(_1370_),
    .C(_1369_),
    .Y(_1371_)
);

AOI21X1 _4915_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1367_),
    .B(_1371_),
    .C(_1353_),
    .Y(_1372_)
);

XNOR2X1 _4916_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1352_),
    .B(_1348_),
    .Y(_1373_)
);

NAND3X1 _4917_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1370_),
    .C(_1355_),
    .Y(_1374_)
);

OAI21X1 _4918_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1366_),
    .B(_1361_),
    .C(_1354_),
    .Y(_1375_)
);

AOI21X1 _4919_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(_1374_),
    .C(_1373_),
    .Y(_1376_)
);

OAI21X1 _4920_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1376_),
    .B(_1372_),
    .C(_1347_),
    .Y(_1377_)
);

AOI21X1 _4921_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1277_),
    .B(_1254_),
    .C(_1280_),
    .Y(_1378_)
);

NAND3X1 _4922_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(_1374_),
    .C(_1373_),
    .Y(_1380_)
);

NOR3X1 _4923_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1361_),
    .B(_1354_),
    .C(_1366_),
    .Y(_1381_)
);

AOI21X1 _4924_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1369_),
    .B(_1370_),
    .C(_1355_),
    .Y(_1382_)
);

OAI21X1 _4925_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1382_),
    .B(_1381_),
    .C(_1353_),
    .Y(_1383_)
);

NAND3X1 _4926_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1378_),
    .B(_1383_),
    .C(_1380_),
    .Y(_1384_)
);

AOI21X1 _4927_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1384_),
    .B(_1377_),
    .C(_1345_),
    .Y(_1385_)
);

OAI21X1 _4928_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1337_),
    .B(_1338_),
    .C(_1340_),
    .Y(_1386_)
);

OAI21X1 _4929_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1343_),
    .C(_1333_),
    .Y(_1387_)
);

NAND2X1 _4930_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1386_),
    .B(_1387_),
    .Y(_1388_)
);

NAND3X1 _4931_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1347_),
    .B(_1383_),
    .C(_1380_),
    .Y(_1389_)
);

OAI21X1 _4932_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1376_),
    .B(_1372_),
    .C(_1378_),
    .Y(_1391_)
);

AOI21X1 _4933_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .B(_1391_),
    .C(_1388_),
    .Y(_1392_)
);

OAI21X1 _4934_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1392_),
    .C(_1332_),
    .Y(_1393_)
);

NOR3X1 _4935_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1290_),
    .B(_1289_),
    .C(_1286_),
    .Y(_1394_)
);

AOI21X1 _4936_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1246_),
    .B(_1291_),
    .C(_1394_),
    .Y(_1395_)
);

NAND3X1 _4937_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1389_),
    .B(_1391_),
    .C(_1388_),
    .Y(_1396_)
);

NOR3X1 _4938_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1372_),
    .B(_1378_),
    .C(_1376_),
    .Y(_1397_)
);

AOI21X1 _4939_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1383_),
    .B(_1380_),
    .C(_1347_),
    .Y(_1398_)
);

OAI21X1 _4940_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1397_),
    .B(_1398_),
    .C(_1345_),
    .Y(_1399_)
);

NAND3X1 _4941_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1395_),
    .B(_1396_),
    .C(_1399_),
    .Y(_1400_)
);

AOI21X1 _4942_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1393_),
    .B(_1400_),
    .C(_1330_),
    .Y(_1402_)
);

INVX2 _4943_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1330_),
    .Y(_1403_)
);

NAND3X1 _4944_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1332_),
    .B(_1396_),
    .C(_1399_),
    .Y(_1404_)
);

OAI21X1 _4945_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1392_),
    .C(_1395_),
    .Y(_1405_)
);

AOI21X1 _4946_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1405_),
    .B(_1404_),
    .C(_1403_),
    .Y(_1406_)
);

OAI21X1 _4947_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1402_),
    .B(_1406_),
    .C(_1327_),
    .Y(_1407_)
);

NAND3X1 _4948_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1405_),
    .C(_1404_),
    .Y(_1408_)
);

NOR3X1 _4949_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1385_),
    .B(_1395_),
    .C(_1392_),
    .Y(_1409_)
);

AOI21X1 _4950_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1396_),
    .B(_1399_),
    .C(_1332_),
    .Y(_1410_)
);

OAI21X1 _4951_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1409_),
    .B(_1410_),
    .C(_1330_),
    .Y(_1411_)
);

NAND3X1 _4952_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1326_),
    .B(_1408_),
    .C(_1411_),
    .Y(_1413_)
);

NAND2X1 _4953_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1407_),
    .B(_1413_),
    .Y(_1414_)
);

XNOR2X1 _4954_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1325_),
    .B(_1414_),
    .Y(\partials[7] [12])
);

NAND2X1 _4955_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1408_),
    .B(_1411_),
    .Y(_1415_)
);

AOI21X1 _4956_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1103_),
    .B(_1106_),
    .C(_1109_),
    .Y(_1416_)
);

NOR3X1 _4957_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_1020_),
    .C(_1113_),
    .Y(_1417_)
);

OAI22X1 _4958_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1008_),
    .B(_1002_),
    .C(_1416_),
    .D(_1417_),
    .Y(_1418_)
);

AOI21X1 _4959_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1215_),
    .B(_1219_),
    .C(_1214_),
    .Y(_1419_)
);

NOR3X1 _4960_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1125_),
    .C(_1212_),
    .Y(_1420_)
);

AOI21X1 _4961_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1305_),
    .B(_1308_),
    .C(_1310_),
    .Y(_1421_)
);

NOR3X1 _4962_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1225_),
    .C(_1315_),
    .Y(_1423_)
);

OAI22X1 _4963_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1419_),
    .B(_1420_),
    .C(_1423_),
    .D(_1421_),
    .Y(_1424_)
);

NOR3X1 _4964_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1418_),
    .B(_1017_),
    .C(_1424_),
    .Y(_1425_)
);

NOR3X1 _4965_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1006_),
    .B(_1007_),
    .C(_918_),
    .Y(_1426_)
);

NOR3X1 _4966_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1112_),
    .B(_1113_),
    .C(_1109_),
    .Y(_1427_)
);

OAI21X1 _4967_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1426_),
    .B(_1427_),
    .C(_1114_),
    .Y(_1428_)
);

NOR3X1 _4968_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1208_),
    .B(_1212_),
    .C(_1214_),
    .Y(_1429_)
);

NOR3X1 _4969_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1313_),
    .B(_1315_),
    .C(_1310_),
    .Y(_1430_)
);

AOI21X1 _4970_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1316_),
    .B(_1429_),
    .C(_1430_),
    .Y(_1431_)
);

OAI21X1 _4971_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1424_),
    .B(_1428_),
    .C(_1431_),
    .Y(_1432_)
);

AND2X2 _4972_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1413_),
    .B(_1407_),
    .Y(_1434_)
);

OAI21X1 _4973_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(_1432_),
    .C(_1434_),
    .Y(_1435_)
);

OAI21X1 _4974_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1327_),
    .B(_1415_),
    .C(_1435_),
    .Y(_1436_)
);

OAI21X1 _4975_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1410_),
    .B(_1330_),
    .C(_1404_),
    .Y(_1437_)
);

INVX1 _4976_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1339_),
    .Y(_1438_)
);

NOR2X1 _4977_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1342_),
    .B(_1438_),
    .Y(_1439_)
);

INVX2 _4978_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1439_),
    .Y(_1440_)
);

OAI21X1 _4979_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1345_),
    .B(_1398_),
    .C(_1389_),
    .Y(_1441_)
);

NAND2X1 _4980_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .B(breg[11]),
    .Y(_1442_)
);

NAND2X1 _4981_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[10]),
    .Y(_1443_)
);

INVX2 _4982_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1443_),
    .Y(_1445_)
);

INVX1 _4983_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1350_),
    .Y(_1446_)
);

OAI21X1 _4984_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1351_),
    .B(_1348_),
    .C(_1446_),
    .Y(_1447_)
);

XNOR2X1 _4985_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1447_),
    .B(_1445_),
    .Y(_1448_)
);

XOR2X1 _4986_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1442_),
    .Y(_1449_)
);

OAI21X1 _4987_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1353_),
    .B(_1382_),
    .C(_1374_),
    .Y(_1450_)
);

NAND2X1 _4988_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[6]),
    .B(areg_7_bF$buf1),
    .Y(_1451_)
);

NAND2X1 _4989_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg[7]),
    .Y(_1452_)
);

NAND2X1 _4990_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[8]),
    .Y(_1453_)
);

NOR2X1 _4991_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(_1453_),
    .Y(_1454_)
);

AND2X2 _4992_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1452_),
    .B(_1453_),
    .Y(_1456_)
);

NOR2X1 _4993_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1454_),
    .B(_1456_),
    .Y(_1457_)
);

XNOR2X1 _4994_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1457_),
    .B(_1451_),
    .Y(_1458_)
);

OAI21X1 _4995_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1360_),
    .B(_1356_),
    .C(_1364_),
    .Y(_1459_)
);

NAND2X1 _4996_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .B(breg[9]),
    .Y(_1460_)
);

INVX2 _4997_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .Y(_1461_)
);

AND2X2 _4998_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[13]),
    .Y(_1462_)
);

NAND2X1 _4999_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1462_),
    .Y(_1463_)
);

INVX2 _5000_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[13]),
    .Y(_1464_)
);

OAI21X1 _5001_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1464_),
    .C(_1358_),
    .Y(_1465_)
);

NAND3X1 _5002_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1461_),
    .B(_1465_),
    .C(_1463_),
    .Y(_1466_)
);

NAND2X1 _5003_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf1),
    .B(breg[13]),
    .Y(_1467_)
);

NOR2X1 _5004_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1467_),
    .Y(_1468_)
);

NOR2X1 _5005_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1363_),
    .B(_1462_),
    .Y(_1469_)
);

OAI21X1 _5006_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1468_),
    .C(_1460_),
    .Y(_1470_)
);

NAND3X1 _5007_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1459_),
    .B(_1466_),
    .C(_1470_),
    .Y(_1471_)
);

AOI21X1 _5008_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1362_),
    .B(_1365_),
    .C(_1359_),
    .Y(_1472_)
);

NOR3X1 _5009_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1460_),
    .B(_1468_),
    .C(_1469_),
    .Y(_1473_)
);

AOI21X1 _5010_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1465_),
    .B(_1463_),
    .C(_1461_),
    .Y(_1474_)
);

OAI21X1 _5011_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1474_),
    .C(_1472_),
    .Y(_1475_)
);

NAND3X1 _5012_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1471_),
    .B(_1475_),
    .C(_1458_),
    .Y(_1477_)
);

XOR2X1 _5013_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1457_),
    .B(_1451_),
    .Y(_1478_)
);

NOR3X1 _5014_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1472_),
    .B(_1474_),
    .C(_1473_),
    .Y(_1479_)
);

AOI21X1 _5015_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1466_),
    .B(_1470_),
    .C(_1459_),
    .Y(_1480_)
);

OAI21X1 _5016_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1479_),
    .B(_1480_),
    .C(_1478_),
    .Y(_1481_)
);

NAND3X1 _5017_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .B(_1481_),
    .C(_1450_),
    .Y(_1482_)
);

AOI21X1 _5018_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1375_),
    .B(_1373_),
    .C(_1381_),
    .Y(_1483_)
);

OAI21X1 _5019_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1473_),
    .B(_1474_),
    .C(_1459_),
    .Y(_1484_)
);

NAND3X1 _5020_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1472_),
    .B(_1466_),
    .C(_1470_),
    .Y(_1485_)
);

AOI21X1 _5021_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1485_),
    .B(_1484_),
    .C(_1478_),
    .Y(_1486_)
);

AOI21X1 _5022_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1471_),
    .B(_1475_),
    .C(_1458_),
    .Y(_1487_)
);

OAI21X1 _5023_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(_1487_),
    .C(_1483_),
    .Y(_1488_)
);

NAND3X1 _5024_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1449_),
    .B(_1488_),
    .C(_1482_),
    .Y(_1489_)
);

XNOR2X1 _5025_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1442_),
    .Y(_1490_)
);

OAI21X1 _5026_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(_1487_),
    .C(_1450_),
    .Y(_1491_)
);

NAND3X1 _5027_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .B(_1481_),
    .C(_1483_),
    .Y(_1492_)
);

NAND3X1 _5028_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1490_),
    .B(_1491_),
    .C(_1492_),
    .Y(_1493_)
);

NAND3X1 _5029_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1489_),
    .B(_1493_),
    .C(_1441_),
    .Y(_1494_)
);

AOI21X1 _5030_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1391_),
    .B(_1388_),
    .C(_1397_),
    .Y(_1495_)
);

AOI21X1 _5031_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1492_),
    .B(_1491_),
    .C(_1490_),
    .Y(_1496_)
);

AOI21X1 _5032_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1482_),
    .B(_1488_),
    .C(_1449_),
    .Y(_1498_)
);

OAI21X1 _5033_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1496_),
    .C(_1495_),
    .Y(_1499_)
);

NAND3X1 _5034_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1494_),
    .C(_1499_),
    .Y(_1500_)
);

NOR3X1 _5035_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1496_),
    .B(_1498_),
    .C(_1495_),
    .Y(_1501_)
);

AOI21X1 _5036_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1493_),
    .B(_1489_),
    .C(_1441_),
    .Y(_1502_)
);

OAI21X1 _5037_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1502_),
    .C(_1439_),
    .Y(_1503_)
);

NAND3X1 _5038_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1500_),
    .B(_1437_),
    .C(_1503_),
    .Y(_1504_)
);

AOI21X1 _5039_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1403_),
    .B(_1405_),
    .C(_1409_),
    .Y(_1505_)
);

OAI21X1 _5040_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1498_),
    .B(_1496_),
    .C(_1441_),
    .Y(_1506_)
);

NAND3X1 _5041_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1489_),
    .B(_1493_),
    .C(_1495_),
    .Y(_1507_)
);

AOI21X1 _5042_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1507_),
    .B(_1506_),
    .C(_1439_),
    .Y(_1510_)
);

AOI21X1 _5043_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1494_),
    .B(_1499_),
    .C(_1440_),
    .Y(_1511_)
);

OAI21X1 _5044_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1510_),
    .B(_1511_),
    .C(_1505_),
    .Y(_1512_)
);

NAND2X1 _5045_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1504_),
    .Y(_1513_)
);

XNOR2X1 _5046_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1436_),
    .B(_1513_),
    .Y(\partials[7] [13])
);

OAI21X1 _5047_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1415_),
    .B(_1327_),
    .C(_1504_),
    .Y(_1514_)
);

NAND2X1 _5048_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1512_),
    .B(_1514_),
    .Y(_1515_)
);

NOR2X1 _5049_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1414_),
    .Y(_1516_)
);

OAI21X1 _5050_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(_1432_),
    .C(_1516_),
    .Y(_1517_)
);

OAI21X1 _5051_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1502_),
    .B(_1439_),
    .C(_1494_),
    .Y(_1518_)
);

NAND2X1 _5052_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1445_),
    .B(_1447_),
    .Y(_1519_)
);

OAI21X1 _5053_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1448_),
    .B(_1442_),
    .C(_1519_),
    .Y(_1520_)
);

INVX2 _5054_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1520_),
    .Y(_1521_)
);

AOI21X1 _5055_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1477_),
    .B(_1481_),
    .C(_1450_),
    .Y(_1522_)
);

OAI21X1 _5056_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1522_),
    .B(_1490_),
    .C(_1482_),
    .Y(_1523_)
);

NAND2X1 _5057_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .B(breg[12]),
    .Y(_1524_)
);

NOR2X1 _5058_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_636_),
    .B(_1273_),
    .Y(_1525_)
);

NAND2X1 _5059_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg[8]),
    .Y(_1526_)
);

OAI22X1 _5060_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1349_),
    .B(_1526_),
    .C(_1456_),
    .D(_1451_),
    .Y(_1527_)
);

XNOR2X1 _5061_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1527_),
    .B(_1525_),
    .Y(_1528_)
);

XNOR2X1 _5062_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1524_),
    .Y(_1531_)
);

OAI21X1 _5063_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1478_),
    .B(_1480_),
    .C(_1471_),
    .Y(_1532_)
);

NAND2X1 _5064_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[7]),
    .B(areg_7_bF$buf0),
    .Y(_1533_)
);

NAND2X1 _5065_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg[9]),
    .Y(_1534_)
);

OAI21X1 _5066_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_1062_),
    .C(_1526_),
    .Y(_1535_)
);

OAI21X1 _5067_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .B(_1534_),
    .C(_1535_),
    .Y(_1536_)
);

XNOR2X1 _5068_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1533_),
    .Y(_1537_)
);

OAI21X1 _5069_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1469_),
    .B(_1460_),
    .C(_1463_),
    .Y(_1538_)
);

NAND2X1 _5070_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg[10]),
    .Y(_1539_)
);

NAND2X1 _5071_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf2),
    .B(breg[14]),
    .Y(_1540_)
);

NOR2X1 _5072_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1467_),
    .B(_1540_),
    .Y(_1542_)
);

AND2X2 _5073_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf1),
    .B(breg[13]),
    .Y(_1543_)
);

AND2X2 _5074_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf0),
    .B(breg[14]),
    .Y(_1544_)
);

NOR2X1 _5075_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1543_),
    .B(_1544_),
    .Y(_1545_)
);

NOR3X1 _5076_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .B(_1542_),
    .C(_1545_),
    .Y(_1546_)
);

INVX2 _5077_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1539_),
    .Y(_1547_)
);

NAND2X1 _5078_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1543_),
    .B(_1544_),
    .Y(_1548_)
);

NAND2X1 _5079_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf4),
    .B(breg[14]),
    .Y(_1549_)
);

OAI21X1 _5080_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_613_),
    .B(_1464_),
    .C(_1549_),
    .Y(_1550_)
);

AOI21X1 _5081_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1550_),
    .B(_1548_),
    .C(_1547_),
    .Y(_1551_)
);

OAI21X1 _5082_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1546_),
    .B(_1551_),
    .C(_1538_),
    .Y(_1553_)
);

AOI21X1 _5083_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1461_),
    .B(_1465_),
    .C(_1468_),
    .Y(_1554_)
);

NAND3X1 _5084_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1550_),
    .C(_1548_),
    .Y(_1555_)
);

OAI21X1 _5085_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1545_),
    .B(_1542_),
    .C(_1539_),
    .Y(_1556_)
);

NAND3X1 _5086_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1554_),
    .B(_1555_),
    .C(_1556_),
    .Y(_1557_)
);

AOI21X1 _5087_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1557_),
    .B(_1553_),
    .C(_1537_),
    .Y(_1558_)
);

XOR2X1 _5088_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1536_),
    .B(_1533_),
    .Y(_1559_)
);

NAND3X1 _5089_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1538_),
    .C(_1556_),
    .Y(_1560_)
);

OAI21X1 _5090_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1546_),
    .B(_1551_),
    .C(_1554_),
    .Y(_1561_)
);

AOI21X1 _5091_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1560_),
    .B(_1561_),
    .C(_1559_),
    .Y(_1562_)
);

OAI21X1 _5092_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .B(_1558_),
    .C(_1532_),
    .Y(_1564_)
);

AOI21X1 _5093_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1475_),
    .B(_1458_),
    .C(_1479_),
    .Y(_1565_)
);

NAND3X1 _5094_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1559_),
    .B(_1560_),
    .C(_1561_),
    .Y(_1566_)
);

NOR3X1 _5095_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1551_),
    .B(_1554_),
    .C(_1546_),
    .Y(_1567_)
);

AOI21X1 _5096_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1555_),
    .B(_1556_),
    .C(_1538_),
    .Y(_1568_)
);

OAI21X1 _5097_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1567_),
    .B(_1568_),
    .C(_1537_),
    .Y(_1569_)
);

NAND3X1 _5098_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .B(_1569_),
    .C(_1565_),
    .Y(_1570_)
);

AOI21X1 _5099_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1564_),
    .B(_1570_),
    .C(_1531_),
    .Y(_1571_)
);

XOR2X1 _5100_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1524_),
    .Y(_1572_)
);

NAND3X1 _5101_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .B(_1569_),
    .C(_1532_),
    .Y(_1573_)
);

OAI21X1 _5102_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .B(_1558_),
    .C(_1565_),
    .Y(_1575_)
);

AOI21X1 _5103_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1575_),
    .B(_1573_),
    .C(_1572_),
    .Y(_1576_)
);

OAI21X1 _5104_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(_1571_),
    .C(_1523_),
    .Y(_1577_)
);

NOR3X1 _5105_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1486_),
    .B(_1487_),
    .C(_1483_),
    .Y(_1578_)
);

AOI21X1 _5106_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1488_),
    .B(_1449_),
    .C(_1578_),
    .Y(_1579_)
);

NAND3X1 _5107_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1572_),
    .B(_1575_),
    .C(_1573_),
    .Y(_1580_)
);

NAND3X1 _5108_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1531_),
    .B(_1564_),
    .C(_1570_),
    .Y(_1581_)
);

NAND3X1 _5109_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1581_),
    .B(_1580_),
    .C(_1579_),
    .Y(_1582_)
);

AOI21X1 _5110_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1582_),
    .B(_1577_),
    .C(_1521_),
    .Y(_1583_)
);

NAND3X1 _5111_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1581_),
    .B(_1580_),
    .C(_1523_),
    .Y(_1584_)
);

OAI21X1 _5112_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(_1571_),
    .C(_1579_),
    .Y(_1586_)
);

AOI21X1 _5113_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1584_),
    .B(_1586_),
    .C(_1520_),
    .Y(_1587_)
);

OAI21X1 _5114_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1583_),
    .B(_1587_),
    .C(_1518_),
    .Y(_1588_)
);

AOI21X1 _5115_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1440_),
    .B(_1499_),
    .C(_1501_),
    .Y(_1589_)
);

NAND3X1 _5116_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1520_),
    .B(_1584_),
    .C(_1586_),
    .Y(_1590_)
);

NOR3X1 _5117_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1576_),
    .B(_1571_),
    .C(_1579_),
    .Y(_1591_)
);

AOI21X1 _5118_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1581_),
    .B(_1580_),
    .C(_1523_),
    .Y(_1592_)
);

OAI21X1 _5119_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1591_),
    .B(_1592_),
    .C(_1521_),
    .Y(_1593_)
);

NAND3X1 _5120_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(_1589_),
    .C(_1593_),
    .Y(_1594_)
);

AOI22X1 _5121_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1594_),
    .C(_1517_),
    .D(_1515_),
    .Y(_1595_)
);

NAND2X1 _5122_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1517_),
    .Y(_1597_)
);

NAND2X1 _5123_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1588_),
    .B(_1594_),
    .Y(_1598_)
);

NOR2X1 _5124_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1598_),
    .B(_1597_),
    .Y(_1599_)
);

NOR2X1 _5125_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1595_),
    .B(_1599_),
    .Y(\partials[7] [14])
);

NOR2X1 _5126_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1587_),
    .B(_1583_),
    .Y(_1600_)
);

AOI21X1 _5127_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1518_),
    .B(_1600_),
    .C(_1595_),
    .Y(_1601_)
);

OAI21X1 _5128_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1592_),
    .B(_1521_),
    .C(_1584_),
    .Y(_1602_)
);

NAND2X1 _5129_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .B(_1527_),
    .Y(_1603_)
);

OAI21X1 _5130_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1528_),
    .B(_1524_),
    .C(_1603_),
    .Y(_1604_)
);

INVX1 _5131_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .Y(_1605_)
);

AOI21X1 _5132_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1566_),
    .B(_1569_),
    .C(_1532_),
    .Y(_1607_)
);

OAI21X1 _5133_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1607_),
    .B(_1531_),
    .C(_1573_),
    .Y(_1608_)
);

NOR2X1 _5134_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1464_),
    .Y(_1609_)
);

NAND2X1 _5135_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[12]),
    .Y(_1610_)
);

OAI22X1 _5136_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1453_),
    .B(_1534_),
    .C(_1536_),
    .D(_1533_),
    .Y(_1611_)
);

AND2X2 _5137_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1611_),
    .B(_1610_),
    .Y(_1612_)
);

NOR2X1 _5138_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1610_),
    .B(_1611_),
    .Y(_1613_)
);

OAI21X1 _5139_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1613_),
    .C(_1609_),
    .Y(_1614_)
);

INVX1 _5140_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1609_),
    .Y(_1615_)
);

INVX1 _5141_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1610_),
    .Y(_1616_)
);

AND2X2 _5142_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1611_),
    .B(_1616_),
    .Y(_1618_)
);

NOR2X1 _5143_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1616_),
    .B(_1611_),
    .Y(_1619_)
);

OAI21X1 _5144_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1619_),
    .C(_1615_),
    .Y(_1620_)
);

NAND2X1 _5145_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1614_),
    .B(_1620_),
    .Y(_1621_)
);

OAI21X1 _5146_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1537_),
    .B(_1568_),
    .C(_1560_),
    .Y(_1622_)
);

NAND2X1 _5147_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg[8]),
    .Y(_1623_)
);

NAND2X1 _5148_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[9]),
    .Y(_1624_)
);

NAND2X1 _5149_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg[10]),
    .Y(_1625_)
);

OAI21X1 _5150_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_1165_),
    .C(_1534_),
    .Y(_1626_)
);

OAI21X1 _5151_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .B(_1625_),
    .C(_1626_),
    .Y(_1627_)
);

XNOR2X1 _5152_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1623_),
    .Y(_1629_)
);

OAI21X1 _5153_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1545_),
    .B(_1539_),
    .C(_1548_),
    .Y(_1630_)
);

NAND2X1 _5154_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg[11]),
    .Y(_1631_)
);

NAND3X1 _5155_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf3),
    .B(breg[15]),
    .C(_1540_),
    .Y(_1632_)
);

NAND2X1 _5156_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_0_bF$buf2),
    .B(breg[15]),
    .Y(_1633_)
);

NAND3X1 _5157_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf0),
    .B(breg[14]),
    .C(_1633_),
    .Y(_1634_)
);

AOI21X1 _5158_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1632_),
    .B(_1634_),
    .C(_1631_),
    .Y(_1635_)
);

INVX1 _5159_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1631_),
    .Y(_1636_)
);

AND2X2 _5160_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf4),
    .B(breg[15]),
    .Y(_1637_)
);

NAND2X1 _5161_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1544_),
    .B(_1637_),
    .Y(_1638_)
);

INVX2 _5162_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[15]),
    .Y(_1640_)
);

OAI21X1 _5163_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_129_),
    .B(_1640_),
    .C(_1540_),
    .Y(_1641_)
);

AOI21X1 _5164_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1641_),
    .B(_1638_),
    .C(_1636_),
    .Y(_1642_)
);

OAI21X1 _5165_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1635_),
    .C(_1630_),
    .Y(_1643_)
);

AOI21X1 _5166_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1547_),
    .B(_1550_),
    .C(_1542_),
    .Y(_1644_)
);

NAND3X1 _5167_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1636_),
    .B(_1641_),
    .C(_1638_),
    .Y(_1645_)
);

NAND3X1 _5168_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1631_),
    .B(_1632_),
    .C(_1634_),
    .Y(_1646_)
);

NAND3X1 _5169_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1644_),
    .B(_1646_),
    .C(_1645_),
    .Y(_1647_)
);

AOI21X1 _5170_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1647_),
    .C(_1629_),
    .Y(_1648_)
);

XOR2X1 _5171_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1627_),
    .B(_1623_),
    .Y(_1649_)
);

NAND3X1 _5172_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1645_),
    .B(_1646_),
    .C(_1630_),
    .Y(_1651_)
);

OAI21X1 _5173_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1642_),
    .B(_1635_),
    .C(_1644_),
    .Y(_1652_)
);

AOI21X1 _5174_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1652_),
    .B(_1651_),
    .C(_1649_),
    .Y(_1653_)
);

OAI21X1 _5175_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(_1648_),
    .C(_1622_),
    .Y(_1654_)
);

AOI21X1 _5176_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1561_),
    .B(_1559_),
    .C(_1567_),
    .Y(_1655_)
);

NAND3X1 _5177_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(_1652_),
    .C(_1649_),
    .Y(_1656_)
);

NAND3X1 _5178_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1643_),
    .B(_1647_),
    .C(_1629_),
    .Y(_1657_)
);

NAND3X1 _5179_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1657_),
    .B(_1656_),
    .C(_1655_),
    .Y(_1658_)
);

AOI21X1 _5180_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1654_),
    .B(_1658_),
    .C(_1621_),
    .Y(_1659_)
);

OAI21X1 _5181_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1612_),
    .B(_1613_),
    .C(_1615_),
    .Y(_1660_)
);

OAI21X1 _5182_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1619_),
    .C(_1609_),
    .Y(_1662_)
);

NAND2X1 _5183_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1660_),
    .B(_1662_),
    .Y(_1663_)
);

NAND3X1 _5184_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1656_),
    .B(_1657_),
    .C(_1622_),
    .Y(_1664_)
);

OAI21X1 _5185_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1653_),
    .B(_1648_),
    .C(_1655_),
    .Y(_1665_)
);

AOI21X1 _5186_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1664_),
    .B(_1665_),
    .C(_1663_),
    .Y(_1666_)
);

OAI21X1 _5187_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1666_),
    .C(_1608_),
    .Y(_1667_)
);

NOR3X1 _5188_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1562_),
    .B(_1558_),
    .C(_1565_),
    .Y(_1668_)
);

AOI21X1 _5189_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1575_),
    .B(_1572_),
    .C(_1668_),
    .Y(_1669_)
);

NAND3X1 _5190_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1664_),
    .B(_1665_),
    .C(_1663_),
    .Y(_1670_)
);

NAND3X1 _5191_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1654_),
    .B(_1658_),
    .C(_1621_),
    .Y(_1671_)
);

NAND3X1 _5192_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1670_),
    .B(_1671_),
    .C(_1669_),
    .Y(_1673_)
);

AOI21X1 _5193_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1673_),
    .B(_1667_),
    .C(_1605_),
    .Y(_1674_)
);

NAND3X1 _5194_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1608_),
    .B(_1670_),
    .C(_1671_),
    .Y(_1675_)
);

OAI21X1 _5195_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1659_),
    .B(_1666_),
    .C(_1669_),
    .Y(_1676_)
);

AOI21X1 _5196_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(_1676_),
    .C(_1604_),
    .Y(_1677_)
);

OAI21X1 _5197_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1674_),
    .B(_1677_),
    .C(_1602_),
    .Y(_1678_)
);

AOI21X1 _5198_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1520_),
    .B(_1586_),
    .C(_1591_),
    .Y(_1679_)
);

NAND3X1 _5199_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .B(_1675_),
    .C(_1676_),
    .Y(_1680_)
);

NAND3X1 _5200_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1605_),
    .B(_1673_),
    .C(_1667_),
    .Y(_1681_)
);

NAND3X1 _5201_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1680_),
    .B(_1681_),
    .C(_1679_),
    .Y(_1682_)
);

NAND2X1 _5202_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1682_),
    .B(_1678_),
    .Y(_1684_)
);

XNOR2X1 _5203_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1601_),
    .B(_1684_),
    .Y(\partials[7] [15])
);

AOI21X1 _5204_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1590_),
    .B(_1593_),
    .C(_1589_),
    .Y(_1685_)
);

NOR3X1 _5205_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1583_),
    .B(_1518_),
    .C(_1587_),
    .Y(_1686_)
);

AOI21X1 _5206_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1680_),
    .B(_1681_),
    .C(_1679_),
    .Y(_1687_)
);

NOR3X1 _5207_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(_1602_),
    .C(_1674_),
    .Y(_1688_)
);

OAI22X1 _5208_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1686_),
    .B(_1685_),
    .C(_1687_),
    .D(_1688_),
    .Y(_1689_)
);

NOR2X1 _5209_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1677_),
    .B(_1674_),
    .Y(_1690_)
);

OAI21X1 _5210_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1501_),
    .B(_1510_),
    .C(_1600_),
    .Y(_1691_)
);

INVX1 _5211_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1690_),
    .Y(_1692_)
);

OAI21X1 _5212_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1692_),
    .B(_1679_),
    .C(_1691_),
    .Y(_1694_)
);

OAI21X1 _5213_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1602_),
    .B(_1690_),
    .C(_1694_),
    .Y(_1695_)
);

OAI21X1 _5214_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1515_),
    .B(_1689_),
    .C(_1695_),
    .Y(_1696_)
);

AND2X2 _5215_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1504_),
    .B(_1512_),
    .Y(_1697_)
);

AOI22X1 _5216_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1678_),
    .B(_1682_),
    .C(_1594_),
    .D(_1588_),
    .Y(_1698_)
);

NAND3X1 _5217_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1697_),
    .B(_1434_),
    .C(_1698_),
    .Y(_1699_)
);

AOI21X1 _5218_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1321_),
    .B(_1323_),
    .C(_1699_),
    .Y(_1700_)
);

NOR2X1 _5219_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1700_),
    .B(_1696_),
    .Y(_1701_)
);

NAND2X1 _5220_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .B(_1680_),
    .Y(_1702_)
);

INVX1 _5221_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1614_),
    .Y(_1703_)
);

NOR2X1 _5222_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1618_),
    .B(_1703_),
    .Y(_1705_)
);

NAND2X1 _5223_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1664_),
    .B(_1670_),
    .Y(_1706_)
);

INVX1 _5224_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[14]),
    .Y(_1707_)
);

NOR2X1 _5225_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_628_),
    .B(_1707_),
    .Y(_1708_)
);

OAI22X1 _5226_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1624_),
    .B(_1625_),
    .C(_1627_),
    .D(_1623_),
    .Y(_1709_)
);

NOR2X1 _5227_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .B(_1709_),
    .Y(_1710_)
);

NAND2X1 _5228_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1708_),
    .B(_1709_),
    .Y(_1711_)
);

INVX2 _5229_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1711_),
    .Y(_1712_)
);

NOR2X1 _5230_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1710_),
    .B(_1712_),
    .Y(_1713_)
);

INVX2 _5231_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1713_),
    .Y(_1714_)
);

NAND2X1 _5232_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1651_),
    .B(_1656_),
    .Y(_1716_)
);

NAND2X1 _5233_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[13]),
    .Y(_1717_)
);

NAND2X1 _5234_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg[10]),
    .Y(_1718_)
);

NOR2X1 _5235_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .B(_1718_),
    .Y(_1719_)
);

AOI22X1 _5236_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf2),
    .B(breg[10]),
    .C(areg_7_bF$buf1),
    .D(breg[9]),
    .Y(_1720_)
);

OAI21X1 _5237_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1719_),
    .B(_1720_),
    .C(_1717_),
    .Y(_1721_)
);

NOR2X1 _5238_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1720_),
    .B(_1719_),
    .Y(_1722_)
);

NAND3X1 _5239_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[13]),
    .C(_1722_),
    .Y(_1723_)
);

NAND2X1 _5240_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1721_),
    .B(_1723_),
    .Y(_1724_)
);

NAND2X1 _5241_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_1_bF$buf3),
    .B(breg[15]),
    .Y(_1725_)
);

OAI21X1 _5242_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1549_),
    .B(_1725_),
    .C(_1645_),
    .Y(_1727_)
);

NOR2X1 _5243_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_1273_),
    .Y(_1728_)
);

INVX1 _5244_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1728_),
    .Y(_1729_)
);

NAND2X1 _5245_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg[15]),
    .Y(_1730_)
);

INVX2 _5246_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf2),
    .Y(_1731_)
);

INVX2 _5247_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(breg[12]),
    .Y(_1732_)
);

OAI21X1 _5248_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1731_),
    .B(_1732_),
    .C(_1725_),
    .Y(_1733_)
);

OAI21X1 _5249_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1358_),
    .B(_1730_),
    .C(_1733_),
    .Y(_1734_)
);

XNOR2X1 _5250_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1734_),
    .B(_1729_),
    .Y(_1735_)
);

NAND2X1 _5251_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_1735_),
    .Y(_1736_)
);

AOI21X1 _5252_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1544_),
    .B(_1637_),
    .C(_1635_),
    .Y(_1738_)
);

XNOR2X1 _5253_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1734_),
    .B(_1728_),
    .Y(_1739_)
);

NAND2X1 _5254_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1739_),
    .Y(_1740_)
);

AOI21X1 _5255_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1740_),
    .B(_1736_),
    .C(_1724_),
    .Y(_1741_)
);

INVX2 _5256_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1724_),
    .Y(_1742_)
);

NAND2X1 _5257_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_1739_),
    .Y(_1743_)
);

NAND2X1 _5258_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1735_),
    .Y(_1744_)
);

AOI21X1 _5259_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1743_),
    .B(_1744_),
    .C(_1742_),
    .Y(_1745_)
);

OAI21X1 _5260_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1745_),
    .B(_1741_),
    .C(_1716_),
    .Y(_1746_)
);

AND2X2 _5261_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1656_),
    .B(_1651_),
    .Y(_1747_)
);

NAND3X1 _5262_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1743_),
    .B(_1744_),
    .C(_1742_),
    .Y(_1749_)
);

NOR2X1 _5263_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1738_),
    .B(_1735_),
    .Y(_1750_)
);

NOR2X1 _5264_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1727_),
    .B(_1739_),
    .Y(_1751_)
);

OAI21X1 _5265_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1750_),
    .B(_1751_),
    .C(_1724_),
    .Y(_1752_)
);

NAND3X1 _5266_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1749_),
    .B(_1752_),
    .C(_1747_),
    .Y(_1753_)
);

AOI21X1 _5267_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1746_),
    .B(_1753_),
    .C(_1714_),
    .Y(_1754_)
);

NAND3X1 _5268_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1716_),
    .B(_1749_),
    .C(_1752_),
    .Y(_1755_)
);

OAI21X1 _5269_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1745_),
    .B(_1741_),
    .C(_1747_),
    .Y(_1756_)
);

AOI21X1 _5270_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1756_),
    .B(_1755_),
    .C(_1713_),
    .Y(_1757_)
);

OAI21X1 _5271_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(_1757_),
    .C(_1706_),
    .Y(_1758_)
);

NOR2X1 _5272_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1648_),
    .B(_1653_),
    .Y(_1760_)
);

AOI21X1 _5273_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1622_),
    .B(_1760_),
    .C(_1659_),
    .Y(_1761_)
);

NAND3X1 _5274_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1713_),
    .B(_1756_),
    .C(_1755_),
    .Y(_1762_)
);

NAND3X1 _5275_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1714_),
    .B(_1746_),
    .C(_1753_),
    .Y(_1763_)
);

NAND3X1 _5276_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1762_),
    .B(_1763_),
    .C(_1761_),
    .Y(_1764_)
);

AOI21X1 _5277_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1758_),
    .B(_1764_),
    .C(_1705_),
    .Y(_1765_)
);

INVX1 _5278_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .Y(_1766_)
);

NAND3X1 _5279_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1762_),
    .B(_1763_),
    .C(_1706_),
    .Y(_1767_)
);

OAI21X1 _5280_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1754_),
    .B(_1757_),
    .C(_1761_),
    .Y(_1768_)
);

AOI21X1 _5281_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1768_),
    .B(_1767_),
    .C(_1766_),
    .Y(_1769_)
);

OAI21X1 _5282_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1765_),
    .B(_1769_),
    .C(_1702_),
    .Y(_1771_)
);

INVX1 _5283_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1675_),
    .Y(_1772_)
);

AOI21X1 _5284_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1604_),
    .B(_1676_),
    .C(_1772_),
    .Y(_1773_)
);

NAND3X1 _5285_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1766_),
    .B(_1768_),
    .C(_1767_),
    .Y(_1774_)
);

NAND3X1 _5286_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1705_),
    .B(_1758_),
    .C(_1764_),
    .Y(_1775_)
);

NAND3X1 _5287_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1773_),
    .B(_1774_),
    .C(_1775_),
    .Y(_1776_)
);

NAND2X1 _5288_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1776_),
    .B(_1771_),
    .Y(_1777_)
);

XNOR2X1 _5289_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .B(_1777_),
    .Y(\partials[7] [16])
);

NAND2X1 _5290_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1774_),
    .B(_1775_),
    .Y(_1778_)
);

OR2X2 _5291_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1778_),
    .B(_1773_),
    .Y(_1779_)
);

AND2X2 _5292_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1771_),
    .B(_1776_),
    .Y(_1781_)
);

OAI21X1 _5293_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .B(_1781_),
    .C(_1779_),
    .Y(_1782_)
);

AND2X2 _5294_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1774_),
    .B(_1767_),
    .Y(_1783_)
);

NOR3X1 _5295_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1741_),
    .B(_1745_),
    .C(_1747_),
    .Y(_1784_)
);

AOI21X1 _5296_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1713_),
    .B(_1756_),
    .C(_1784_),
    .Y(_1785_)
);

OAI21X1 _5297_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1534_),
    .B(_1718_),
    .C(_1723_),
    .Y(_1786_)
);

AOI21X1 _5298_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1744_),
    .B(_1742_),
    .C(_1750_),
    .Y(_1787_)
);

NAND2X1 _5299_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .B(breg[15]),
    .Y(_1788_)
);

AOI22X1 _5300_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[14]),
    .C(areg_7_bF$buf0),
    .D(breg[10]),
    .Y(_1789_)
);

NAND2X1 _5301_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg[14]),
    .Y(_1790_)
);

NOR2X1 _5302_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1443_),
    .B(_1790_),
    .Y(_1792_)
);

OAI21X1 _5303_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1792_),
    .B(_1789_),
    .C(_1788_),
    .Y(_1793_)
);

NOR2X1 _5304_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1789_),
    .B(_1792_),
    .Y(_1794_)
);

NAND3X1 _5305_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[2]),
    .B(breg[15]),
    .C(_1794_),
    .Y(_1795_)
);

NAND2X1 _5306_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1793_),
    .B(_1795_),
    .Y(_1796_)
);

INVX2 _5307_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1796_),
    .Y(_1797_)
);

NAND2X1 _5308_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf1),
    .B(breg[12]),
    .Y(_1798_)
);

NOR2X1 _5309_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1725_),
    .B(_1798_),
    .Y(_1799_)
);

AOI21X1 _5310_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1728_),
    .B(_1733_),
    .C(_1799_),
    .Y(_1800_)
);

NOR2X1 _5311_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_1273_),
    .Y(_1801_)
);

INVX2 _5312_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1801_),
    .Y(_1803_)
);

NAND2X1 _5313_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[13]),
    .Y(_1804_)
);

NAND2X1 _5314_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf0),
    .B(breg[13]),
    .Y(_1805_)
);

OAI21X1 _5315_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1048_),
    .B(_1732_),
    .C(_1805_),
    .Y(_1806_)
);

OAI21X1 _5316_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .B(_1804_),
    .C(_1806_),
    .Y(_1807_)
);

XNOR2X1 _5317_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(_1803_),
    .Y(_1808_)
);

NAND2X1 _5318_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .B(_1808_),
    .Y(_1809_)
);

INVX1 _5319_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .Y(_1810_)
);

XNOR2X1 _5320_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1807_),
    .B(_1801_),
    .Y(_1811_)
);

NAND2X1 _5321_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .B(_1811_),
    .Y(_1812_)
);

AOI21X1 _5322_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1812_),
    .B(_1809_),
    .C(_1797_),
    .Y(_1814_)
);

NOR2X1 _5323_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1810_),
    .B(_1811_),
    .Y(_1815_)
);

NOR2X1 _5324_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1800_),
    .B(_1808_),
    .Y(_1816_)
);

NOR3X1 _5325_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_1796_),
    .C(_1816_),
    .Y(_1817_)
);

OAI21X1 _5326_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1817_),
    .B(_1814_),
    .C(_1787_),
    .Y(_1818_)
);

OAI21X1 _5327_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1751_),
    .B(_1724_),
    .C(_1743_),
    .Y(_1819_)
);

OAI21X1 _5328_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1816_),
    .B(_1815_),
    .C(_1796_),
    .Y(_1820_)
);

NAND3X1 _5329_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1812_),
    .C(_1797_),
    .Y(_1821_)
);

NAND3X1 _5330_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1821_),
    .B(_1819_),
    .C(_1820_),
    .Y(_1822_)
);

AOI21X1 _5331_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1822_),
    .B(_1818_),
    .C(_1786_),
    .Y(_1823_)
);

INVX2 _5332_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .Y(_1825_)
);

AOI21X1 _5333_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1821_),
    .B(_1820_),
    .C(_1819_),
    .Y(_1826_)
);

NOR3X1 _5334_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1787_),
    .B(_1814_),
    .C(_1817_),
    .Y(_1827_)
);

NOR3X1 _5335_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1825_),
    .B(_1826_),
    .C(_1827_),
    .Y(_1828_)
);

OAI21X1 _5336_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1828_),
    .B(_1823_),
    .C(_1785_),
    .Y(_1829_)
);

INVX1 _5337_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1756_),
    .Y(_1830_)
);

OAI21X1 _5338_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1830_),
    .B(_1714_),
    .C(_1755_),
    .Y(_1831_)
);

OAI21X1 _5339_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1827_),
    .B(_1826_),
    .C(_1825_),
    .Y(_1832_)
);

NAND3X1 _5340_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .B(_1822_),
    .C(_1818_),
    .Y(_1833_)
);

NAND3X1 _5341_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1832_),
    .B(_1833_),
    .C(_1831_),
    .Y(_1834_)
);

AOI21X1 _5342_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1834_),
    .B(_1829_),
    .C(_1712_),
    .Y(_1836_)
);

AOI21X1 _5343_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1833_),
    .B(_1832_),
    .C(_1831_),
    .Y(_1837_)
);

NOR3X1 _5344_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1785_),
    .B(_1823_),
    .C(_1828_),
    .Y(_1838_)
);

NOR3X1 _5345_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1711_),
    .B(_1837_),
    .C(_1838_),
    .Y(_1839_)
);

OAI21X1 _5346_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1839_),
    .B(_1836_),
    .C(_1783_),
    .Y(_1840_)
);

NAND2X1 _5347_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1767_),
    .B(_1774_),
    .Y(_1841_)
);

OAI21X1 _5348_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1838_),
    .B(_1837_),
    .C(_1711_),
    .Y(_1842_)
);

NAND3X1 _5349_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(_1834_),
    .C(_1829_),
    .Y(_1843_)
);

NAND3X1 _5350_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1842_),
    .B(_1843_),
    .C(_1841_),
    .Y(_1844_)
);

AND2X2 _5351_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .B(_1844_),
    .Y(_1845_)
);

XOR2X1 _5352_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1782_),
    .B(_1845_),
    .Y(\partials[7] [17])
);

NAND3X1 _5353_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1844_),
    .B(_1840_),
    .C(_1777_),
    .Y(_1847_)
);

OAI21X1 _5354_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1773_),
    .B(_1778_),
    .C(_1844_),
    .Y(_1848_)
);

NAND2X1 _5355_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1840_),
    .B(_1848_),
    .Y(_1849_)
);

OAI21X1 _5356_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .B(_1847_),
    .C(_1849_),
    .Y(_1850_)
);

AOI21X1 _5357_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1786_),
    .B(_1818_),
    .C(_1827_),
    .Y(_1851_)
);

OAI21X1 _5358_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1443_),
    .B(_1790_),
    .C(_1795_),
    .Y(_1852_)
);

AOI21X1 _5359_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1809_),
    .B(_1797_),
    .C(_1816_),
    .Y(_1853_)
);

INVX1 _5360_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1525_),
    .Y(_1854_)
);

NAND2X1 _5361_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf2),
    .B(breg[15]),
    .Y(_1855_)
);

NOR2X1 _5362_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .B(_1854_),
    .Y(_1857_)
);

AOI22X1 _5363_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[3]),
    .B(breg[15]),
    .C(areg_7_bF$buf1),
    .D(breg[11]),
    .Y(_1858_)
);

NOR2X1 _5364_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1858_),
    .B(_1857_),
    .Y(_1859_)
);

OAI22X1 _5365_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1798_),
    .B(_1804_),
    .C(_1807_),
    .D(_1803_),
    .Y(_1860_)
);

INVX1 _5366_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1860_),
    .Y(_1861_)
);

NAND2X1 _5367_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[14]),
    .Y(_1862_)
);

OAI21X1 _5368_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1731_),
    .B(_1707_),
    .C(_1804_),
    .Y(_1863_)
);

OAI21X1 _5369_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1805_),
    .B(_1862_),
    .C(_1863_),
    .Y(_1864_)
);

OAI21X1 _5370_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_1732_),
    .C(_1864_),
    .Y(_1865_)
);

NOR2X1 _5371_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_1732_),
    .Y(_1866_)
);

NAND2X1 _5372_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_4_bF$buf3),
    .B(breg[14]),
    .Y(_1868_)
);

OR2X2 _5373_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1804_),
    .B(_1868_),
    .Y(_1869_)
);

NAND3X1 _5374_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1866_),
    .B(_1863_),
    .C(_1869_),
    .Y(_1870_)
);

NAND2X1 _5375_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .B(_1865_),
    .Y(_1871_)
);

NAND2X1 _5376_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1871_),
    .B(_1861_),
    .Y(_1872_)
);

AND2X2 _5377_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1865_),
    .B(_1870_),
    .Y(_1873_)
);

NAND2X1 _5378_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1860_),
    .B(_1873_),
    .Y(_1874_)
);

AOI21X1 _5379_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1872_),
    .B(_1874_),
    .C(_1859_),
    .Y(_1875_)
);

INVX2 _5380_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1859_),
    .Y(_1876_)
);

NOR2X1 _5381_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1860_),
    .B(_1873_),
    .Y(_1877_)
);

NOR2X1 _5382_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1871_),
    .B(_1861_),
    .Y(_1879_)
);

NOR3X1 _5383_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1876_),
    .B(_1879_),
    .C(_1877_),
    .Y(_1880_)
);

OAI21X1 _5384_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1880_),
    .B(_1875_),
    .C(_1853_),
    .Y(_1881_)
);

OAI21X1 _5385_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1815_),
    .B(_1796_),
    .C(_1812_),
    .Y(_1882_)
);

OAI21X1 _5386_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1877_),
    .B(_1879_),
    .C(_1876_),
    .Y(_1883_)
);

NAND3X1 _5387_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1859_),
    .B(_1872_),
    .C(_1874_),
    .Y(_1884_)
);

NAND3X1 _5388_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1882_),
    .C(_1883_),
    .Y(_1885_)
);

AOI21X1 _5389_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1885_),
    .B(_1881_),
    .C(_1852_),
    .Y(_1886_)
);

INVX2 _5390_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .Y(_1887_)
);

AOI21X1 _5391_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1884_),
    .B(_1883_),
    .C(_1882_),
    .Y(_1888_)
);

NOR3X1 _5392_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1853_),
    .B(_1875_),
    .C(_1880_),
    .Y(_1890_)
);

NOR3X1 _5393_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1887_),
    .B(_1888_),
    .C(_1890_),
    .Y(_1891_)
);

OAI21X1 _5394_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1891_),
    .B(_1886_),
    .C(_1851_),
    .Y(_1892_)
);

OAI21X1 _5395_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1826_),
    .B(_1825_),
    .C(_1822_),
    .Y(_1893_)
);

OAI21X1 _5396_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1890_),
    .B(_1888_),
    .C(_1887_),
    .Y(_1894_)
);

NAND3X1 _5397_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_1885_),
    .C(_1881_),
    .Y(_1895_)
);

NAND3X1 _5398_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1893_),
    .B(_1895_),
    .C(_1894_),
    .Y(_1896_)
);

NAND2X1 _5399_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1896_),
    .B(_1892_),
    .Y(_1897_)
);

OAI21X1 _5400_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1839_),
    .B(_1838_),
    .C(_1897_),
    .Y(_1898_)
);

AOI21X1 _5401_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1712_),
    .B(_1829_),
    .C(_1838_),
    .Y(_1899_)
);

NAND3X1 _5402_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1892_),
    .B(_1896_),
    .C(_1899_),
    .Y(_1901_)
);

NAND2X1 _5403_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1898_),
    .Y(_1902_)
);

INVX2 _5404_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1902_),
    .Y(_1903_)
);

XNOR2X1 _5405_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1850_),
    .B(_1903_),
    .Y(\partials[7] [18])
);

NOR2X1 _5406_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1897_),
    .B(_1899_),
    .Y(_1904_)
);

INVX1 _5407_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1847_),
    .Y(_1905_)
);

OAI21X1 _5408_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1696_),
    .B(_1700_),
    .C(_1905_),
    .Y(_1906_)
);

AOI21X1 _5409_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1849_),
    .B(_1906_),
    .C(_1903_),
    .Y(_1907_)
);

OAI21X1 _5410_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1888_),
    .B(_1887_),
    .C(_1885_),
    .Y(_1908_)
);

INVX2 _5411_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1857_),
    .Y(_1909_)
);

OAI21X1 _5412_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1877_),
    .B(_1876_),
    .C(_1874_),
    .Y(_1911_)
);

INVX1 _5413_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf0),
    .Y(_1912_)
);

NOR2X1 _5414_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1912_),
    .B(_1732_),
    .Y(_1913_)
);

INVX1 _5415_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1913_),
    .Y(_1914_)
);

OAI21X1 _5416_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1805_),
    .B(_1862_),
    .C(_1870_),
    .Y(_1915_)
);

NAND2X1 _5417_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf1),
    .B(breg[13]),
    .Y(_1916_)
);

NAND2X1 _5418_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg[5]),
    .B(breg[15]),
    .Y(_1917_)
);

OAI21X1 _5419_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1731_),
    .B(_1640_),
    .C(_1862_),
    .Y(_1918_)
);

OAI21X1 _5420_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(_1917_),
    .C(_1918_),
    .Y(_1919_)
);

XOR2X1 _5421_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1916_),
    .Y(_1920_)
);

NOR2X1 _5422_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1915_),
    .B(_1920_),
    .Y(_1922_)
);

AND2X2 _5423_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1870_),
    .B(_1869_),
    .Y(_1923_)
);

XNOR2X1 _5424_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1919_),
    .B(_1916_),
    .Y(_1924_)
);

NOR2X1 _5425_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .B(_1924_),
    .Y(_1925_)
);

OAI21X1 _5426_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1922_),
    .B(_1925_),
    .C(_1914_),
    .Y(_1926_)
);

NAND2X1 _5427_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1923_),
    .B(_1924_),
    .Y(_1927_)
);

NAND2X1 _5428_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1915_),
    .B(_1920_),
    .Y(_1928_)
);

NAND3X1 _5429_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1913_),
    .B(_1927_),
    .C(_1928_),
    .Y(_1929_)
);

AOI21X1 _5430_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1929_),
    .B(_1926_),
    .C(_1911_),
    .Y(_1930_)
);

AOI21X1 _5431_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1859_),
    .B(_1872_),
    .C(_1879_),
    .Y(_1931_)
);

AOI21X1 _5432_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1927_),
    .B(_1928_),
    .C(_1913_),
    .Y(_1933_)
);

INVX2 _5433_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1929_),
    .Y(_1934_)
);

NOR3X1 _5434_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1931_),
    .B(_1933_),
    .C(_1934_),
    .Y(_1935_)
);

OAI21X1 _5435_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1935_),
    .B(_1930_),
    .C(_1909_),
    .Y(_1936_)
);

OAI21X1 _5436_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1934_),
    .B(_1933_),
    .C(_1931_),
    .Y(_1937_)
);

NAND3X1 _5437_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1926_),
    .B(_1929_),
    .C(_1911_),
    .Y(_1938_)
);

NAND3X1 _5438_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1857_),
    .B(_1938_),
    .C(_1937_),
    .Y(_1939_)
);

AOI21X1 _5439_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1939_),
    .B(_1936_),
    .C(_1908_),
    .Y(_1940_)
);

AOI21X1 _5440_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1852_),
    .B(_1881_),
    .C(_1890_),
    .Y(_1941_)
);

AOI21X1 _5441_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1938_),
    .B(_1937_),
    .C(_1857_),
    .Y(_1942_)
);

NOR3X1 _5442_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1909_),
    .B(_1930_),
    .C(_1935_),
    .Y(_1944_)
);

NOR3X1 _5443_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1942_),
    .B(_1941_),
    .C(_1944_),
    .Y(_1945_)
);

OAI21X1 _5444_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1945_),
    .B(_1940_),
    .C(_1896_),
    .Y(_1946_)
);

NOR3X1 _5445_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1851_),
    .B(_1886_),
    .C(_1891_),
    .Y(_1947_)
);

OAI21X1 _5446_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1944_),
    .B(_1942_),
    .C(_1941_),
    .Y(_1948_)
);

NAND3X1 _5447_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1908_),
    .B(_1939_),
    .C(_1936_),
    .Y(_1949_)
);

NAND3X1 _5448_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .B(_1948_),
    .C(_1947_),
    .Y(_1950_)
);

NAND2X1 _5449_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1950_),
    .B(_1946_),
    .Y(_1951_)
);

OAI21X1 _5450_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1907_),
    .B(_1904_),
    .C(_1951_),
    .Y(_1952_)
);

OR2X2 _5451_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1899_),
    .B(_1897_),
    .Y(_1953_)
);

OAI21X1 _5452_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1513_),
    .B(_1413_),
    .C(_1504_),
    .Y(_1955_)
);

OAI21X1 _5453_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1674_),
    .B(_1677_),
    .C(_1679_),
    .Y(_1956_)
);

AOI22X1 _5454_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1956_),
    .B(_1694_),
    .C(_1955_),
    .D(_1698_),
    .Y(_1957_)
);

NOR3X1 _5455_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1414_),
    .B(_1513_),
    .C(_1689_),
    .Y(_1958_)
);

OAI21X1 _5456_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1425_),
    .B(_1432_),
    .C(_1958_),
    .Y(_1959_)
);

AOI21X1 _5457_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1957_),
    .B(_1959_),
    .C(_1847_),
    .Y(_1960_)
);

AND2X2 _5458_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1848_),
    .B(_1840_),
    .Y(_1961_)
);

OAI21X1 _5459_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1960_),
    .B(_1961_),
    .C(_1902_),
    .Y(_1962_)
);

AND2X2 _5460_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1946_),
    .B(_1950_),
    .Y(_1963_)
);

NAND3X1 _5461_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1953_),
    .B(_1963_),
    .C(_1962_),
    .Y(_1964_)
);

NAND2X1 _5462_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1952_),
    .B(_1964_),
    .Y(\partials[7] [19])
);

AOI21X1 _5463_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1901_),
    .B(_1898_),
    .C(_1951_),
    .Y(_1966_)
);

NAND3X1 _5464_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1777_),
    .B(_1966_),
    .C(_1845_),
    .Y(_1967_)
);

OAI21X1 _5465_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1953_),
    .B(_1951_),
    .C(_1950_),
    .Y(_1968_)
);

AOI21X1 _5466_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1966_),
    .B(_1961_),
    .C(_1968_),
    .Y(_1969_)
);

OAI21X1 _5467_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1701_),
    .B(_1967_),
    .C(_1969_),
    .Y(_1970_)
);

OAI21X1 _5468_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1930_),
    .B(_1909_),
    .C(_1938_),
    .Y(_1971_)
);

OAI21X1 _5469_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1922_),
    .B(_1914_),
    .C(_1928_),
    .Y(_1972_)
);

OAI22X1 _5470_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1868_),
    .B(_1917_),
    .C(_1919_),
    .D(_1916_),
    .Y(_1973_)
);

NAND2X1 _5471_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_7_bF$buf3),
    .B(breg[13]),
    .Y(_1974_)
);

NAND2X1 _5472_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf0),
    .B(breg[14]),
    .Y(_1976_)
);

NOR2X1 _5473_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_1976_),
    .Y(_1977_)
);

AND2X2 _5474_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1917_),
    .B(_1976_),
    .Y(_1978_)
);

NOR2X1 _5475_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1977_),
    .B(_1978_),
    .Y(_1979_)
);

XNOR2X1 _5476_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1979_),
    .B(_1974_),
    .Y(_1980_)
);

XOR2X1 _5477_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1980_),
    .B(_1973_),
    .Y(_1981_)
);

XOR2X1 _5478_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1972_),
    .B(_1981_),
    .Y(_1982_)
);

XNOR2X1 _5479_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1971_),
    .B(_1982_),
    .Y(_1983_)
);

NAND2X1 _5480_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .B(_1983_),
    .Y(_1984_)
);

NOR2X1 _5481_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1949_),
    .B(_1983_),
    .Y(_1985_)
);

INVX2 _5482_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1985_),
    .Y(_1986_)
);

NAND2X1 _5483_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1984_),
    .B(_1986_),
    .Y(_1987_)
);

XNOR2X1 _5484_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1970_),
    .B(_1987_),
    .Y(\partials[7] [20])
);

AOI21X1 _5485_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1957_),
    .B(_1959_),
    .C(_1967_),
    .Y(_1988_)
);

NAND2X1 _5486_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1897_),
    .B(_1899_),
    .Y(_1989_)
);

NAND3X1 _5487_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1989_),
    .B(_1953_),
    .C(_1963_),
    .Y(_1990_)
);

INVX1 _5488_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1968_),
    .Y(_1991_)
);

OAI21X1 _5489_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1849_),
    .B(_1990_),
    .C(_1991_),
    .Y(_1992_)
);

INVX1 _5490_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1987_),
    .Y(_1993_)
);

OAI21X1 _5491_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(_1992_),
    .C(_1993_),
    .Y(_1994_)
);

OAI21X1 _5492_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1944_),
    .B(_1935_),
    .C(_1982_),
    .Y(_1996_)
);

OAI21X1 _5493_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1934_),
    .B(_1925_),
    .C(_1981_),
    .Y(_1997_)
);

NAND2X1 _5494_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1973_),
    .B(_1980_),
    .Y(_1998_)
);

INVX1 _5495_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1977_),
    .Y(_1999_)
);

OAI21X1 _5496_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1978_),
    .B(_1974_),
    .C(_1999_),
    .Y(_2000_)
);

OR2X2 _5497_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1855_),
    .B(_1976_),
    .Y(_2001_)
);

OAI21X1 _5498_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_773_),
    .B(_1640_),
    .C(_1790_),
    .Y(_2002_)
);

AND2X2 _5499_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2001_),
    .B(_2002_),
    .Y(_2003_)
);

NAND2X1 _5500_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_2000_),
    .Y(_2004_)
);

INVX1 _5501_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .Y(_2005_)
);

NOR2X1 _5502_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2003_),
    .B(_2000_),
    .Y(_2008_)
);

OAI21X1 _5503_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2005_),
    .B(_2008_),
    .C(_1998_),
    .Y(_2009_)
);

NOR2X1 _5504_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2008_),
    .B(_2005_),
    .Y(_2010_)
);

NAND3X1 _5505_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1973_),
    .B(_1980_),
    .C(_2010_),
    .Y(_2011_)
);

NAND2X1 _5506_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2009_),
    .B(_2011_),
    .Y(_2012_)
);

XOR2X1 _5507_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1997_),
    .B(_2012_),
    .Y(_2013_)
);

INVX1 _5508_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2013_),
    .Y(_2014_)
);

NAND2X1 _5509_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2014_),
    .B(_1996_),
    .Y(_2015_)
);

OR2X2 _5510_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1996_),
    .B(_2014_),
    .Y(_2016_)
);

NAND2X1 _5511_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2015_),
    .B(_2016_),
    .Y(_2017_)
);

INVX1 _5512_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .Y(_2018_)
);

NAND3X1 _5513_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1986_),
    .B(_2018_),
    .C(_1994_),
    .Y(_2019_)
);

NOR2X1 _5514_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1990_),
    .B(_1847_),
    .Y(_2020_)
);

OAI21X1 _5515_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1696_),
    .B(_1700_),
    .C(_2020_),
    .Y(_2021_)
);

AOI21X1 _5516_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1969_),
    .B(_2021_),
    .C(_1987_),
    .Y(_2022_)
);

OAI21X1 _5517_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2022_),
    .B(_1985_),
    .C(_2017_),
    .Y(_2023_)
);

NAND2X1 _5518_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2023_),
    .B(_2019_),
    .Y(\partials[7] [21])
);

NOR2X1 _5519_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_1987_),
    .Y(_2024_)
);

OAI21X1 _5520_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1988_),
    .B(_1992_),
    .C(_2024_),
    .Y(_2025_)
);

OAI21X1 _5521_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2017_),
    .B(_1986_),
    .C(_2016_),
    .Y(_2026_)
);

INVX1 _5522_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2026_),
    .Y(_2029_)
);

AOI21X1 _5523_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(areg_6_bF$buf3),
    .B(breg[14]),
    .C(_1855_),
    .Y(_2030_)
);

XNOR2X1 _5524_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(_2030_),
    .Y(_2031_)
);

OAI21X1 _5525_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1997_),
    .B(_2012_),
    .C(_2011_),
    .Y(_2032_)
);

XNOR2X1 _5526_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2032_),
    .B(_2031_),
    .Y(_2033_)
);

INVX1 _5527_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2033_),
    .Y(_2034_)
);

NAND3X1 _5528_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2029_),
    .B(_2034_),
    .C(_2025_),
    .Y(_2035_)
);

INVX1 _5529_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2024_),
    .Y(_2036_)
);

AOI21X1 _5530_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_1969_),
    .B(_2021_),
    .C(_2036_),
    .Y(_2037_)
);

OAI21X1 _5531_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .B(_2026_),
    .C(_2033_),
    .Y(_2038_)
);

NAND2X1 _5532_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2038_),
    .B(_2035_),
    .Y(\partials[7] [22])
);

OAI21X1 _5533_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2037_),
    .B(_2026_),
    .C(_2034_),
    .Y(_2040_)
);

OAI21X1 _5534_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2004_),
    .B(_1855_),
    .C(_2001_),
    .Y(_2041_)
);

AOI21X1 _5535_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2031_),
    .B(_2032_),
    .C(_2041_),
    .Y(_2042_)
);

NAND2X1 _5536_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2042_),
    .B(_2040_),
    .Y(\partials[7] [23])
);

BUFX2 _5537_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[0]),
    .Y(y[0])
);

BUFX2 _5538_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[1]),
    .Y(y[1])
);

BUFX2 _5539_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[2]),
    .Y(y[2])
);

BUFX2 _5540_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[3]),
    .Y(y[3])
);

BUFX2 _5541_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[4]),
    .Y(y[4])
);

BUFX2 _5542_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[5]),
    .Y(y[5])
);

BUFX2 _5543_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[6]),
    .Y(y[6])
);

BUFX2 _5544_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[7]),
    .Y(y[7])
);

BUFX2 _5545_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[8]),
    .Y(y[8])
);

BUFX2 _5546_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[9]),
    .Y(y[9])
);

BUFX2 _5547_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[10]),
    .Y(y[10])
);

BUFX2 _5548_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[11]),
    .Y(y[11])
);

BUFX2 _5549_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[12]),
    .Y(y[12])
);

BUFX2 _5550_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[13]),
    .Y(y[13])
);

BUFX2 _5551_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[14]),
    .Y(y[14])
);

BUFX2 _5552_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[15]),
    .Y(y[15])
);

BUFX2 _5553_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[16]),
    .Y(y[16])
);

BUFX2 _5554_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[17]),
    .Y(y[17])
);

BUFX2 _5555_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[18]),
    .Y(y[18])
);

BUFX2 _5556_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[19]),
    .Y(y[19])
);

BUFX2 _5557_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[20]),
    .Y(y[20])
);

BUFX2 _5558_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[21]),
    .Y(y[21])
);

BUFX2 _5559_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[22]),
    .Y(y[22])
);

BUFX2 _5560_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[23]),
    .Y(y[23])
);

BUFX2 _5561_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[24]),
    .Y(y[24])
);

BUFX2 _5562_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[25]),
    .Y(y[25])
);

BUFX2 _5563_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[26]),
    .Y(y[26])
);

BUFX2 _5564_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[27]),
    .Y(y[27])
);

BUFX2 _5565_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[28]),
    .Y(y[28])
);

BUFX2 _5566_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[29]),
    .Y(y[29])
);

BUFX2 _5567_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[30]),
    .Y(y[30])
);

BUFX2 _5568_ (
    .gnd(gnd),
    .vdd(vdd),
    .A(_2744_[31]),
    .Y(y[31])
);

DFFPOSX1 _5569_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[0] [0]),
    .Q(\partials[15] [0])
);

DFFPOSX1 _5570_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[7] [1]),
    .Q(\partials[15] [1])
);

DFFPOSX1 _5571_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[7] [2]),
    .Q(\partials[15] [2])
);

DFFPOSX1 _5572_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[7] [3]),
    .Q(\partials[15] [3])
);

DFFPOSX1 _5573_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[7] [4]),
    .Q(\partials[15] [4])
);

DFFPOSX1 _5574_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[7] [5]),
    .Q(\partials[15] [5])
);

DFFPOSX1 _5575_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(\partials[7] [6]),
    .Q(\partials[15] [6])
);

DFFPOSX1 _5576_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(\partials[7] [7]),
    .Q(\partials[15] [7])
);

DFFPOSX1 _5577_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(\partials[7] [8]),
    .Q(\preg[7] [8])
);

DFFPOSX1 _5578_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(\partials[7] [9]),
    .Q(\preg[7] [9])
);

DFFPOSX1 _5579_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[7] [10]),
    .Q(\preg[7] [10])
);

DFFPOSX1 _5580_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[7] [11]),
    .Q(\preg[7] [11])
);

DFFPOSX1 _5581_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[7] [12]),
    .Q(\preg[7] [12])
);

DFFPOSX1 _5582_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[7] [13]),
    .Q(\preg[7] [13])
);

DFFPOSX1 _5583_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[7] [14]),
    .Q(\preg[7] [14])
);

DFFPOSX1 _5584_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[7] [15]),
    .Q(\preg[7] [15])
);

DFFPOSX1 _5585_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(\partials[7] [16]),
    .Q(\preg[7] [16])
);

DFFPOSX1 _5586_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(\partials[7] [17]),
    .Q(\preg[7] [17])
);

DFFPOSX1 _5587_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(\partials[7] [18]),
    .Q(\preg[7] [18])
);

DFFPOSX1 _5588_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(\partials[7] [19]),
    .Q(\preg[7] [19])
);

DFFPOSX1 _5589_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[7] [20]),
    .Q(\preg[7] [20])
);

DFFPOSX1 _5590_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[7] [21]),
    .Q(\preg[7] [21])
);

DFFPOSX1 _5591_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[7] [22]),
    .Q(\preg[7] [22])
);

DFFPOSX1 _5592_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[7] [23]),
    .Q(\preg[7] [23])
);

DFFPOSX1 _5593_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[15] [0]),
    .Q(_2744_[0])
);

DFFPOSX1 _5594_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[15] [1]),
    .Q(_2744_[1])
);

DFFPOSX1 _5595_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(\partials[15] [2]),
    .Q(_2744_[2])
);

DFFPOSX1 _5596_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(\partials[15] [3]),
    .Q(_2744_[3])
);

DFFPOSX1 _5597_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(\partials[15] [4]),
    .Q(_2744_[4])
);

DFFPOSX1 _5598_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(\partials[15] [5]),
    .Q(_2744_[5])
);

DFFPOSX1 _5599_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[15] [6]),
    .Q(_2744_[6])
);

DFFPOSX1 _5600_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[15] [7]),
    .Q(_2744_[7])
);

DFFPOSX1 _5601_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[15] [8]),
    .Q(_2744_[8])
);

DFFPOSX1 _5602_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[15] [9]),
    .Q(_2744_[9])
);

DFFPOSX1 _5603_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[15] [10]),
    .Q(_2744_[10])
);

DFFPOSX1 _5604_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[15] [11]),
    .Q(_2744_[11])
);

DFFPOSX1 _5605_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(\partials[15] [12]),
    .Q(_2744_[12])
);

DFFPOSX1 _5606_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(\partials[15] [13]),
    .Q(_2744_[13])
);

DFFPOSX1 _5607_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(\partials[15] [14]),
    .Q(_2744_[14])
);

DFFPOSX1 _5608_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(\partials[15] [15]),
    .Q(_2744_[15])
);

DFFPOSX1 _5609_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[15] [16]),
    .Q(_2744_[16])
);

DFFPOSX1 _5610_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[15] [17]),
    .Q(_2744_[17])
);

DFFPOSX1 _5611_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[15] [18]),
    .Q(_2744_[18])
);

DFFPOSX1 _5612_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[15] [19]),
    .Q(_2744_[19])
);

DFFPOSX1 _5613_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[15] [20]),
    .Q(_2744_[20])
);

DFFPOSX1 _5614_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[15] [21]),
    .Q(_2744_[21])
);

DFFPOSX1 _5615_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(\partials[15] [22]),
    .Q(_2744_[22])
);

DFFPOSX1 _5616_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(\partials[15] [23]),
    .Q(_2744_[23])
);

DFFPOSX1 _5617_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(\partials[15] [24]),
    .Q(_2744_[24])
);

DFFPOSX1 _5618_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(\partials[15] [25]),
    .Q(_2744_[25])
);

DFFPOSX1 _5619_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(\partials[15] [26]),
    .Q(_2744_[26])
);

DFFPOSX1 _5620_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(\partials[15] [27]),
    .Q(_2744_[27])
);

DFFPOSX1 _5621_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(\partials[15] [28]),
    .Q(_2744_[28])
);

DFFPOSX1 _5622_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(\partials[15] [29]),
    .Q(_2744_[29])
);

DFFPOSX1 _5623_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(\partials[15] [30]),
    .Q(_2744_[30])
);

DFFPOSX1 _5624_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(\partials[15] [31]),
    .Q(_2744_[31])
);

DFFPOSX1 _5625_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(areg[8]),
    .Q(aregp1[8])
);

DFFPOSX1 _5626_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(areg[9]),
    .Q(aregp1[9])
);

DFFPOSX1 _5627_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(areg[10]),
    .Q(aregp1[10])
);

DFFPOSX1 _5628_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(areg[11]),
    .Q(aregp1[11])
);

DFFPOSX1 _5629_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(areg[12]),
    .Q(aregp1[12])
);

DFFPOSX1 _5630_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(areg[13]),
    .Q(aregp1[13])
);

DFFPOSX1 _5631_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(areg[14]),
    .Q(aregp1[14])
);

DFFPOSX1 _5632_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(areg[15]),
    .Q(aregp1[15])
);

DFFPOSX1 _5633_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(breg[0]),
    .Q(bregp1[0])
);

DFFPOSX1 _5634_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(breg[1]),
    .Q(bregp1[1])
);

DFFPOSX1 _5635_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(breg[2]),
    .Q(bregp1[2])
);

DFFPOSX1 _5636_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(breg[3]),
    .Q(bregp1[3])
);

DFFPOSX1 _5637_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(breg[4]),
    .Q(bregp1[4])
);

DFFPOSX1 _5638_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(breg[5]),
    .Q(bregp1[5])
);

DFFPOSX1 _5639_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(breg[6]),
    .Q(bregp1[6])
);

DFFPOSX1 _5640_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(breg[7]),
    .Q(bregp1[7])
);

DFFPOSX1 _5641_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(breg[8]),
    .Q(bregp1[8])
);

DFFPOSX1 _5642_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(breg[9]),
    .Q(bregp1[9])
);

DFFPOSX1 _5643_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(breg[10]),
    .Q(bregp1[10])
);

DFFPOSX1 _5644_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(breg[11]),
    .Q(bregp1[11])
);

DFFPOSX1 _5645_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(breg[12]),
    .Q(bregp1[12])
);

DFFPOSX1 _5646_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(breg[13]),
    .Q(bregp1[13])
);

DFFPOSX1 _5647_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(breg[14]),
    .Q(bregp1[14])
);

DFFPOSX1 _5648_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(breg[15]),
    .Q(bregp1[15])
);

DFFPOSX1 _5649_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(a[0]),
    .Q(areg[0])
);

DFFPOSX1 _5650_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(a[1]),
    .Q(areg[1])
);

DFFPOSX1 _5651_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(a[2]),
    .Q(areg[2])
);

DFFPOSX1 _5652_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(a[3]),
    .Q(areg[3])
);

DFFPOSX1 _5653_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(a[4]),
    .Q(areg[4])
);

DFFPOSX1 _5654_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(a[5]),
    .Q(areg[5])
);

DFFPOSX1 _5655_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(a[6]),
    .Q(areg[6])
);

DFFPOSX1 _5656_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(a[7]),
    .Q(areg[7])
);

DFFPOSX1 _5657_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(a[8]),
    .Q(areg[8])
);

DFFPOSX1 _5658_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(a[9]),
    .Q(areg[9])
);

DFFPOSX1 _5659_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(a[10]),
    .Q(areg[10])
);

DFFPOSX1 _5660_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(a[11]),
    .Q(areg[11])
);

DFFPOSX1 _5661_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(a[12]),
    .Q(areg[12])
);

DFFPOSX1 _5662_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(a[13]),
    .Q(areg[13])
);

DFFPOSX1 _5663_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(a[14]),
    .Q(areg[14])
);

DFFPOSX1 _5664_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(a[15]),
    .Q(areg[15])
);

DFFPOSX1 _5665_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(b[0]),
    .Q(breg[0])
);

DFFPOSX1 _5666_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(b[1]),
    .Q(breg[1])
);

DFFPOSX1 _5667_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(b[2]),
    .Q(breg[2])
);

DFFPOSX1 _5668_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(b[3]),
    .Q(breg[3])
);

DFFPOSX1 _5669_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(b[4]),
    .Q(breg[4])
);

DFFPOSX1 _5670_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(b[5]),
    .Q(breg[5])
);

DFFPOSX1 _5671_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf7),
    .D(b[6]),
    .Q(breg[6])
);

DFFPOSX1 _5672_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf6),
    .D(b[7]),
    .Q(breg[7])
);

DFFPOSX1 _5673_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf5),
    .D(b[8]),
    .Q(breg[8])
);

DFFPOSX1 _5674_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf4),
    .D(b[9]),
    .Q(breg[9])
);

DFFPOSX1 _5675_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf3),
    .D(b[10]),
    .Q(breg[10])
);

DFFPOSX1 _5676_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf2),
    .D(b[11]),
    .Q(breg[11])
);

DFFPOSX1 _5677_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf1),
    .D(b[12]),
    .Q(breg[12])
);

DFFPOSX1 _5678_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf0),
    .D(b[13]),
    .Q(breg[13])
);

DFFPOSX1 _5679_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf9),
    .D(b[14]),
    .Q(breg[14])
);

DFFPOSX1 _5680_ (
    .gnd(gnd),
    .vdd(vdd),
    .CLK(clk_bF$buf8),
    .D(b[15]),
    .Q(breg[15])
);

endmodule
