/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module multiplierCarry(
    input [7:0] a,
    input [7:0] b,
    input clk,
    output [15:0] y
);

wire [7:0] a ;
wire [7:0] b ;
wire [15:0] y ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _19_ ;
wire _512_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _415_ ;
wire _95_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _262_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _165_ ;
wire _394_ ;
wire _259_ ;
wire _488_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _412_ ;
wire _92_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _162_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _197_ ;
wire [7:0] _7_ ;
wire _503_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _215_ ;
wire _444_ ;
wire _253_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _479_ ;
wire _288_ ;
wire [7:0] _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _212_ ;
wire _441_ ;
wire _250_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _153_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire [7:0] _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _150_ ;
wire _206_ ;
wire _435_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _338_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _279_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _203_ ;
wire _432_ ;
wire _241_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _335_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire _238_ ;
wire _467_ ;
wire _276_ ;
wire _33_ ;
wire _179_ ;
wire _71_ ;
wire _200_ ;
wire _523_ ;
wire _103_ ;
wire _332_ ;
wire _68_ ;
wire _141_ ;
wire _370_ ;
wire _426_ ;
wire _235_ ;
wire _464_ ;
wire _273_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _176_ ;
wire _499_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _423_ ;
wire _232_ ;
wire _461_ ;
wire _517_ ;
wire _270_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _173_ ;
wire _229_ ;
wire _458_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _420_ ;
wire _514_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _170_ ;
wire _226_ ;
wire _455_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _167_ ;
wire _396_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _320_ ;
wire _56_ ;
wire _414_ ;
wire _94_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _261_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire [7:0] breg ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _220_ ;
wire [15:0] _9_ ;
wire _505_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _161_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire [7:0] _6_ ;
wire _502_ ;
wire [7:0] areg ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire _214_ ;
wire _443_ ;
wire _252_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire [7:0] _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _211_ ;
wire _440_ ;
wire _305_ ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _152_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire [7:0] _0_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _205_ ;
wire _434_ ;
wire _243_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _337_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _278_ ;
wire _35_ ;
wire _73_ ;
wire _202_ ;
wire _431_ ;
wire _240_ ;
wire _525_ ;
wire _105_ ;
wire _334_ ;
wire _143_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _237_ ;
wire _466_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _178_ ;
wire _70_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _331_ ;
wire _67_ ;
wire [15:0] _560_ ;
wire _140_ ;
wire _425_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _272_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _175_ ;
wire _269_ ;
wire _498_ ;
wire _26_ ;
wire _64_ ;
wire _422_ ;
wire _231_ ;
wire _460_ ;
wire _516_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _172_ ;
wire _228_ ;
wire _457_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _513_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire _225_ ;
wire _454_ ;
wire _263_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _413_ ;
wire _93_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _260_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _163_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire [6:0] _8_ ;
wire _504_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _160_ ;
wire _216_ ;
wire _445_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire [7:0] _5_ ;
wire _501_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _213_ ;
wire _442_ ;
wire _251_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire [7:0] _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _210_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _151_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire _339_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _204_ ;
wire _433_ ;
wire _242_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _336_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _239_ ;
wire _468_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _201_ ;
wire _430_ ;
wire _524_ ;
wire _104_ ;
wire _333_ ;
wire _69_ ;
wire _142_ ;
wire _371_ ;
wire _427_ ;
wire _180_ ;
wire _236_ ;
wire _465_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _177_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _330_ ;
wire _66_ ;
wire _424_ ;
wire _233_ ;
wire _462_ ;
wire _518_ ;
wire _271_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _174_ ;
wire _459_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _421_ ;
wire _230_ ;
wire _515_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _171_ ;
wire _227_ ;
wire _456_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

CLKBUF1 CLKBUF1_insert4 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert3 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert2 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert1 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert0 (
    .A(clk),
    .Y(clk_bF$buf4)
);

NAND3X1 _1000_ (
    .A(_386_),
    .B(_381_),
    .C(_382_),
    .Y(_387_)
);

INVX1 _1001_ (
    .A(_381_),
    .Y(_388_)
);

NOR2X1 _1002_ (
    .A(_367_),
    .B(_380_),
    .Y(_389_)
);

INVX1 _1003_ (
    .A(_386_),
    .Y(_390_)
);

OAI21X1 _1004_ (
    .A(_388_),
    .B(_389_),
    .C(_390_),
    .Y(_391_)
);

AOI21X1 _1005_ (
    .A(_387_),
    .B(_391_),
    .C(_366_),
    .Y(_392_)
);

OAI21X1 _1006_ (
    .A(_388_),
    .B(_389_),
    .C(_386_),
    .Y(_393_)
);

NAND3X1 _1007_ (
    .A(_390_),
    .B(_381_),
    .C(_382_),
    .Y(_394_)
);

AOI21X1 _1008_ (
    .A(_394_),
    .B(_393_),
    .C(_365_),
    .Y(_396_)
);

OAI21X1 _1009_ (
    .A(_338_),
    .B(_335_),
    .C(_329_),
    .Y(_397_)
);

INVX2 _1010_ (
    .A(_397_),
    .Y(_398_)
);

OAI21X1 _1011_ (
    .A(_396_),
    .B(_392_),
    .C(_398_),
    .Y(_399_)
);

OR2X2 _1012_ (
    .A(_396_),
    .B(_398_),
    .Y(_400_)
);

OAI21X1 _1013_ (
    .A(_400_),
    .B(_392_),
    .C(_399_),
    .Y(_401_)
);

NAND3X1 _1014_ (
    .A(_360_),
    .B(_401_),
    .C(_364_),
    .Y(_402_)
);

INVX1 _1015_ (
    .A(_295_),
    .Y(_403_)
);

AOI21X1 _1016_ (
    .A(_355_),
    .B(_358_),
    .C(_359_),
    .Y(_404_)
);

OAI21X1 _1017_ (
    .A(_404_),
    .B(_403_),
    .C(_360_),
    .Y(_405_)
);

NOR2X1 _1018_ (
    .A(_392_),
    .B(_396_),
    .Y(_407_)
);

XNOR2X1 _1019_ (
    .A(_407_),
    .B(_398_),
    .Y(_408_)
);

NAND2X1 _1020_ (
    .A(_408_),
    .B(_405_),
    .Y(_409_)
);

NAND2X1 _1021_ (
    .A(_402_),
    .B(_409_),
    .Y(_410_)
);

XNOR2X1 _1022_ (
    .A(_410_),
    .B(_363_),
    .Y(_9_[10])
);

INVX1 _1023_ (
    .A(_392_),
    .Y(_411_)
);

OAI21X1 _1024_ (
    .A(_396_),
    .B(_398_),
    .C(_411_),
    .Y(_412_)
);

OAI21X1 _1025_ (
    .A(_405_),
    .B(_408_),
    .C(_363_),
    .Y(_413_)
);

NOR2X1 _1026_ (
    .A(_559_),
    .B(_265_),
    .Y(_414_)
);

NAND2X1 _1027_ (
    .A(breg[7]),
    .B(areg[4]),
    .Y(_415_)
);

OAI21X1 _1028_ (
    .A(_370_),
    .B(_371_),
    .C(_374_),
    .Y(_417_)
);

OAI21X1 _1029_ (
    .A(_150_),
    .B(_540_),
    .C(_417_),
    .Y(_418_)
);

OAI21X1 _1030_ (
    .A(_372_),
    .B(_374_),
    .C(_418_),
    .Y(_419_)
);

OAI21X1 _1031_ (
    .A(_305_),
    .B(_308_),
    .C(_419_),
    .Y(_420_)
);

INVX1 _1032_ (
    .A(_419_),
    .Y(_421_)
);

NAND3X1 _1033_ (
    .A(breg[6]),
    .B(areg[5]),
    .C(_421_),
    .Y(_422_)
);

NAND2X1 _1034_ (
    .A(_420_),
    .B(_422_),
    .Y(_423_)
);

XNOR2X1 _1035_ (
    .A(_423_),
    .B(_415_),
    .Y(_424_)
);

OAI21X1 _1036_ (
    .A(_379_),
    .B(_368_),
    .C(_376_),
    .Y(_425_)
);

NAND2X1 _1037_ (
    .A(_368_),
    .B(_379_),
    .Y(_426_)
);

NAND2X1 _1038_ (
    .A(_426_),
    .B(_425_),
    .Y(_428_)
);

NOR2X1 _1039_ (
    .A(_46_),
    .B(_287_),
    .Y(_429_)
);

XNOR2X1 _1040_ (
    .A(_428_),
    .B(_429_),
    .Y(_430_)
);

XOR2X1 _1041_ (
    .A(_430_),
    .B(_424_),
    .Y(_431_)
);

NAND2X1 _1042_ (
    .A(_414_),
    .B(_431_),
    .Y(_432_)
);

OR2X2 _1043_ (
    .A(_431_),
    .B(_414_),
    .Y(_433_)
);

NAND2X1 _1044_ (
    .A(_432_),
    .B(_433_),
    .Y(_434_)
);

OAI21X1 _1045_ (
    .A(_389_),
    .B(_386_),
    .C(_381_),
    .Y(_435_)
);

XNOR2X1 _1046_ (
    .A(_434_),
    .B(_435_),
    .Y(_436_)
);

INVX1 _1047_ (
    .A(_436_),
    .Y(_437_)
);

NAND3X1 _1048_ (
    .A(_409_),
    .B(_437_),
    .C(_413_),
    .Y(_439_)
);

INVX1 _1049_ (
    .A(_363_),
    .Y(_440_)
);

NAND2X1 _1050_ (
    .A(_440_),
    .B(_409_),
    .Y(_441_)
);

NAND3X1 _1051_ (
    .A(_402_),
    .B(_436_),
    .C(_441_),
    .Y(_442_)
);

NAND2X1 _1052_ (
    .A(_439_),
    .B(_442_),
    .Y(_443_)
);

XNOR2X1 _1053_ (
    .A(_443_),
    .B(_412_),
    .Y(_9_[11])
);

INVX1 _1054_ (
    .A(_433_),
    .Y(_444_)
);

INVX1 _1055_ (
    .A(_435_),
    .Y(_445_)
);

OAI21X1 _1056_ (
    .A(_444_),
    .B(_445_),
    .C(_432_),
    .Y(_446_)
);

NAND2X1 _1057_ (
    .A(_412_),
    .B(_439_),
    .Y(_447_)
);

NOR2X1 _1058_ (
    .A(_150_),
    .B(_308_),
    .Y(_449_)
);

OAI21X1 _1059_ (
    .A(_150_),
    .B(_25_),
    .C(_422_),
    .Y(_450_)
);

NAND2X1 _1060_ (
    .A(_420_),
    .B(_450_),
    .Y(_451_)
);

OAI21X1 _1061_ (
    .A(_305_),
    .B(_287_),
    .C(_451_),
    .Y(_452_)
);

INVX1 _1062_ (
    .A(_451_),
    .Y(_453_)
);

NAND3X1 _1063_ (
    .A(breg[6]),
    .B(areg[6]),
    .C(_453_),
    .Y(_454_)
);

NAND2X1 _1064_ (
    .A(_452_),
    .B(_454_),
    .Y(_455_)
);

XOR2X1 _1065_ (
    .A(_455_),
    .B(_449_),
    .Y(_456_)
);

NAND2X1 _1066_ (
    .A(_429_),
    .B(_428_),
    .Y(_457_)
);

NAND2X1 _1067_ (
    .A(_424_),
    .B(_457_),
    .Y(_458_)
);

OAI21X1 _1068_ (
    .A(_428_),
    .B(_429_),
    .C(_458_),
    .Y(_460_)
);

OAI21X1 _1069_ (
    .A(_46_),
    .B(_265_),
    .C(_460_),
    .Y(_461_)
);

NOR2X1 _1070_ (
    .A(_46_),
    .B(_265_),
    .Y(_462_)
);

INVX1 _1071_ (
    .A(_462_),
    .Y(_463_)
);

NOR2X1 _1072_ (
    .A(_463_),
    .B(_460_),
    .Y(_464_)
);

INVX1 _1073_ (
    .A(_464_),
    .Y(_465_)
);

NAND2X1 _1074_ (
    .A(_461_),
    .B(_465_),
    .Y(_466_)
);

XNOR2X1 _1075_ (
    .A(_466_),
    .B(_456_),
    .Y(_467_)
);

NAND3X1 _1076_ (
    .A(_442_),
    .B(_467_),
    .C(_447_),
    .Y(_468_)
);

INVX1 _1077_ (
    .A(_412_),
    .Y(_469_)
);

AOI21X1 _1078_ (
    .A(_360_),
    .B(_364_),
    .C(_401_),
    .Y(_470_)
);

AOI21X1 _1079_ (
    .A(_363_),
    .B(_402_),
    .C(_470_),
    .Y(_471_)
);

OAI21X1 _1080_ (
    .A(_471_),
    .B(_437_),
    .C(_469_),
    .Y(_472_)
);

INVX1 _1081_ (
    .A(_467_),
    .Y(_473_)
);

NAND3X1 _1082_ (
    .A(_439_),
    .B(_473_),
    .C(_472_),
    .Y(_474_)
);

NAND2X1 _1083_ (
    .A(_474_),
    .B(_468_),
    .Y(_475_)
);

XNOR2X1 _1084_ (
    .A(_475_),
    .B(_446_),
    .Y(_9_[12])
);

INVX1 _1085_ (
    .A(_461_),
    .Y(_476_)
);

OAI21X1 _1086_ (
    .A(_456_),
    .B(_476_),
    .C(_465_),
    .Y(_477_)
);

INVX1 _1087_ (
    .A(_446_),
    .Y(_478_)
);

AOI21X1 _1088_ (
    .A(_439_),
    .B(_472_),
    .C(_473_),
    .Y(_480_)
);

OAI21X1 _1089_ (
    .A(_480_),
    .B(_478_),
    .C(_474_),
    .Y(_481_)
);

NOR2X1 _1090_ (
    .A(_150_),
    .B(_287_),
    .Y(_482_)
);

INVX1 _1091_ (
    .A(_482_),
    .Y(_483_)
);

OAI21X1 _1092_ (
    .A(_150_),
    .B(_308_),
    .C(_454_),
    .Y(_484_)
);

NAND2X1 _1093_ (
    .A(_452_),
    .B(_484_),
    .Y(_485_)
);

OAI21X1 _1094_ (
    .A(_305_),
    .B(_265_),
    .C(_485_),
    .Y(_486_)
);

NOR2X1 _1095_ (
    .A(_305_),
    .B(_265_),
    .Y(_487_)
);

INVX1 _1096_ (
    .A(_487_),
    .Y(_488_)
);

NOR2X1 _1097_ (
    .A(_488_),
    .B(_485_),
    .Y(_489_)
);

INVX1 _1098_ (
    .A(_489_),
    .Y(_492_)
);

NAND2X1 _1099_ (
    .A(_486_),
    .B(_492_),
    .Y(_493_)
);

XNOR2X1 _1100_ (
    .A(_493_),
    .B(_483_),
    .Y(_494_)
);

INVX2 _1101_ (
    .A(_494_),
    .Y(_495_)
);

NOR2X1 _1102_ (
    .A(_495_),
    .B(_481_),
    .Y(_496_)
);

NAND2X1 _1103_ (
    .A(_446_),
    .B(_468_),
    .Y(_497_)
);

AOI21X1 _1104_ (
    .A(_474_),
    .B(_497_),
    .C(_494_),
    .Y(_498_)
);

OAI21X1 _1105_ (
    .A(_496_),
    .B(_498_),
    .C(_477_),
    .Y(_499_)
);

INVX1 _1106_ (
    .A(_477_),
    .Y(_500_)
);

NAND3X1 _1107_ (
    .A(_474_),
    .B(_494_),
    .C(_497_),
    .Y(_501_)
);

NAND2X1 _1108_ (
    .A(_495_),
    .B(_481_),
    .Y(_503_)
);

NAND3X1 _1109_ (
    .A(_500_),
    .B(_501_),
    .C(_503_),
    .Y(_504_)
);

NAND2X1 _1110_ (
    .A(_504_),
    .B(_499_),
    .Y(_9_[13])
);

AOI21X1 _1111_ (
    .A(_442_),
    .B(_447_),
    .C(_467_),
    .Y(_505_)
);

AOI21X1 _1112_ (
    .A(_446_),
    .B(_468_),
    .C(_505_),
    .Y(_506_)
);

OAI21X1 _1113_ (
    .A(_506_),
    .B(_494_),
    .C(_500_),
    .Y(_507_)
);

NOR2X1 _1114_ (
    .A(_150_),
    .B(_265_),
    .Y(_508_)
);

INVX1 _1115_ (
    .A(_508_),
    .Y(_509_)
);

AOI21X1 _1116_ (
    .A(_482_),
    .B(_486_),
    .C(_489_),
    .Y(_510_)
);

OR2X2 _1117_ (
    .A(_510_),
    .B(_509_),
    .Y(_511_)
);

OAI21X1 _1118_ (
    .A(_150_),
    .B(_265_),
    .C(_510_),
    .Y(_513_)
);

AND2X2 _1119_ (
    .A(_511_),
    .B(_513_),
    .Y(_514_)
);

INVX1 _1120_ (
    .A(_514_),
    .Y(_515_)
);

NAND3X1 _1121_ (
    .A(_501_),
    .B(_515_),
    .C(_507_),
    .Y(_516_)
);

OAI21X1 _1122_ (
    .A(_481_),
    .B(_495_),
    .C(_477_),
    .Y(_517_)
);

NAND3X1 _1123_ (
    .A(_503_),
    .B(_514_),
    .C(_517_),
    .Y(_518_)
);

NAND2X1 _1124_ (
    .A(_516_),
    .B(_518_),
    .Y(_9_[14])
);

AOI21X1 _1125_ (
    .A(_477_),
    .B(_501_),
    .C(_498_),
    .Y(_519_)
);

OAI21X1 _1126_ (
    .A(_519_),
    .B(_509_),
    .C(_511_),
    .Y(_8_[6])
);

BUFX2 _1127_ (
    .A(_560_[0]),
    .Y(y[0])
);

BUFX2 _1128_ (
    .A(_560_[1]),
    .Y(y[1])
);

BUFX2 _1129_ (
    .A(_560_[2]),
    .Y(y[2])
);

BUFX2 _1130_ (
    .A(_560_[3]),
    .Y(y[3])
);

BUFX2 _1131_ (
    .A(_560_[4]),
    .Y(y[4])
);

BUFX2 _1132_ (
    .A(_560_[5]),
    .Y(y[5])
);

BUFX2 _1133_ (
    .A(_560_[6]),
    .Y(y[6])
);

BUFX2 _1134_ (
    .A(_560_[7]),
    .Y(y[7])
);

BUFX2 _1135_ (
    .A(_560_[8]),
    .Y(y[8])
);

BUFX2 _1136_ (
    .A(_560_[9]),
    .Y(y[9])
);

BUFX2 _1137_ (
    .A(_560_[10]),
    .Y(y[10])
);

BUFX2 _1138_ (
    .A(_560_[11]),
    .Y(y[11])
);

BUFX2 _1139_ (
    .A(_560_[12]),
    .Y(y[12])
);

BUFX2 _1140_ (
    .A(_560_[13]),
    .Y(y[13])
);

BUFX2 _1141_ (
    .A(_560_[14]),
    .Y(y[14])
);

BUFX2 _1142_ (
    .A(_560_[15]),
    .Y(y[15])
);

DFFPOSX1 _1143_ (
    .CLK(clk_bF$buf4),
    .D(_9_[8]),
    .Q(_560_[8])
);

DFFPOSX1 _1144_ (
    .CLK(clk_bF$buf3),
    .D(_9_[9]),
    .Q(_560_[9])
);

DFFPOSX1 _1145_ (
    .CLK(clk_bF$buf2),
    .D(_9_[10]),
    .Q(_560_[10])
);

DFFPOSX1 _1146_ (
    .CLK(clk_bF$buf1),
    .D(_9_[11]),
    .Q(_560_[11])
);

DFFPOSX1 _1147_ (
    .CLK(clk_bF$buf0),
    .D(_9_[12]),
    .Q(_560_[12])
);

DFFPOSX1 _1148_ (
    .CLK(clk_bF$buf4),
    .D(_9_[13]),
    .Q(_560_[13])
);

DFFPOSX1 _1149_ (
    .CLK(clk_bF$buf3),
    .D(_9_[14]),
    .Q(_560_[14])
);

DFFPOSX1 _1150_ (
    .CLK(clk_bF$buf2),
    .D(_8_[6]),
    .Q(_560_[15])
);

DFFPOSX1 _1151_ (
    .CLK(clk_bF$buf1),
    .D(a[0]),
    .Q(areg[0])
);

DFFPOSX1 _1152_ (
    .CLK(clk_bF$buf0),
    .D(a[1]),
    .Q(areg[1])
);

DFFPOSX1 _1153_ (
    .CLK(clk_bF$buf4),
    .D(a[2]),
    .Q(areg[2])
);

DFFPOSX1 _1154_ (
    .CLK(clk_bF$buf3),
    .D(a[3]),
    .Q(areg[3])
);

DFFPOSX1 _1155_ (
    .CLK(clk_bF$buf2),
    .D(a[4]),
    .Q(areg[4])
);

DFFPOSX1 _1156_ (
    .CLK(clk_bF$buf1),
    .D(a[5]),
    .Q(areg[5])
);

DFFPOSX1 _1157_ (
    .CLK(clk_bF$buf0),
    .D(a[6]),
    .Q(areg[6])
);

DFFPOSX1 _1158_ (
    .CLK(clk_bF$buf4),
    .D(a[7]),
    .Q(areg[7])
);

DFFPOSX1 _1159_ (
    .CLK(clk_bF$buf3),
    .D(b[0]),
    .Q(breg[0])
);

DFFPOSX1 _1160_ (
    .CLK(clk_bF$buf2),
    .D(b[1]),
    .Q(breg[1])
);

DFFPOSX1 _1161_ (
    .CLK(clk_bF$buf1),
    .D(b[2]),
    .Q(breg[2])
);

DFFPOSX1 _1162_ (
    .CLK(clk_bF$buf0),
    .D(b[3]),
    .Q(breg[3])
);

DFFPOSX1 _1163_ (
    .CLK(clk_bF$buf4),
    .D(b[4]),
    .Q(breg[4])
);

DFFPOSX1 _1164_ (
    .CLK(clk_bF$buf3),
    .D(b[5]),
    .Q(breg[5])
);

DFFPOSX1 _1165_ (
    .CLK(clk_bF$buf2),
    .D(b[6]),
    .Q(breg[6])
);

DFFPOSX1 _1166_ (
    .CLK(clk_bF$buf1),
    .D(b[7]),
    .Q(breg[7])
);

DFFPOSX1 _1167_ (
    .CLK(clk_bF$buf0),
    .D(_0_[0]),
    .Q(_560_[0])
);

DFFPOSX1 _1168_ (
    .CLK(clk_bF$buf4),
    .D(_7_[0]),
    .Q(_560_[1])
);

DFFPOSX1 _1169_ (
    .CLK(clk_bF$buf3),
    .D(_1_[0]),
    .Q(_560_[2])
);

DFFPOSX1 _1170_ (
    .CLK(clk_bF$buf2),
    .D(_2_[0]),
    .Q(_560_[3])
);

DFFPOSX1 _1171_ (
    .CLK(clk_bF$buf1),
    .D(_3_[0]),
    .Q(_560_[4])
);

DFFPOSX1 _1172_ (
    .CLK(clk_bF$buf0),
    .D(_4_[0]),
    .Q(_560_[5])
);

DFFPOSX1 _1173_ (
    .CLK(clk_bF$buf4),
    .D(_5_[0]),
    .Q(_560_[6])
);

DFFPOSX1 _1174_ (
    .CLK(clk_bF$buf3),
    .D(_6_[0]),
    .Q(_560_[7])
);

INVX1 _561_ (
    .A(areg[0]),
    .Y(_243_)
);

INVX4 _562_ (
    .A(breg[0]),
    .Y(_244_)
);

NOR2X1 _563_ (
    .A(_243_),
    .B(_244_),
    .Y(_0_[0])
);

INVX4 _564_ (
    .A(areg[7]),
    .Y(_265_)
);

NOR2X1 _565_ (
    .A(_244_),
    .B(_265_),
    .Y(_276_)
);

INVX4 _566_ (
    .A(areg[6]),
    .Y(_287_)
);

NOR2X1 _567_ (
    .A(_244_),
    .B(_287_),
    .Y(_297_)
);

INVX4 _568_ (
    .A(areg[5]),
    .Y(_308_)
);

INVX4 _569_ (
    .A(breg[1]),
    .Y(_319_)
);

NOR2X1 _570_ (
    .A(_308_),
    .B(_319_),
    .Y(_330_)
);

INVX2 _571_ (
    .A(_330_),
    .Y(_341_)
);

INVX4 _572_ (
    .A(areg[2]),
    .Y(_352_)
);

INVX4 _573_ (
    .A(breg[2]),
    .Y(_362_)
);

NOR2X1 _574_ (
    .A(_352_),
    .B(_362_),
    .Y(_373_)
);

INVX2 _575_ (
    .A(_373_),
    .Y(_384_)
);

NAND2X1 _576_ (
    .A(areg[0]),
    .B(breg[3]),
    .Y(_395_)
);

NAND2X1 _577_ (
    .A(areg[1]),
    .B(breg[2]),
    .Y(_406_)
);

NAND2X1 _578_ (
    .A(areg[1]),
    .B(breg[3]),
    .Y(_416_)
);

NAND2X1 _579_ (
    .A(areg[0]),
    .B(breg[4]),
    .Y(_427_)
);

NOR2X1 _580_ (
    .A(_416_),
    .B(_427_),
    .Y(_438_)
);

AND2X2 _581_ (
    .A(areg[1]),
    .B(breg[3]),
    .Y(_448_)
);

AND2X2 _582_ (
    .A(areg[0]),
    .B(breg[4]),
    .Y(_459_)
);

NOR2X1 _583_ (
    .A(_448_),
    .B(_459_),
    .Y(_479_)
);

OAI22X1 _584_ (
    .A(_395_),
    .B(_406_),
    .C(_479_),
    .D(_438_),
    .Y(_490_)
);

NAND2X1 _585_ (
    .A(areg[0]),
    .B(breg[2]),
    .Y(_491_)
);

INVX1 _586_ (
    .A(_491_),
    .Y(_502_)
);

NAND3X1 _587_ (
    .A(_427_),
    .B(_448_),
    .C(_502_),
    .Y(_512_)
);

NAND3X1 _588_ (
    .A(_384_),
    .B(_512_),
    .C(_490_),
    .Y(_520_)
);

NOR2X1 _589_ (
    .A(_395_),
    .B(_406_),
    .Y(_521_)
);

NAND2X1 _590_ (
    .A(_448_),
    .B(_459_),
    .Y(_522_)
);

INVX2 _591_ (
    .A(areg[1]),
    .Y(_523_)
);

INVX4 _592_ (
    .A(breg[3]),
    .Y(_524_)
);

OAI21X1 _593_ (
    .A(_523_),
    .B(_524_),
    .C(_427_),
    .Y(_525_)
);

AOI21X1 _594_ (
    .A(_525_),
    .B(_522_),
    .C(_521_),
    .Y(_526_)
);

INVX1 _595_ (
    .A(_512_),
    .Y(_527_)
);

OAI21X1 _596_ (
    .A(_527_),
    .B(_526_),
    .C(_373_),
    .Y(_528_)
);

AND2X2 _597_ (
    .A(areg[0]),
    .B(breg[1]),
    .Y(_529_)
);

INVX1 _598_ (
    .A(_529_),
    .Y(_530_)
);

AND2X2 _599_ (
    .A(areg[0]),
    .B(breg[3]),
    .Y(_531_)
);

AND2X2 _600_ (
    .A(areg[1]),
    .B(breg[2]),
    .Y(_532_)
);

NOR2X1 _601_ (
    .A(_531_),
    .B(_532_),
    .Y(_533_)
);

OAI22X1 _602_ (
    .A(_406_),
    .B(_530_),
    .C(_533_),
    .D(_521_),
    .Y(_534_)
);

NAND3X1 _603_ (
    .A(_395_),
    .B(_532_),
    .C(_529_),
    .Y(_535_)
);

OAI21X1 _604_ (
    .A(_352_),
    .B(_319_),
    .C(_535_),
    .Y(_536_)
);

NAND2X1 _605_ (
    .A(_536_),
    .B(_534_),
    .Y(_537_)
);

AOI21X1 _606_ (
    .A(_520_),
    .B(_528_),
    .C(_537_),
    .Y(_538_)
);

NAND3X1 _607_ (
    .A(_537_),
    .B(_520_),
    .C(_528_),
    .Y(_539_)
);

INVX4 _608_ (
    .A(areg[3]),
    .Y(_540_)
);

NOR2X1 _609_ (
    .A(_540_),
    .B(_319_),
    .Y(_541_)
);

AOI21X1 _610_ (
    .A(_541_),
    .B(_539_),
    .C(_538_),
    .Y(_542_)
);

NOR2X1 _611_ (
    .A(_540_),
    .B(_362_),
    .Y(_543_)
);

INVX2 _612_ (
    .A(_543_),
    .Y(_544_)
);

OAI21X1 _613_ (
    .A(_352_),
    .B(_362_),
    .C(_512_),
    .Y(_545_)
);

NAND2X1 _614_ (
    .A(_490_),
    .B(_545_),
    .Y(_546_)
);

NOR2X1 _615_ (
    .A(_352_),
    .B(_524_),
    .Y(_547_)
);

INVX2 _616_ (
    .A(_547_),
    .Y(_548_)
);

NAND2X1 _617_ (
    .A(areg[1]),
    .B(breg[4]),
    .Y(_549_)
);

NAND2X1 _618_ (
    .A(areg[0]),
    .B(breg[5]),
    .Y(_550_)
);

NOR2X1 _619_ (
    .A(_549_),
    .B(_550_),
    .Y(_551_)
);

AND2X2 _620_ (
    .A(_549_),
    .B(_550_),
    .Y(_552_)
);

OAI21X1 _621_ (
    .A(_552_),
    .B(_551_),
    .C(_522_),
    .Y(_553_)
);

AND2X2 _622_ (
    .A(areg[1]),
    .B(breg[4]),
    .Y(_554_)
);

NAND3X1 _623_ (
    .A(_550_),
    .B(_531_),
    .C(_554_),
    .Y(_555_)
);

NAND3X1 _624_ (
    .A(_548_),
    .B(_555_),
    .C(_553_),
    .Y(_556_)
);

AND2X2 _625_ (
    .A(areg[0]),
    .B(breg[5]),
    .Y(_557_)
);

NAND2X1 _626_ (
    .A(_554_),
    .B(_557_),
    .Y(_558_)
);

INVX4 _627_ (
    .A(breg[4]),
    .Y(_559_)
);

OAI21X1 _628_ (
    .A(_523_),
    .B(_559_),
    .C(_550_),
    .Y(_10_)
);

AOI21X1 _629_ (
    .A(_10_),
    .B(_558_),
    .C(_438_),
    .Y(_11_)
);

INVX2 _630_ (
    .A(_555_),
    .Y(_12_)
);

OAI21X1 _631_ (
    .A(_11_),
    .B(_12_),
    .C(_547_),
    .Y(_13_)
);

NAND3X1 _632_ (
    .A(_556_),
    .B(_13_),
    .C(_546_),
    .Y(_14_)
);

OAI21X1 _633_ (
    .A(_526_),
    .B(_384_),
    .C(_512_),
    .Y(_15_)
);

OAI21X1 _634_ (
    .A(_11_),
    .B(_12_),
    .C(_548_),
    .Y(_16_)
);

NAND3X1 _635_ (
    .A(_547_),
    .B(_555_),
    .C(_553_),
    .Y(_17_)
);

NAND3X1 _636_ (
    .A(_17_),
    .B(_15_),
    .C(_16_),
    .Y(_18_)
);

NAND3X1 _637_ (
    .A(_544_),
    .B(_18_),
    .C(_14_),
    .Y(_19_)
);

AOI21X1 _638_ (
    .A(_17_),
    .B(_16_),
    .C(_15_),
    .Y(_20_)
);

AOI21X1 _639_ (
    .A(_556_),
    .B(_13_),
    .C(_546_),
    .Y(_21_)
);

OAI21X1 _640_ (
    .A(_20_),
    .B(_21_),
    .C(_543_),
    .Y(_22_)
);

AOI21X1 _641_ (
    .A(_19_),
    .B(_22_),
    .C(_542_),
    .Y(_23_)
);

NAND3X1 _642_ (
    .A(_19_),
    .B(_22_),
    .C(_542_),
    .Y(_24_)
);

INVX4 _643_ (
    .A(areg[4]),
    .Y(_25_)
);

NOR2X1 _644_ (
    .A(_25_),
    .B(_319_),
    .Y(_26_)
);

AOI21X1 _645_ (
    .A(_26_),
    .B(_24_),
    .C(_23_),
    .Y(_27_)
);

NOR2X1 _646_ (
    .A(_25_),
    .B(_362_),
    .Y(_28_)
);

INVX2 _647_ (
    .A(_28_),
    .Y(_29_)
);

AOI21X1 _648_ (
    .A(_543_),
    .B(_14_),
    .C(_21_),
    .Y(_30_)
);

NOR2X1 _649_ (
    .A(_540_),
    .B(_524_),
    .Y(_31_)
);

INVX2 _650_ (
    .A(_31_),
    .Y(_32_)
);

AOI21X1 _651_ (
    .A(_547_),
    .B(_553_),
    .C(_12_),
    .Y(_33_)
);

NOR2X1 _652_ (
    .A(_352_),
    .B(_559_),
    .Y(_34_)
);

INVX2 _653_ (
    .A(_34_),
    .Y(_35_)
);

NAND2X1 _654_ (
    .A(areg[1]),
    .B(breg[5]),
    .Y(_36_)
);

NAND2X1 _655_ (
    .A(areg[0]),
    .B(breg[6]),
    .Y(_37_)
);

NOR2X1 _656_ (
    .A(_36_),
    .B(_37_),
    .Y(_38_)
);

AND2X2 _657_ (
    .A(_36_),
    .B(_37_),
    .Y(_39_)
);

OAI21X1 _658_ (
    .A(_39_),
    .B(_38_),
    .C(_558_),
    .Y(_40_)
);

AND2X2 _659_ (
    .A(areg[1]),
    .B(breg[5]),
    .Y(_41_)
);

NAND3X1 _660_ (
    .A(_37_),
    .B(_459_),
    .C(_41_),
    .Y(_42_)
);

NAND3X1 _661_ (
    .A(_35_),
    .B(_42_),
    .C(_40_),
    .Y(_43_)
);

AND2X2 _662_ (
    .A(areg[0]),
    .B(breg[6]),
    .Y(_44_)
);

NAND2X1 _663_ (
    .A(_41_),
    .B(_44_),
    .Y(_45_)
);

INVX4 _664_ (
    .A(breg[5]),
    .Y(_46_)
);

OAI21X1 _665_ (
    .A(_523_),
    .B(_46_),
    .C(_37_),
    .Y(_47_)
);

AOI21X1 _666_ (
    .A(_47_),
    .B(_45_),
    .C(_551_),
    .Y(_48_)
);

INVX2 _667_ (
    .A(_42_),
    .Y(_49_)
);

OAI21X1 _668_ (
    .A(_48_),
    .B(_49_),
    .C(_34_),
    .Y(_50_)
);

NAND3X1 _669_ (
    .A(_43_),
    .B(_33_),
    .C(_50_),
    .Y(_51_)
);

OAI21X1 _670_ (
    .A(_11_),
    .B(_548_),
    .C(_555_),
    .Y(_52_)
);

OAI21X1 _671_ (
    .A(_48_),
    .B(_49_),
    .C(_35_),
    .Y(_53_)
);

NAND3X1 _672_ (
    .A(_34_),
    .B(_42_),
    .C(_40_),
    .Y(_54_)
);

NAND3X1 _673_ (
    .A(_54_),
    .B(_52_),
    .C(_53_),
    .Y(_55_)
);

NAND3X1 _674_ (
    .A(_32_),
    .B(_51_),
    .C(_55_),
    .Y(_56_)
);

AOI21X1 _675_ (
    .A(_54_),
    .B(_53_),
    .C(_52_),
    .Y(_57_)
);

AOI21X1 _676_ (
    .A(_43_),
    .B(_50_),
    .C(_33_),
    .Y(_58_)
);

OAI21X1 _677_ (
    .A(_57_),
    .B(_58_),
    .C(_31_),
    .Y(_59_)
);

NAND3X1 _678_ (
    .A(_56_),
    .B(_30_),
    .C(_59_),
    .Y(_60_)
);

OAI21X1 _679_ (
    .A(_20_),
    .B(_544_),
    .C(_18_),
    .Y(_61_)
);

OAI21X1 _680_ (
    .A(_57_),
    .B(_58_),
    .C(_32_),
    .Y(_62_)
);

NAND3X1 _681_ (
    .A(_31_),
    .B(_51_),
    .C(_55_),
    .Y(_63_)
);

NAND3X1 _682_ (
    .A(_63_),
    .B(_61_),
    .C(_62_),
    .Y(_64_)
);

NAND3X1 _683_ (
    .A(_29_),
    .B(_60_),
    .C(_64_),
    .Y(_65_)
);

AOI21X1 _684_ (
    .A(_63_),
    .B(_62_),
    .C(_61_),
    .Y(_66_)
);

AOI21X1 _685_ (
    .A(_56_),
    .B(_59_),
    .C(_30_),
    .Y(_67_)
);

OAI21X1 _686_ (
    .A(_66_),
    .B(_67_),
    .C(_28_),
    .Y(_68_)
);

NAND3X1 _687_ (
    .A(_65_),
    .B(_27_),
    .C(_68_),
    .Y(_69_)
);

OAI21X1 _688_ (
    .A(_527_),
    .B(_526_),
    .C(_384_),
    .Y(_70_)
);

NAND3X1 _689_ (
    .A(_373_),
    .B(_512_),
    .C(_490_),
    .Y(_71_)
);

AND2X2 _690_ (
    .A(_534_),
    .B(_536_),
    .Y(_72_)
);

NAND3X1 _691_ (
    .A(_71_),
    .B(_70_),
    .C(_72_),
    .Y(_73_)
);

AOI21X1 _692_ (
    .A(_71_),
    .B(_70_),
    .C(_72_),
    .Y(_74_)
);

INVX1 _693_ (
    .A(_541_),
    .Y(_75_)
);

OAI21X1 _694_ (
    .A(_74_),
    .B(_75_),
    .C(_73_),
    .Y(_76_)
);

OAI21X1 _695_ (
    .A(_20_),
    .B(_21_),
    .C(_544_),
    .Y(_77_)
);

NAND3X1 _696_ (
    .A(_543_),
    .B(_18_),
    .C(_14_),
    .Y(_78_)
);

NAND3X1 _697_ (
    .A(_78_),
    .B(_77_),
    .C(_76_),
    .Y(_79_)
);

AOI21X1 _698_ (
    .A(_78_),
    .B(_77_),
    .C(_76_),
    .Y(_80_)
);

INVX1 _699_ (
    .A(_26_),
    .Y(_81_)
);

OAI21X1 _700_ (
    .A(_80_),
    .B(_81_),
    .C(_79_),
    .Y(_82_)
);

OAI21X1 _701_ (
    .A(_66_),
    .B(_67_),
    .C(_29_),
    .Y(_83_)
);

NAND3X1 _702_ (
    .A(_28_),
    .B(_60_),
    .C(_64_),
    .Y(_84_)
);

NAND3X1 _703_ (
    .A(_84_),
    .B(_82_),
    .C(_83_),
    .Y(_85_)
);

NAND3X1 _704_ (
    .A(_341_),
    .B(_69_),
    .C(_85_),
    .Y(_86_)
);

AOI21X1 _705_ (
    .A(_84_),
    .B(_83_),
    .C(_82_),
    .Y(_87_)
);

AOI21X1 _706_ (
    .A(_65_),
    .B(_68_),
    .C(_27_),
    .Y(_88_)
);

OAI21X1 _707_ (
    .A(_87_),
    .B(_88_),
    .C(_330_),
    .Y(_89_)
);

NOR2X1 _708_ (
    .A(_244_),
    .B(_308_),
    .Y(_90_)
);

INVX1 _709_ (
    .A(_90_),
    .Y(_91_)
);

OAI21X1 _710_ (
    .A(_23_),
    .B(_80_),
    .C(_26_),
    .Y(_92_)
);

NAND3X1 _711_ (
    .A(_81_),
    .B(_24_),
    .C(_79_),
    .Y(_93_)
);

NAND3X1 _712_ (
    .A(_91_),
    .B(_93_),
    .C(_92_),
    .Y(_94_)
);

NOR2X1 _713_ (
    .A(_244_),
    .B(_25_),
    .Y(_95_)
);

OAI21X1 _714_ (
    .A(_538_),
    .B(_74_),
    .C(_75_),
    .Y(_96_)
);

NAND3X1 _715_ (
    .A(_541_),
    .B(_539_),
    .C(_73_),
    .Y(_97_)
);

AOI21X1 _716_ (
    .A(_97_),
    .B(_96_),
    .C(_95_),
    .Y(_98_)
);

NOR2X1 _717_ (
    .A(_352_),
    .B(_319_),
    .Y(_99_)
);

NAND2X1 _718_ (
    .A(_535_),
    .B(_534_),
    .Y(_100_)
);

XOR2X1 _719_ (
    .A(_100_),
    .B(_99_),
    .Y(_101_)
);

OAI21X1 _720_ (
    .A(_244_),
    .B(_540_),
    .C(_101_),
    .Y(_102_)
);

OAI21X1 _721_ (
    .A(_523_),
    .B(_319_),
    .C(_491_),
    .Y(_103_)
);

OAI21X1 _722_ (
    .A(_530_),
    .B(_406_),
    .C(_103_),
    .Y(_104_)
);

OAI21X1 _723_ (
    .A(_244_),
    .B(_352_),
    .C(_104_),
    .Y(_105_)
);

NOR2X1 _724_ (
    .A(_244_),
    .B(_523_),
    .Y(_106_)
);

NAND2X1 _725_ (
    .A(_529_),
    .B(_106_),
    .Y(_107_)
);

INVX2 _726_ (
    .A(_107_),
    .Y(_108_)
);

NOR2X1 _727_ (
    .A(_244_),
    .B(_352_),
    .Y(_109_)
);

INVX1 _728_ (
    .A(_109_),
    .Y(_110_)
);

NOR2X1 _729_ (
    .A(_110_),
    .B(_104_),
    .Y(_111_)
);

OAI21X1 _730_ (
    .A(_111_),
    .B(_108_),
    .C(_105_),
    .Y(_112_)
);

INVX2 _731_ (
    .A(_112_),
    .Y(_113_)
);

NOR2X1 _732_ (
    .A(_244_),
    .B(_540_),
    .Y(_114_)
);

INVX1 _733_ (
    .A(_114_),
    .Y(_115_)
);

NOR2X1 _734_ (
    .A(_115_),
    .B(_101_),
    .Y(_116_)
);

OAI21X1 _735_ (
    .A(_116_),
    .B(_113_),
    .C(_102_),
    .Y(_117_)
);

NAND3X1 _736_ (
    .A(_95_),
    .B(_97_),
    .C(_96_),
    .Y(_118_)
);

AOI21X1 _737_ (
    .A(_118_),
    .B(_117_),
    .C(_98_),
    .Y(_119_)
);

AOI21X1 _738_ (
    .A(_93_),
    .B(_92_),
    .C(_91_),
    .Y(_120_)
);

OAI21X1 _739_ (
    .A(_120_),
    .B(_119_),
    .C(_94_),
    .Y(_121_)
);

NAND3X1 _740_ (
    .A(_86_),
    .B(_121_),
    .C(_89_),
    .Y(_122_)
);

AOI21X1 _741_ (
    .A(_86_),
    .B(_89_),
    .C(_121_),
    .Y(_123_)
);

AOI21X1 _742_ (
    .A(_297_),
    .B(_122_),
    .C(_123_),
    .Y(_124_)
);

NOR2X1 _743_ (
    .A(_287_),
    .B(_319_),
    .Y(_125_)
);

INVX2 _744_ (
    .A(_125_),
    .Y(_126_)
);

AOI21X1 _745_ (
    .A(_330_),
    .B(_69_),
    .C(_88_),
    .Y(_127_)
);

NOR2X1 _746_ (
    .A(_308_),
    .B(_362_),
    .Y(_128_)
);

INVX2 _747_ (
    .A(_128_),
    .Y(_129_)
);

AOI21X1 _748_ (
    .A(_28_),
    .B(_60_),
    .C(_67_),
    .Y(_130_)
);

NOR2X1 _749_ (
    .A(_25_),
    .B(_524_),
    .Y(_131_)
);

INVX2 _750_ (
    .A(_131_),
    .Y(_132_)
);

AOI21X1 _751_ (
    .A(_31_),
    .B(_51_),
    .C(_58_),
    .Y(_133_)
);

NOR2X1 _752_ (
    .A(_540_),
    .B(_559_),
    .Y(_134_)
);

INVX2 _753_ (
    .A(_134_),
    .Y(_135_)
);

AOI21X1 _754_ (
    .A(_34_),
    .B(_40_),
    .C(_49_),
    .Y(_136_)
);

NOR2X1 _755_ (
    .A(_352_),
    .B(_46_),
    .Y(_137_)
);

INVX2 _756_ (
    .A(_137_),
    .Y(_138_)
);

NAND2X1 _757_ (
    .A(breg[7]),
    .B(areg[1]),
    .Y(_139_)
);

NOR2X1 _758_ (
    .A(_37_),
    .B(_139_),
    .Y(_140_)
);

NAND2X1 _759_ (
    .A(areg[1]),
    .B(breg[6]),
    .Y(_141_)
);

NAND2X1 _760_ (
    .A(areg[0]),
    .B(breg[7]),
    .Y(_142_)
);

AND2X2 _761_ (
    .A(_141_),
    .B(_142_),
    .Y(_143_)
);

OAI21X1 _762_ (
    .A(_143_),
    .B(_140_),
    .C(_45_),
    .Y(_144_)
);

AND2X2 _763_ (
    .A(areg[1]),
    .B(breg[6]),
    .Y(_145_)
);

NAND3X1 _764_ (
    .A(_142_),
    .B(_557_),
    .C(_145_),
    .Y(_146_)
);

NAND3X1 _765_ (
    .A(_138_),
    .B(_146_),
    .C(_144_),
    .Y(_147_)
);

AND2X2 _766_ (
    .A(breg[7]),
    .B(areg[1]),
    .Y(_148_)
);

NAND2X1 _767_ (
    .A(_44_),
    .B(_148_),
    .Y(_149_)
);

INVX4 _768_ (
    .A(breg[7]),
    .Y(_150_)
);

OAI21X1 _769_ (
    .A(_243_),
    .B(_150_),
    .C(_141_),
    .Y(_151_)
);

AOI21X1 _770_ (
    .A(_151_),
    .B(_149_),
    .C(_38_),
    .Y(_152_)
);

INVX1 _771_ (
    .A(_146_),
    .Y(_153_)
);

OAI21X1 _772_ (
    .A(_152_),
    .B(_153_),
    .C(_137_),
    .Y(_154_)
);

NAND3X1 _773_ (
    .A(_147_),
    .B(_136_),
    .C(_154_),
    .Y(_155_)
);

OAI21X1 _774_ (
    .A(_48_),
    .B(_35_),
    .C(_42_),
    .Y(_156_)
);

OAI21X1 _775_ (
    .A(_152_),
    .B(_153_),
    .C(_138_),
    .Y(_157_)
);

NAND3X1 _776_ (
    .A(_137_),
    .B(_146_),
    .C(_144_),
    .Y(_158_)
);

NAND3X1 _777_ (
    .A(_158_),
    .B(_156_),
    .C(_157_),
    .Y(_159_)
);

NAND3X1 _778_ (
    .A(_135_),
    .B(_155_),
    .C(_159_),
    .Y(_160_)
);

AOI21X1 _779_ (
    .A(_158_),
    .B(_157_),
    .C(_156_),
    .Y(_161_)
);

AOI21X1 _780_ (
    .A(_147_),
    .B(_154_),
    .C(_136_),
    .Y(_162_)
);

OAI21X1 _781_ (
    .A(_161_),
    .B(_162_),
    .C(_134_),
    .Y(_163_)
);

NAND3X1 _782_ (
    .A(_160_),
    .B(_133_),
    .C(_163_),
    .Y(_164_)
);

OAI21X1 _783_ (
    .A(_57_),
    .B(_32_),
    .C(_55_),
    .Y(_165_)
);

OAI21X1 _784_ (
    .A(_161_),
    .B(_162_),
    .C(_135_),
    .Y(_166_)
);

NAND3X1 _785_ (
    .A(_134_),
    .B(_155_),
    .C(_159_),
    .Y(_167_)
);

NAND3X1 _786_ (
    .A(_167_),
    .B(_165_),
    .C(_166_),
    .Y(_168_)
);

NAND3X1 _787_ (
    .A(_132_),
    .B(_164_),
    .C(_168_),
    .Y(_169_)
);

AOI21X1 _788_ (
    .A(_167_),
    .B(_166_),
    .C(_165_),
    .Y(_170_)
);

AOI21X1 _789_ (
    .A(_160_),
    .B(_163_),
    .C(_133_),
    .Y(_171_)
);

OAI21X1 _790_ (
    .A(_170_),
    .B(_171_),
    .C(_131_),
    .Y(_172_)
);

NAND3X1 _791_ (
    .A(_130_),
    .B(_169_),
    .C(_172_),
    .Y(_173_)
);

OAI21X1 _792_ (
    .A(_66_),
    .B(_29_),
    .C(_64_),
    .Y(_174_)
);

OAI21X1 _793_ (
    .A(_170_),
    .B(_171_),
    .C(_132_),
    .Y(_175_)
);

NAND3X1 _794_ (
    .A(_131_),
    .B(_164_),
    .C(_168_),
    .Y(_176_)
);

NAND3X1 _795_ (
    .A(_176_),
    .B(_174_),
    .C(_175_),
    .Y(_177_)
);

NAND3X1 _796_ (
    .A(_129_),
    .B(_173_),
    .C(_177_),
    .Y(_178_)
);

AOI21X1 _797_ (
    .A(_176_),
    .B(_175_),
    .C(_174_),
    .Y(_179_)
);

AOI21X1 _798_ (
    .A(_169_),
    .B(_172_),
    .C(_130_),
    .Y(_180_)
);

OAI21X1 _799_ (
    .A(_179_),
    .B(_180_),
    .C(_128_),
    .Y(_181_)
);

NAND3X1 _800_ (
    .A(_127_),
    .B(_178_),
    .C(_181_),
    .Y(_182_)
);

OAI21X1 _801_ (
    .A(_87_),
    .B(_341_),
    .C(_85_),
    .Y(_183_)
);

OAI21X1 _802_ (
    .A(_179_),
    .B(_180_),
    .C(_129_),
    .Y(_184_)
);

NAND3X1 _803_ (
    .A(_128_),
    .B(_173_),
    .C(_177_),
    .Y(_185_)
);

NAND3X1 _804_ (
    .A(_185_),
    .B(_183_),
    .C(_184_),
    .Y(_186_)
);

NAND3X1 _805_ (
    .A(_126_),
    .B(_182_),
    .C(_186_),
    .Y(_187_)
);

AOI21X1 _806_ (
    .A(_185_),
    .B(_184_),
    .C(_183_),
    .Y(_188_)
);

AOI21X1 _807_ (
    .A(_178_),
    .B(_181_),
    .C(_127_),
    .Y(_189_)
);

OAI21X1 _808_ (
    .A(_188_),
    .B(_189_),
    .C(_125_),
    .Y(_190_)
);

NAND3X1 _809_ (
    .A(_124_),
    .B(_187_),
    .C(_190_),
    .Y(_191_)
);

OAI21X1 _810_ (
    .A(_87_),
    .B(_88_),
    .C(_341_),
    .Y(_192_)
);

NAND3X1 _811_ (
    .A(_330_),
    .B(_69_),
    .C(_85_),
    .Y(_193_)
);

AOI21X1 _812_ (
    .A(_193_),
    .B(_192_),
    .C(_297_),
    .Y(_194_)
);

NAND3X1 _813_ (
    .A(_297_),
    .B(_193_),
    .C(_192_),
    .Y(_195_)
);

AOI21X1 _814_ (
    .A(_121_),
    .B(_195_),
    .C(_194_),
    .Y(_196_)
);

OAI21X1 _815_ (
    .A(_188_),
    .B(_189_),
    .C(_126_),
    .Y(_197_)
);

NAND3X1 _816_ (
    .A(_125_),
    .B(_182_),
    .C(_186_),
    .Y(_198_)
);

NAND3X1 _817_ (
    .A(_196_),
    .B(_198_),
    .C(_197_),
    .Y(_199_)
);

NAND2X1 _818_ (
    .A(_191_),
    .B(_199_),
    .Y(_200_)
);

XNOR2X1 _819_ (
    .A(_200_),
    .B(_276_),
    .Y(_6_[0])
);

NAND2X1 _820_ (
    .A(_86_),
    .B(_89_),
    .Y(_201_)
);

XNOR2X1 _821_ (
    .A(_201_),
    .B(_297_),
    .Y(_202_)
);

XOR2X1 _822_ (
    .A(_202_),
    .B(_121_),
    .Y(_5_[0])
);

INVX1 _823_ (
    .A(_120_),
    .Y(_203_)
);

NAND2X1 _824_ (
    .A(_94_),
    .B(_203_),
    .Y(_204_)
);

XNOR2X1 _825_ (
    .A(_204_),
    .B(_119_),
    .Y(_4_[0])
);

INVX1 _826_ (
    .A(_98_),
    .Y(_205_)
);

NAND2X1 _827_ (
    .A(_118_),
    .B(_205_),
    .Y(_206_)
);

XOR2X1 _828_ (
    .A(_206_),
    .B(_117_),
    .Y(_3_[0])
);

INVX1 _829_ (
    .A(_116_),
    .Y(_207_)
);

NAND2X1 _830_ (
    .A(_102_),
    .B(_207_),
    .Y(_208_)
);

XNOR2X1 _831_ (
    .A(_208_),
    .B(_113_),
    .Y(_2_[0])
);

INVX1 _832_ (
    .A(_111_),
    .Y(_209_)
);

NAND2X1 _833_ (
    .A(_105_),
    .B(_209_),
    .Y(_210_)
);

XNOR2X1 _834_ (
    .A(_210_),
    .B(_108_),
    .Y(_1_[0])
);

NOR2X1 _835_ (
    .A(_529_),
    .B(_106_),
    .Y(_211_)
);

NOR2X1 _836_ (
    .A(_211_),
    .B(_108_),
    .Y(_7_[0])
);

OAI21X1 _837_ (
    .A(_188_),
    .B(_126_),
    .C(_186_),
    .Y(_212_)
);

NOR2X1 _838_ (
    .A(_362_),
    .B(_287_),
    .Y(_213_)
);

NOR2X1 _839_ (
    .A(_524_),
    .B(_308_),
    .Y(_214_)
);

NOR2X1 _840_ (
    .A(_559_),
    .B(_25_),
    .Y(_215_)
);

INVX1 _841_ (
    .A(_215_),
    .Y(_216_)
);

NOR2X1 _842_ (
    .A(_46_),
    .B(_540_),
    .Y(_217_)
);

AOI22X1 _843_ (
    .A(breg[7]),
    .B(areg[1]),
    .C(breg[6]),
    .D(areg[2]),
    .Y(_218_)
);

NAND2X1 _844_ (
    .A(breg[7]),
    .B(areg[2]),
    .Y(_219_)
);

NOR2X1 _845_ (
    .A(_141_),
    .B(_219_),
    .Y(_220_)
);

OAI21X1 _846_ (
    .A(_220_),
    .B(_218_),
    .C(_149_),
    .Y(_221_)
);

NAND2X1 _847_ (
    .A(breg[6]),
    .B(areg[2]),
    .Y(_222_)
);

NAND3X1 _848_ (
    .A(_222_),
    .B(_44_),
    .C(_148_),
    .Y(_223_)
);

NAND3X1 _849_ (
    .A(_217_),
    .B(_223_),
    .C(_221_),
    .Y(_224_)
);

INVX1 _850_ (
    .A(_217_),
    .Y(_225_)
);

OAI21X1 _851_ (
    .A(_220_),
    .B(_218_),
    .C(_140_),
    .Y(_226_)
);

INVX1 _852_ (
    .A(_218_),
    .Y(_227_)
);

OR2X2 _853_ (
    .A(_139_),
    .B(_222_),
    .Y(_228_)
);

NAND3X1 _854_ (
    .A(_227_),
    .B(_149_),
    .C(_228_),
    .Y(_229_)
);

NAND3X1 _855_ (
    .A(_225_),
    .B(_226_),
    .C(_229_),
    .Y(_230_)
);

OAI21X1 _856_ (
    .A(_352_),
    .B(_46_),
    .C(_146_),
    .Y(_231_)
);

NAND2X1 _857_ (
    .A(_231_),
    .B(_144_),
    .Y(_232_)
);

NAND3X1 _858_ (
    .A(_224_),
    .B(_232_),
    .C(_230_),
    .Y(_233_)
);

NAND3X1 _859_ (
    .A(_225_),
    .B(_223_),
    .C(_221_),
    .Y(_234_)
);

NAND3X1 _860_ (
    .A(_217_),
    .B(_226_),
    .C(_229_),
    .Y(_235_)
);

OAI21X1 _861_ (
    .A(_152_),
    .B(_138_),
    .C(_146_),
    .Y(_236_)
);

NAND3X1 _862_ (
    .A(_234_),
    .B(_235_),
    .C(_236_),
    .Y(_237_)
);

AOI21X1 _863_ (
    .A(_233_),
    .B(_237_),
    .C(_216_),
    .Y(_238_)
);

NAND3X1 _864_ (
    .A(_234_),
    .B(_232_),
    .C(_235_),
    .Y(_239_)
);

NAND3X1 _865_ (
    .A(_224_),
    .B(_230_),
    .C(_236_),
    .Y(_240_)
);

AOI21X1 _866_ (
    .A(_239_),
    .B(_240_),
    .C(_215_),
    .Y(_241_)
);

AOI21X1 _867_ (
    .A(_134_),
    .B(_155_),
    .C(_162_),
    .Y(_242_)
);

OAI21X1 _868_ (
    .A(_238_),
    .B(_241_),
    .C(_242_),
    .Y(_245_)
);

NAND3X1 _869_ (
    .A(_215_),
    .B(_239_),
    .C(_240_),
    .Y(_246_)
);

NAND3X1 _870_ (
    .A(_216_),
    .B(_233_),
    .C(_237_),
    .Y(_247_)
);

OAI21X1 _871_ (
    .A(_161_),
    .B(_135_),
    .C(_159_),
    .Y(_248_)
);

NAND3X1 _872_ (
    .A(_246_),
    .B(_247_),
    .C(_248_),
    .Y(_249_)
);

NAND3X1 _873_ (
    .A(_214_),
    .B(_249_),
    .C(_245_),
    .Y(_250_)
);

INVX2 _874_ (
    .A(_214_),
    .Y(_251_)
);

NAND3X1 _875_ (
    .A(_246_),
    .B(_247_),
    .C(_242_),
    .Y(_252_)
);

OAI21X1 _876_ (
    .A(_238_),
    .B(_241_),
    .C(_248_),
    .Y(_253_)
);

NAND3X1 _877_ (
    .A(_251_),
    .B(_252_),
    .C(_253_),
    .Y(_254_)
);

AOI21X1 _878_ (
    .A(_131_),
    .B(_164_),
    .C(_171_),
    .Y(_255_)
);

AOI21X1 _879_ (
    .A(_250_),
    .B(_254_),
    .C(_255_),
    .Y(_256_)
);

NAND3X1 _880_ (
    .A(_251_),
    .B(_249_),
    .C(_245_),
    .Y(_257_)
);

NAND3X1 _881_ (
    .A(_214_),
    .B(_252_),
    .C(_253_),
    .Y(_258_)
);

OAI21X1 _882_ (
    .A(_170_),
    .B(_132_),
    .C(_168_),
    .Y(_259_)
);

AOI21X1 _883_ (
    .A(_257_),
    .B(_258_),
    .C(_259_),
    .Y(_260_)
);

OAI21X1 _884_ (
    .A(_260_),
    .B(_256_),
    .C(_213_),
    .Y(_261_)
);

INVX2 _885_ (
    .A(_213_),
    .Y(_262_)
);

AOI21X1 _886_ (
    .A(_252_),
    .B(_253_),
    .C(_251_),
    .Y(_263_)
);

AOI21X1 _887_ (
    .A(_249_),
    .B(_245_),
    .C(_214_),
    .Y(_264_)
);

OAI21X1 _888_ (
    .A(_263_),
    .B(_264_),
    .C(_259_),
    .Y(_266_)
);

NAND3X1 _889_ (
    .A(_250_),
    .B(_254_),
    .C(_255_),
    .Y(_267_)
);

NAND3X1 _890_ (
    .A(_262_),
    .B(_267_),
    .C(_266_),
    .Y(_268_)
);

AOI21X1 _891_ (
    .A(_128_),
    .B(_173_),
    .C(_180_),
    .Y(_269_)
);

NAND3X1 _892_ (
    .A(_268_),
    .B(_261_),
    .C(_269_),
    .Y(_270_)
);

AOI21X1 _893_ (
    .A(_267_),
    .B(_266_),
    .C(_262_),
    .Y(_271_)
);

NOR3X1 _894_ (
    .A(_256_),
    .B(_213_),
    .C(_260_),
    .Y(_272_)
);

OAI21X1 _895_ (
    .A(_179_),
    .B(_129_),
    .C(_177_),
    .Y(_273_)
);

OAI21X1 _896_ (
    .A(_272_),
    .B(_271_),
    .C(_273_),
    .Y(_274_)
);

NOR2X1 _897_ (
    .A(_319_),
    .B(_265_),
    .Y(_275_)
);

AOI21X1 _898_ (
    .A(_270_),
    .B(_274_),
    .C(_275_),
    .Y(_277_)
);

OAI21X1 _899_ (
    .A(_260_),
    .B(_256_),
    .C(_262_),
    .Y(_278_)
);

NAND3X1 _900_ (
    .A(_213_),
    .B(_267_),
    .C(_266_),
    .Y(_279_)
);

NAND3X1 _901_ (
    .A(_279_),
    .B(_278_),
    .C(_269_),
    .Y(_280_)
);

NAND3X1 _902_ (
    .A(_261_),
    .B(_268_),
    .C(_273_),
    .Y(_281_)
);

INVX2 _903_ (
    .A(_275_),
    .Y(_282_)
);

AOI21X1 _904_ (
    .A(_280_),
    .B(_281_),
    .C(_282_),
    .Y(_283_)
);

OAI21X1 _905_ (
    .A(_277_),
    .B(_283_),
    .C(_212_),
    .Y(_284_)
);

AOI21X1 _906_ (
    .A(_125_),
    .B(_182_),
    .C(_189_),
    .Y(_285_)
);

NAND3X1 _907_ (
    .A(_282_),
    .B(_280_),
    .C(_281_),
    .Y(_286_)
);

NAND3X1 _908_ (
    .A(_270_),
    .B(_275_),
    .C(_274_),
    .Y(_288_)
);

NAND3X1 _909_ (
    .A(_286_),
    .B(_285_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _910_ (
    .A(_289_),
    .B(_284_),
    .Y(_290_)
);

AOI21X1 _911_ (
    .A(_187_),
    .B(_190_),
    .C(_124_),
    .Y(_291_)
);

AOI21X1 _912_ (
    .A(_276_),
    .B(_191_),
    .C(_291_),
    .Y(_292_)
);

XOR2X1 _913_ (
    .A(_292_),
    .B(_290_),
    .Y(_9_[8])
);

NAND2X1 _914_ (
    .A(_270_),
    .B(_274_),
    .Y(_293_)
);

OAI21X1 _915_ (
    .A(_212_),
    .B(_275_),
    .C(_293_),
    .Y(_294_)
);

OAI21X1 _916_ (
    .A(_285_),
    .B(_282_),
    .C(_294_),
    .Y(_295_)
);

NOR2X1 _917_ (
    .A(_362_),
    .B(_265_),
    .Y(_296_)
);

INVX1 _918_ (
    .A(_296_),
    .Y(_298_)
);

NOR2X1 _919_ (
    .A(_524_),
    .B(_287_),
    .Y(_299_)
);

NOR2X1 _920_ (
    .A(_559_),
    .B(_308_),
    .Y(_300_)
);

NAND2X1 _921_ (
    .A(_230_),
    .B(_236_),
    .Y(_301_)
);

NOR2X1 _922_ (
    .A(_46_),
    .B(_25_),
    .Y(_302_)
);

OAI21X1 _923_ (
    .A(_141_),
    .B(_219_),
    .C(_149_),
    .Y(_303_)
);

NAND2X1 _924_ (
    .A(breg[7]),
    .B(areg[3]),
    .Y(_304_)
);

INVX4 _925_ (
    .A(breg[6]),
    .Y(_305_)
);

OAI21X1 _926_ (
    .A(_305_),
    .B(_540_),
    .C(_219_),
    .Y(_306_)
);

OAI21X1 _927_ (
    .A(_222_),
    .B(_304_),
    .C(_306_),
    .Y(_307_)
);

XNOR2X1 _928_ (
    .A(_303_),
    .B(_307_),
    .Y(_309_)
);

NAND2X1 _929_ (
    .A(_302_),
    .B(_309_),
    .Y(_310_)
);

XOR2X1 _930_ (
    .A(_303_),
    .B(_307_),
    .Y(_311_)
);

OAI21X1 _931_ (
    .A(_46_),
    .B(_25_),
    .C(_311_),
    .Y(_312_)
);

NAND2X1 _932_ (
    .A(_310_),
    .B(_312_),
    .Y(_313_)
);

NAND3X1 _933_ (
    .A(_224_),
    .B(_301_),
    .C(_313_),
    .Y(_314_)
);

NAND2X1 _934_ (
    .A(_224_),
    .B(_301_),
    .Y(_315_)
);

NAND3X1 _935_ (
    .A(_310_),
    .B(_312_),
    .C(_315_),
    .Y(_316_)
);

NAND3X1 _936_ (
    .A(_300_),
    .B(_316_),
    .C(_314_),
    .Y(_317_)
);

INVX1 _937_ (
    .A(_300_),
    .Y(_318_)
);

OR2X2 _938_ (
    .A(_313_),
    .B(_315_),
    .Y(_320_)
);

NAND2X1 _939_ (
    .A(_315_),
    .B(_313_),
    .Y(_321_)
);

NAND3X1 _940_ (
    .A(_318_),
    .B(_321_),
    .C(_320_),
    .Y(_322_)
);

OAI21X1 _941_ (
    .A(_242_),
    .B(_241_),
    .C(_246_),
    .Y(_323_)
);

INVX2 _942_ (
    .A(_323_),
    .Y(_324_)
);

AOI21X1 _943_ (
    .A(_317_),
    .B(_322_),
    .C(_324_),
    .Y(_325_)
);

NAND3X1 _944_ (
    .A(_318_),
    .B(_316_),
    .C(_314_),
    .Y(_326_)
);

NAND3X1 _945_ (
    .A(_300_),
    .B(_321_),
    .C(_320_),
    .Y(_327_)
);

AOI21X1 _946_ (
    .A(_326_),
    .B(_327_),
    .C(_323_),
    .Y(_328_)
);

OAI21X1 _947_ (
    .A(_325_),
    .B(_328_),
    .C(_299_),
    .Y(_329_)
);

INVX1 _948_ (
    .A(_299_),
    .Y(_331_)
);

NAND3X1 _949_ (
    .A(_326_),
    .B(_323_),
    .C(_327_),
    .Y(_332_)
);

NAND3X1 _950_ (
    .A(_317_),
    .B(_324_),
    .C(_322_),
    .Y(_333_)
);

NAND3X1 _951_ (
    .A(_331_),
    .B(_333_),
    .C(_332_),
    .Y(_334_)
);

OAI21X1 _952_ (
    .A(_259_),
    .B(_263_),
    .C(_254_),
    .Y(_335_)
);

NAND3X1 _953_ (
    .A(_334_),
    .B(_335_),
    .C(_329_),
    .Y(_336_)
);

AOI21X1 _954_ (
    .A(_333_),
    .B(_332_),
    .C(_331_),
    .Y(_337_)
);

NOR3X1 _955_ (
    .A(_325_),
    .B(_299_),
    .C(_328_),
    .Y(_338_)
);

INVX1 _956_ (
    .A(_335_),
    .Y(_339_)
);

OAI21X1 _957_ (
    .A(_338_),
    .B(_337_),
    .C(_339_),
    .Y(_340_)
);

AOI21X1 _958_ (
    .A(_336_),
    .B(_340_),
    .C(_298_),
    .Y(_342_)
);

OAI21X1 _959_ (
    .A(_338_),
    .B(_337_),
    .C(_335_),
    .Y(_343_)
);

NAND3X1 _960_ (
    .A(_334_),
    .B(_339_),
    .C(_329_),
    .Y(_344_)
);

AOI21X1 _961_ (
    .A(_344_),
    .B(_343_),
    .C(_296_),
    .Y(_345_)
);

OAI21X1 _962_ (
    .A(_272_),
    .B(_269_),
    .C(_261_),
    .Y(_346_)
);

INVX1 _963_ (
    .A(_346_),
    .Y(_347_)
);

OAI21X1 _964_ (
    .A(_342_),
    .B(_345_),
    .C(_347_),
    .Y(_348_)
);

NAND3X1 _965_ (
    .A(_296_),
    .B(_344_),
    .C(_343_),
    .Y(_349_)
);

NAND3X1 _966_ (
    .A(_298_),
    .B(_336_),
    .C(_340_),
    .Y(_350_)
);

NAND3X1 _967_ (
    .A(_346_),
    .B(_349_),
    .C(_350_),
    .Y(_351_)
);

NAND2X1 _968_ (
    .A(_351_),
    .B(_348_),
    .Y(_353_)
);

OAI21X1 _969_ (
    .A(_292_),
    .B(_290_),
    .C(_353_),
    .Y(_354_)
);

AND2X2 _970_ (
    .A(_284_),
    .B(_289_),
    .Y(_355_)
);

INVX1 _971_ (
    .A(_276_),
    .Y(_356_)
);

AOI21X1 _972_ (
    .A(_198_),
    .B(_197_),
    .C(_196_),
    .Y(_357_)
);

OAI21X1 _973_ (
    .A(_357_),
    .B(_356_),
    .C(_199_),
    .Y(_358_)
);

AND2X2 _974_ (
    .A(_348_),
    .B(_351_),
    .Y(_359_)
);

NAND3X1 _975_ (
    .A(_355_),
    .B(_358_),
    .C(_359_),
    .Y(_360_)
);

NAND2X1 _976_ (
    .A(_354_),
    .B(_360_),
    .Y(_361_)
);

XNOR2X1 _977_ (
    .A(_361_),
    .B(_295_),
    .Y(_9_[9])
);

OAI21X1 _978_ (
    .A(_345_),
    .B(_347_),
    .C(_349_),
    .Y(_363_)
);

NAND2X1 _979_ (
    .A(_295_),
    .B(_354_),
    .Y(_364_)
);

NOR2X1 _980_ (
    .A(_524_),
    .B(_265_),
    .Y(_365_)
);

INVX1 _981_ (
    .A(_365_),
    .Y(_366_)
);

NOR2X1 _982_ (
    .A(_559_),
    .B(_287_),
    .Y(_367_)
);

NOR2X1 _983_ (
    .A(_46_),
    .B(_308_),
    .Y(_368_)
);

NAND2X1 _984_ (
    .A(breg[6]),
    .B(areg[3]),
    .Y(_369_)
);

AOI21X1 _985_ (
    .A(_149_),
    .B(_228_),
    .C(_369_),
    .Y(_370_)
);

OAI21X1 _986_ (
    .A(_219_),
    .B(_369_),
    .C(_228_),
    .Y(_371_)
);

OR2X2 _987_ (
    .A(_370_),
    .B(_371_),
    .Y(_372_)
);

NOR2X1 _988_ (
    .A(_305_),
    .B(_25_),
    .Y(_374_)
);

XNOR2X1 _989_ (
    .A(_372_),
    .B(_374_),
    .Y(_375_)
);

XOR2X1 _990_ (
    .A(_375_),
    .B(_304_),
    .Y(_376_)
);

XNOR2X1 _991_ (
    .A(_376_),
    .B(_368_),
    .Y(_377_)
);

OAI21X1 _992_ (
    .A(_302_),
    .B(_309_),
    .C(_315_),
    .Y(_378_)
);

NAND2X1 _993_ (
    .A(_310_),
    .B(_378_),
    .Y(_379_)
);

XNOR2X1 _994_ (
    .A(_377_),
    .B(_379_),
    .Y(_380_)
);

NAND2X1 _995_ (
    .A(_367_),
    .B(_380_),
    .Y(_381_)
);

OR2X2 _996_ (
    .A(_380_),
    .B(_367_),
    .Y(_382_)
);

NAND2X1 _997_ (
    .A(_321_),
    .B(_320_),
    .Y(_383_)
);

NAND2X1 _998_ (
    .A(_324_),
    .B(_317_),
    .Y(_385_)
);

OAI21X1 _999_ (
    .A(_300_),
    .B(_383_),
    .C(_385_),
    .Y(_386_)
);

endmodule
